magic
tech sky130A
magscale 1 2
timestamp 1672517212
<< obsli1 >>
rect 1104 2159 48852 51697
<< obsm1 >>
rect 1026 2128 48852 51728
<< metal2 >>
rect 1030 53200 1086 54000
rect 2870 53200 2926 54000
rect 4710 53200 4766 54000
rect 6550 53200 6606 54000
rect 8390 53200 8446 54000
rect 10230 53200 10286 54000
rect 12070 53200 12126 54000
rect 13910 53200 13966 54000
rect 15750 53200 15806 54000
rect 17590 53200 17646 54000
rect 19430 53200 19486 54000
rect 21270 53200 21326 54000
rect 23110 53200 23166 54000
rect 24950 53200 25006 54000
rect 26790 53200 26846 54000
rect 28630 53200 28686 54000
rect 30470 53200 30526 54000
rect 32310 53200 32366 54000
rect 34150 53200 34206 54000
rect 35990 53200 36046 54000
rect 37830 53200 37886 54000
rect 39670 53200 39726 54000
rect 41510 53200 41566 54000
rect 43350 53200 43406 54000
rect 45190 53200 45246 54000
rect 47030 53200 47086 54000
rect 48870 53200 48926 54000
<< obsm2 >>
rect 1142 53144 2814 53258
rect 2982 53144 4654 53258
rect 4822 53144 6494 53258
rect 6662 53144 8334 53258
rect 8502 53144 10174 53258
rect 10342 53144 12014 53258
rect 12182 53144 13854 53258
rect 14022 53144 15694 53258
rect 15862 53144 17534 53258
rect 17702 53144 19374 53258
rect 19542 53144 21214 53258
rect 21382 53144 23054 53258
rect 23222 53144 24894 53258
rect 25062 53144 26734 53258
rect 26902 53144 28574 53258
rect 28742 53144 30414 53258
rect 30582 53144 32254 53258
rect 32422 53144 34094 53258
rect 34262 53144 35934 53258
rect 36102 53144 37774 53258
rect 37942 53144 39614 53258
rect 39782 53144 41454 53258
rect 41622 53144 43294 53258
rect 43462 53144 45134 53258
rect 45302 53144 46974 53258
rect 47142 53144 48374 53258
rect 1032 1799 48374 53144
<< metal3 >>
rect 0 51960 800 52080
rect 0 50736 800 50856
rect 49200 50872 50000 50992
rect 49200 49784 50000 49904
rect 0 49512 800 49632
rect 49200 48696 50000 48816
rect 0 48288 800 48408
rect 49200 47608 50000 47728
rect 0 47064 800 47184
rect 49200 46520 50000 46640
rect 0 45840 800 45960
rect 49200 45432 50000 45552
rect 0 44616 800 44736
rect 49200 44344 50000 44464
rect 0 43392 800 43512
rect 49200 43256 50000 43376
rect 0 42168 800 42288
rect 49200 42168 50000 42288
rect 0 40944 800 41064
rect 49200 41080 50000 41200
rect 49200 39992 50000 40112
rect 0 39720 800 39840
rect 49200 38904 50000 39024
rect 0 38496 800 38616
rect 49200 37816 50000 37936
rect 0 37272 800 37392
rect 49200 36728 50000 36848
rect 0 36048 800 36168
rect 49200 35640 50000 35760
rect 0 34824 800 34944
rect 49200 34552 50000 34672
rect 0 33600 800 33720
rect 49200 33464 50000 33584
rect 0 32376 800 32496
rect 49200 32376 50000 32496
rect 0 31152 800 31272
rect 49200 31288 50000 31408
rect 49200 30200 50000 30320
rect 0 29928 800 30048
rect 49200 29112 50000 29232
rect 0 28704 800 28824
rect 49200 28024 50000 28144
rect 0 27480 800 27600
rect 49200 26936 50000 27056
rect 0 26256 800 26376
rect 49200 25848 50000 25968
rect 0 25032 800 25152
rect 49200 24760 50000 24880
rect 0 23808 800 23928
rect 49200 23672 50000 23792
rect 0 22584 800 22704
rect 49200 22584 50000 22704
rect 0 21360 800 21480
rect 49200 21496 50000 21616
rect 49200 20408 50000 20528
rect 0 20136 800 20256
rect 49200 19320 50000 19440
rect 0 18912 800 19032
rect 49200 18232 50000 18352
rect 0 17688 800 17808
rect 49200 17144 50000 17264
rect 0 16464 800 16584
rect 49200 16056 50000 16176
rect 0 15240 800 15360
rect 49200 14968 50000 15088
rect 0 14016 800 14136
rect 49200 13880 50000 14000
rect 0 12792 800 12912
rect 49200 12792 50000 12912
rect 0 11568 800 11688
rect 49200 11704 50000 11824
rect 49200 10616 50000 10736
rect 0 10344 800 10464
rect 49200 9528 50000 9648
rect 0 9120 800 9240
rect 49200 8440 50000 8560
rect 0 7896 800 8016
rect 49200 7352 50000 7472
rect 0 6672 800 6792
rect 49200 6264 50000 6384
rect 0 5448 800 5568
rect 49200 5176 50000 5296
rect 0 4224 800 4344
rect 49200 4088 50000 4208
rect 0 3000 800 3120
rect 49200 3000 50000 3120
rect 0 1776 800 1896
<< obsm3 >>
rect 800 51072 49200 51713
rect 800 50936 49120 51072
rect 880 50792 49120 50936
rect 880 50656 49200 50792
rect 800 49984 49200 50656
rect 800 49712 49120 49984
rect 880 49704 49120 49712
rect 880 49432 49200 49704
rect 800 48896 49200 49432
rect 800 48616 49120 48896
rect 800 48488 49200 48616
rect 880 48208 49200 48488
rect 800 47808 49200 48208
rect 800 47528 49120 47808
rect 800 47264 49200 47528
rect 880 46984 49200 47264
rect 800 46720 49200 46984
rect 800 46440 49120 46720
rect 800 46040 49200 46440
rect 880 45760 49200 46040
rect 800 45632 49200 45760
rect 800 45352 49120 45632
rect 800 44816 49200 45352
rect 880 44544 49200 44816
rect 880 44536 49120 44544
rect 800 44264 49120 44536
rect 800 43592 49200 44264
rect 880 43456 49200 43592
rect 880 43312 49120 43456
rect 800 43176 49120 43312
rect 800 42368 49200 43176
rect 880 42088 49120 42368
rect 800 41280 49200 42088
rect 800 41144 49120 41280
rect 880 41000 49120 41144
rect 880 40864 49200 41000
rect 800 40192 49200 40864
rect 800 39920 49120 40192
rect 880 39912 49120 39920
rect 880 39640 49200 39912
rect 800 39104 49200 39640
rect 800 38824 49120 39104
rect 800 38696 49200 38824
rect 880 38416 49200 38696
rect 800 38016 49200 38416
rect 800 37736 49120 38016
rect 800 37472 49200 37736
rect 880 37192 49200 37472
rect 800 36928 49200 37192
rect 800 36648 49120 36928
rect 800 36248 49200 36648
rect 880 35968 49200 36248
rect 800 35840 49200 35968
rect 800 35560 49120 35840
rect 800 35024 49200 35560
rect 880 34752 49200 35024
rect 880 34744 49120 34752
rect 800 34472 49120 34744
rect 800 33800 49200 34472
rect 880 33664 49200 33800
rect 880 33520 49120 33664
rect 800 33384 49120 33520
rect 800 32576 49200 33384
rect 880 32296 49120 32576
rect 800 31488 49200 32296
rect 800 31352 49120 31488
rect 880 31208 49120 31352
rect 880 31072 49200 31208
rect 800 30400 49200 31072
rect 800 30128 49120 30400
rect 880 30120 49120 30128
rect 880 29848 49200 30120
rect 800 29312 49200 29848
rect 800 29032 49120 29312
rect 800 28904 49200 29032
rect 880 28624 49200 28904
rect 800 28224 49200 28624
rect 800 27944 49120 28224
rect 800 27680 49200 27944
rect 880 27400 49200 27680
rect 800 27136 49200 27400
rect 800 26856 49120 27136
rect 800 26456 49200 26856
rect 880 26176 49200 26456
rect 800 26048 49200 26176
rect 800 25768 49120 26048
rect 800 25232 49200 25768
rect 880 24960 49200 25232
rect 880 24952 49120 24960
rect 800 24680 49120 24952
rect 800 24008 49200 24680
rect 880 23872 49200 24008
rect 880 23728 49120 23872
rect 800 23592 49120 23728
rect 800 22784 49200 23592
rect 880 22504 49120 22784
rect 800 21696 49200 22504
rect 800 21560 49120 21696
rect 880 21416 49120 21560
rect 880 21280 49200 21416
rect 800 20608 49200 21280
rect 800 20336 49120 20608
rect 880 20328 49120 20336
rect 880 20056 49200 20328
rect 800 19520 49200 20056
rect 800 19240 49120 19520
rect 800 19112 49200 19240
rect 880 18832 49200 19112
rect 800 18432 49200 18832
rect 800 18152 49120 18432
rect 800 17888 49200 18152
rect 880 17608 49200 17888
rect 800 17344 49200 17608
rect 800 17064 49120 17344
rect 800 16664 49200 17064
rect 880 16384 49200 16664
rect 800 16256 49200 16384
rect 800 15976 49120 16256
rect 800 15440 49200 15976
rect 880 15168 49200 15440
rect 880 15160 49120 15168
rect 800 14888 49120 15160
rect 800 14216 49200 14888
rect 880 14080 49200 14216
rect 880 13936 49120 14080
rect 800 13800 49120 13936
rect 800 12992 49200 13800
rect 880 12712 49120 12992
rect 800 11904 49200 12712
rect 800 11768 49120 11904
rect 880 11624 49120 11768
rect 880 11488 49200 11624
rect 800 10816 49200 11488
rect 800 10544 49120 10816
rect 880 10536 49120 10544
rect 880 10264 49200 10536
rect 800 9728 49200 10264
rect 800 9448 49120 9728
rect 800 9320 49200 9448
rect 880 9040 49200 9320
rect 800 8640 49200 9040
rect 800 8360 49120 8640
rect 800 8096 49200 8360
rect 880 7816 49200 8096
rect 800 7552 49200 7816
rect 800 7272 49120 7552
rect 800 6872 49200 7272
rect 880 6592 49200 6872
rect 800 6464 49200 6592
rect 800 6184 49120 6464
rect 800 5648 49200 6184
rect 880 5376 49200 5648
rect 880 5368 49120 5376
rect 800 5096 49120 5368
rect 800 4424 49200 5096
rect 880 4288 49200 4424
rect 880 4144 49120 4288
rect 800 4008 49120 4144
rect 800 3200 49200 4008
rect 880 2920 49120 3200
rect 800 1976 49200 2920
rect 880 1803 49200 1976
<< metal4 >>
rect 4208 2128 4528 51728
rect 19568 2128 19888 51728
rect 34928 2128 35248 51728
<< labels >>
rlabel metal3 s 49200 3000 50000 3120 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 49200 35640 50000 35760 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 49200 38904 50000 39024 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 49200 42168 50000 42288 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 45432 50000 45552 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 49200 48696 50000 48816 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 48870 53200 48926 54000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 43350 53200 43406 54000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 37830 53200 37886 54000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 32310 53200 32366 54000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 26790 53200 26846 54000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 49200 6264 50000 6384 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 21270 53200 21326 54000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 15750 53200 15806 54000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 10230 53200 10286 54000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 4710 53200 4766 54000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 49200 9528 50000 9648 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 49200 12792 50000 12912 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 49200 16056 50000 16176 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 49200 19320 50000 19440 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 49200 22584 50000 22704 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 49200 25848 50000 25968 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 49200 29112 50000 29232 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 49200 32376 50000 32496 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 49200 5176 50000 5296 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 49200 37816 50000 37936 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 49200 41080 50000 41200 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 49200 44344 50000 44464 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 49200 47608 50000 47728 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 49200 50872 50000 50992 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 45190 53200 45246 54000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39670 53200 39726 54000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 34150 53200 34206 54000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 28630 53200 28686 54000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 23110 53200 23166 54000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 49200 8440 50000 8560 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 17590 53200 17646 54000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 12070 53200 12126 54000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 6550 53200 6606 54000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 1030 53200 1086 54000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 49200 11704 50000 11824 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 49200 14968 50000 15088 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 49200 18232 50000 18352 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 49200 21496 50000 21616 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 49200 24760 50000 24880 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 49200 28024 50000 28144 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 49200 31288 50000 31408 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 49200 34552 50000 34672 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 49200 4088 50000 4208 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 49200 36728 50000 36848 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 49200 39992 50000 40112 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 49200 43256 50000 43376 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 49200 46520 50000 46640 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 49200 49784 50000 49904 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 47030 53200 47086 54000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 41510 53200 41566 54000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 35990 53200 36046 54000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 30470 53200 30526 54000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 24950 53200 25006 54000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 49200 7352 50000 7472 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 19430 53200 19486 54000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 13910 53200 13966 54000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 8390 53200 8446 54000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 2870 53200 2926 54000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 49200 10616 50000 10736 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 49200 13880 50000 14000 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 49200 17144 50000 17264 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 49200 20408 50000 20528 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 49200 23672 50000 23792 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 49200 26936 50000 27056 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 49200 30200 50000 30320 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 49200 33464 50000 33584 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4208 2128 4528 51728 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 51728 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 51728 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 50000 54000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 739722
string GDS_FILE /home/runner/work/tiny_user_project_vgaclock_mpw8/tiny_user_project_vgaclock_mpw8/openlane/tiny_user_project/runs/22_12_31_20_05/results/signoff/tiny_user_project.magic.gds
string GDS_START 23768
<< end >>

