VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 270.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 15.000 250.000 15.600 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 178.200 250.000 178.800 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 194.520 250.000 195.120 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 210.840 250.000 211.440 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 227.160 250.000 227.760 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 243.480 250.000 244.080 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 266.000 244.630 270.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 266.000 217.030 270.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 266.000 189.430 270.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 266.000 161.830 270.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 266.000 134.230 270.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 31.320 250.000 31.920 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 266.000 106.630 270.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 266.000 79.030 270.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 266.000 51.430 270.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 266.000 23.830 270.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 47.640 250.000 48.240 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 63.960 250.000 64.560 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 80.280 250.000 80.880 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 96.600 250.000 97.200 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 112.920 250.000 113.520 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 129.240 250.000 129.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 145.560 250.000 146.160 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 161.880 250.000 162.480 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 25.880 250.000 26.480 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 189.080 250.000 189.680 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 205.400 250.000 206.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 221.720 250.000 222.320 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 238.040 250.000 238.640 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 254.360 250.000 254.960 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 266.000 226.230 270.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 266.000 198.630 270.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 266.000 171.030 270.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 266.000 143.430 270.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 266.000 115.830 270.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 42.200 250.000 42.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 266.000 88.230 270.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 266.000 60.630 270.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 266.000 33.030 270.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 266.000 5.430 270.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 58.520 250.000 59.120 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 74.840 250.000 75.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 91.160 250.000 91.760 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 107.480 250.000 108.080 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 123.800 250.000 124.400 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 140.120 250.000 140.720 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 156.440 250.000 157.040 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 172.760 250.000 173.360 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 20.440 250.000 21.040 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 183.640 250.000 184.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 199.960 250.000 200.560 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 216.280 250.000 216.880 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 232.600 250.000 233.200 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 248.920 250.000 249.520 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 266.000 235.430 270.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 266.000 207.830 270.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 266.000 180.230 270.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 266.000 152.630 270.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 266.000 125.030 270.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 36.760 250.000 37.360 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 266.000 97.430 270.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 266.000 69.830 270.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 266.000 42.230 270.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 266.000 14.630 270.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 53.080 250.000 53.680 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 69.400 250.000 70.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 85.720 250.000 86.320 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 102.040 250.000 102.640 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 118.360 250.000 118.960 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 134.680 250.000 135.280 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 151.000 250.000 151.600 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 167.320 250.000 167.920 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 258.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 258.640 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 258.640 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 258.485 ;
      LAYER met1 ;
        RECT 5.130 10.640 244.260 258.640 ;
      LAYER met2 ;
        RECT 5.710 265.720 14.070 266.290 ;
        RECT 14.910 265.720 23.270 266.290 ;
        RECT 24.110 265.720 32.470 266.290 ;
        RECT 33.310 265.720 41.670 266.290 ;
        RECT 42.510 265.720 50.870 266.290 ;
        RECT 51.710 265.720 60.070 266.290 ;
        RECT 60.910 265.720 69.270 266.290 ;
        RECT 70.110 265.720 78.470 266.290 ;
        RECT 79.310 265.720 87.670 266.290 ;
        RECT 88.510 265.720 96.870 266.290 ;
        RECT 97.710 265.720 106.070 266.290 ;
        RECT 106.910 265.720 115.270 266.290 ;
        RECT 116.110 265.720 124.470 266.290 ;
        RECT 125.310 265.720 133.670 266.290 ;
        RECT 134.510 265.720 142.870 266.290 ;
        RECT 143.710 265.720 152.070 266.290 ;
        RECT 152.910 265.720 161.270 266.290 ;
        RECT 162.110 265.720 170.470 266.290 ;
        RECT 171.310 265.720 179.670 266.290 ;
        RECT 180.510 265.720 188.870 266.290 ;
        RECT 189.710 265.720 198.070 266.290 ;
        RECT 198.910 265.720 207.270 266.290 ;
        RECT 208.110 265.720 216.470 266.290 ;
        RECT 217.310 265.720 225.670 266.290 ;
        RECT 226.510 265.720 234.870 266.290 ;
        RECT 235.710 265.720 241.870 266.290 ;
        RECT 5.160 8.995 241.870 265.720 ;
      LAYER met3 ;
        RECT 4.000 255.360 246.000 258.565 ;
        RECT 4.000 254.680 245.600 255.360 ;
        RECT 4.400 253.960 245.600 254.680 ;
        RECT 4.400 253.280 246.000 253.960 ;
        RECT 4.000 249.920 246.000 253.280 ;
        RECT 4.000 248.560 245.600 249.920 ;
        RECT 4.400 248.520 245.600 248.560 ;
        RECT 4.400 247.160 246.000 248.520 ;
        RECT 4.000 244.480 246.000 247.160 ;
        RECT 4.000 243.080 245.600 244.480 ;
        RECT 4.000 242.440 246.000 243.080 ;
        RECT 4.400 241.040 246.000 242.440 ;
        RECT 4.000 239.040 246.000 241.040 ;
        RECT 4.000 237.640 245.600 239.040 ;
        RECT 4.000 236.320 246.000 237.640 ;
        RECT 4.400 234.920 246.000 236.320 ;
        RECT 4.000 233.600 246.000 234.920 ;
        RECT 4.000 232.200 245.600 233.600 ;
        RECT 4.000 230.200 246.000 232.200 ;
        RECT 4.400 228.800 246.000 230.200 ;
        RECT 4.000 228.160 246.000 228.800 ;
        RECT 4.000 226.760 245.600 228.160 ;
        RECT 4.000 224.080 246.000 226.760 ;
        RECT 4.400 222.720 246.000 224.080 ;
        RECT 4.400 222.680 245.600 222.720 ;
        RECT 4.000 221.320 245.600 222.680 ;
        RECT 4.000 217.960 246.000 221.320 ;
        RECT 4.400 217.280 246.000 217.960 ;
        RECT 4.400 216.560 245.600 217.280 ;
        RECT 4.000 215.880 245.600 216.560 ;
        RECT 4.000 211.840 246.000 215.880 ;
        RECT 4.400 210.440 245.600 211.840 ;
        RECT 4.000 206.400 246.000 210.440 ;
        RECT 4.000 205.720 245.600 206.400 ;
        RECT 4.400 205.000 245.600 205.720 ;
        RECT 4.400 204.320 246.000 205.000 ;
        RECT 4.000 200.960 246.000 204.320 ;
        RECT 4.000 199.600 245.600 200.960 ;
        RECT 4.400 199.560 245.600 199.600 ;
        RECT 4.400 198.200 246.000 199.560 ;
        RECT 4.000 195.520 246.000 198.200 ;
        RECT 4.000 194.120 245.600 195.520 ;
        RECT 4.000 193.480 246.000 194.120 ;
        RECT 4.400 192.080 246.000 193.480 ;
        RECT 4.000 190.080 246.000 192.080 ;
        RECT 4.000 188.680 245.600 190.080 ;
        RECT 4.000 187.360 246.000 188.680 ;
        RECT 4.400 185.960 246.000 187.360 ;
        RECT 4.000 184.640 246.000 185.960 ;
        RECT 4.000 183.240 245.600 184.640 ;
        RECT 4.000 181.240 246.000 183.240 ;
        RECT 4.400 179.840 246.000 181.240 ;
        RECT 4.000 179.200 246.000 179.840 ;
        RECT 4.000 177.800 245.600 179.200 ;
        RECT 4.000 175.120 246.000 177.800 ;
        RECT 4.400 173.760 246.000 175.120 ;
        RECT 4.400 173.720 245.600 173.760 ;
        RECT 4.000 172.360 245.600 173.720 ;
        RECT 4.000 169.000 246.000 172.360 ;
        RECT 4.400 168.320 246.000 169.000 ;
        RECT 4.400 167.600 245.600 168.320 ;
        RECT 4.000 166.920 245.600 167.600 ;
        RECT 4.000 162.880 246.000 166.920 ;
        RECT 4.400 161.480 245.600 162.880 ;
        RECT 4.000 157.440 246.000 161.480 ;
        RECT 4.000 156.760 245.600 157.440 ;
        RECT 4.400 156.040 245.600 156.760 ;
        RECT 4.400 155.360 246.000 156.040 ;
        RECT 4.000 152.000 246.000 155.360 ;
        RECT 4.000 150.640 245.600 152.000 ;
        RECT 4.400 150.600 245.600 150.640 ;
        RECT 4.400 149.240 246.000 150.600 ;
        RECT 4.000 146.560 246.000 149.240 ;
        RECT 4.000 145.160 245.600 146.560 ;
        RECT 4.000 144.520 246.000 145.160 ;
        RECT 4.400 143.120 246.000 144.520 ;
        RECT 4.000 141.120 246.000 143.120 ;
        RECT 4.000 139.720 245.600 141.120 ;
        RECT 4.000 138.400 246.000 139.720 ;
        RECT 4.400 137.000 246.000 138.400 ;
        RECT 4.000 135.680 246.000 137.000 ;
        RECT 4.000 134.280 245.600 135.680 ;
        RECT 4.000 132.280 246.000 134.280 ;
        RECT 4.400 130.880 246.000 132.280 ;
        RECT 4.000 130.240 246.000 130.880 ;
        RECT 4.000 128.840 245.600 130.240 ;
        RECT 4.000 126.160 246.000 128.840 ;
        RECT 4.400 124.800 246.000 126.160 ;
        RECT 4.400 124.760 245.600 124.800 ;
        RECT 4.000 123.400 245.600 124.760 ;
        RECT 4.000 120.040 246.000 123.400 ;
        RECT 4.400 119.360 246.000 120.040 ;
        RECT 4.400 118.640 245.600 119.360 ;
        RECT 4.000 117.960 245.600 118.640 ;
        RECT 4.000 113.920 246.000 117.960 ;
        RECT 4.400 112.520 245.600 113.920 ;
        RECT 4.000 108.480 246.000 112.520 ;
        RECT 4.000 107.800 245.600 108.480 ;
        RECT 4.400 107.080 245.600 107.800 ;
        RECT 4.400 106.400 246.000 107.080 ;
        RECT 4.000 103.040 246.000 106.400 ;
        RECT 4.000 101.680 245.600 103.040 ;
        RECT 4.400 101.640 245.600 101.680 ;
        RECT 4.400 100.280 246.000 101.640 ;
        RECT 4.000 97.600 246.000 100.280 ;
        RECT 4.000 96.200 245.600 97.600 ;
        RECT 4.000 95.560 246.000 96.200 ;
        RECT 4.400 94.160 246.000 95.560 ;
        RECT 4.000 92.160 246.000 94.160 ;
        RECT 4.000 90.760 245.600 92.160 ;
        RECT 4.000 89.440 246.000 90.760 ;
        RECT 4.400 88.040 246.000 89.440 ;
        RECT 4.000 86.720 246.000 88.040 ;
        RECT 4.000 85.320 245.600 86.720 ;
        RECT 4.000 83.320 246.000 85.320 ;
        RECT 4.400 81.920 246.000 83.320 ;
        RECT 4.000 81.280 246.000 81.920 ;
        RECT 4.000 79.880 245.600 81.280 ;
        RECT 4.000 77.200 246.000 79.880 ;
        RECT 4.400 75.840 246.000 77.200 ;
        RECT 4.400 75.800 245.600 75.840 ;
        RECT 4.000 74.440 245.600 75.800 ;
        RECT 4.000 71.080 246.000 74.440 ;
        RECT 4.400 70.400 246.000 71.080 ;
        RECT 4.400 69.680 245.600 70.400 ;
        RECT 4.000 69.000 245.600 69.680 ;
        RECT 4.000 64.960 246.000 69.000 ;
        RECT 4.400 63.560 245.600 64.960 ;
        RECT 4.000 59.520 246.000 63.560 ;
        RECT 4.000 58.840 245.600 59.520 ;
        RECT 4.400 58.120 245.600 58.840 ;
        RECT 4.400 57.440 246.000 58.120 ;
        RECT 4.000 54.080 246.000 57.440 ;
        RECT 4.000 52.720 245.600 54.080 ;
        RECT 4.400 52.680 245.600 52.720 ;
        RECT 4.400 51.320 246.000 52.680 ;
        RECT 4.000 48.640 246.000 51.320 ;
        RECT 4.000 47.240 245.600 48.640 ;
        RECT 4.000 46.600 246.000 47.240 ;
        RECT 4.400 45.200 246.000 46.600 ;
        RECT 4.000 43.200 246.000 45.200 ;
        RECT 4.000 41.800 245.600 43.200 ;
        RECT 4.000 40.480 246.000 41.800 ;
        RECT 4.400 39.080 246.000 40.480 ;
        RECT 4.000 37.760 246.000 39.080 ;
        RECT 4.000 36.360 245.600 37.760 ;
        RECT 4.000 34.360 246.000 36.360 ;
        RECT 4.400 32.960 246.000 34.360 ;
        RECT 4.000 32.320 246.000 32.960 ;
        RECT 4.000 30.920 245.600 32.320 ;
        RECT 4.000 28.240 246.000 30.920 ;
        RECT 4.400 26.880 246.000 28.240 ;
        RECT 4.400 26.840 245.600 26.880 ;
        RECT 4.000 25.480 245.600 26.840 ;
        RECT 4.000 22.120 246.000 25.480 ;
        RECT 4.400 21.440 246.000 22.120 ;
        RECT 4.400 20.720 245.600 21.440 ;
        RECT 4.000 20.040 245.600 20.720 ;
        RECT 4.000 16.000 246.000 20.040 ;
        RECT 4.400 14.600 245.600 16.000 ;
        RECT 4.000 9.880 246.000 14.600 ;
        RECT 4.400 9.015 246.000 9.880 ;
  END
END tiny_user_project
END LIBRARY

