VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 165.030 BY 175.750 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 12.280 165.030 12.880 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 114.280 165.030 114.880 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 124.480 165.030 125.080 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 134.680 165.030 135.280 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 144.880 165.030 145.480 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 155.080 165.030 155.680 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 171.750 160.450 175.750 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 171.750 142.510 175.750 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 171.750 124.570 175.750 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 171.750 106.630 175.750 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 171.750 88.690 175.750 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 22.480 165.030 23.080 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 171.750 70.750 175.750 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 171.750 52.810 175.750 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 171.750 34.870 175.750 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 171.750 16.930 175.750 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 32.680 165.030 33.280 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 42.880 165.030 43.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 53.080 165.030 53.680 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 63.280 165.030 63.880 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 73.480 165.030 74.080 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 83.680 165.030 84.280 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 93.880 165.030 94.480 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 104.080 165.030 104.680 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 19.080 165.030 19.680 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 121.080 165.030 121.680 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 131.280 165.030 131.880 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 141.480 165.030 142.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 151.680 165.030 152.280 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 161.880 165.030 162.480 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 171.750 148.490 175.750 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 171.750 130.550 175.750 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 171.750 112.610 175.750 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 171.750 94.670 175.750 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 171.750 76.730 175.750 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 29.280 165.030 29.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 171.750 58.790 175.750 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 171.750 40.850 175.750 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 171.750 22.910 175.750 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 171.750 4.970 175.750 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 39.480 165.030 40.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 49.680 165.030 50.280 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 59.880 165.030 60.480 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 70.080 165.030 70.680 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 80.280 165.030 80.880 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 90.480 165.030 91.080 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 100.680 165.030 101.280 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 110.880 165.030 111.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 15.680 165.030 16.280 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 117.680 165.030 118.280 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 127.880 165.030 128.480 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 138.080 165.030 138.680 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 148.280 165.030 148.880 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 158.480 165.030 159.080 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 171.750 154.470 175.750 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 171.750 136.530 175.750 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 171.750 118.590 175.750 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 171.750 100.650 175.750 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 171.750 82.710 175.750 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 25.880 165.030 26.480 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 171.750 64.770 175.750 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 171.750 46.830 175.750 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 171.750 28.890 175.750 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 171.750 10.950 175.750 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 36.080 165.030 36.680 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 46.280 165.030 46.880 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 56.480 165.030 57.080 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 66.680 165.030 67.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 76.880 165.030 77.480 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 87.080 165.030 87.680 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 97.280 165.030 97.880 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 161.030 107.480 165.030 108.080 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.925 10.640 25.525 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.335 10.640 63.935 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.745 10.640 102.345 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.155 10.640 140.755 163.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 43.130 10.640 44.730 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.540 10.640 83.140 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.950 10.640 121.550 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.360 10.640 159.960 163.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 159.160 163.285 ;
      LAYER met1 ;
        RECT 4.670 10.640 164.980 167.580 ;
      LAYER met2 ;
        RECT 5.250 171.470 10.390 174.605 ;
        RECT 11.230 171.470 16.370 174.605 ;
        RECT 17.210 171.470 22.350 174.605 ;
        RECT 23.190 171.470 28.330 174.605 ;
        RECT 29.170 171.470 34.310 174.605 ;
        RECT 35.150 171.470 40.290 174.605 ;
        RECT 41.130 171.470 46.270 174.605 ;
        RECT 47.110 171.470 52.250 174.605 ;
        RECT 53.090 171.470 58.230 174.605 ;
        RECT 59.070 171.470 64.210 174.605 ;
        RECT 65.050 171.470 70.190 174.605 ;
        RECT 71.030 171.470 76.170 174.605 ;
        RECT 77.010 171.470 82.150 174.605 ;
        RECT 82.990 171.470 88.130 174.605 ;
        RECT 88.970 171.470 94.110 174.605 ;
        RECT 94.950 171.470 100.090 174.605 ;
        RECT 100.930 171.470 106.070 174.605 ;
        RECT 106.910 171.470 112.050 174.605 ;
        RECT 112.890 171.470 118.030 174.605 ;
        RECT 118.870 171.470 124.010 174.605 ;
        RECT 124.850 171.470 129.990 174.605 ;
        RECT 130.830 171.470 135.970 174.605 ;
        RECT 136.810 171.470 141.950 174.605 ;
        RECT 142.790 171.470 147.930 174.605 ;
        RECT 148.770 171.470 153.910 174.605 ;
        RECT 154.750 171.470 159.890 174.605 ;
        RECT 160.730 171.470 164.980 174.605 ;
        RECT 4.700 3.555 164.980 171.470 ;
      LAYER met3 ;
        RECT 4.000 171.720 164.155 174.585 ;
        RECT 4.400 170.320 164.155 171.720 ;
        RECT 4.000 167.640 164.155 170.320 ;
        RECT 4.400 166.240 164.155 167.640 ;
        RECT 4.000 163.560 164.155 166.240 ;
        RECT 4.400 162.880 164.155 163.560 ;
        RECT 4.400 162.160 160.630 162.880 ;
        RECT 4.000 161.480 160.630 162.160 ;
        RECT 4.000 159.480 164.155 161.480 ;
        RECT 4.400 158.080 160.630 159.480 ;
        RECT 4.000 156.080 164.155 158.080 ;
        RECT 4.000 155.400 160.630 156.080 ;
        RECT 4.400 154.680 160.630 155.400 ;
        RECT 4.400 154.000 164.155 154.680 ;
        RECT 4.000 152.680 164.155 154.000 ;
        RECT 4.000 151.320 160.630 152.680 ;
        RECT 4.400 151.280 160.630 151.320 ;
        RECT 4.400 149.920 164.155 151.280 ;
        RECT 4.000 149.280 164.155 149.920 ;
        RECT 4.000 147.880 160.630 149.280 ;
        RECT 4.000 147.240 164.155 147.880 ;
        RECT 4.400 145.880 164.155 147.240 ;
        RECT 4.400 145.840 160.630 145.880 ;
        RECT 4.000 144.480 160.630 145.840 ;
        RECT 4.000 143.160 164.155 144.480 ;
        RECT 4.400 142.480 164.155 143.160 ;
        RECT 4.400 141.760 160.630 142.480 ;
        RECT 4.000 141.080 160.630 141.760 ;
        RECT 4.000 139.080 164.155 141.080 ;
        RECT 4.400 137.680 160.630 139.080 ;
        RECT 4.000 135.680 164.155 137.680 ;
        RECT 4.000 135.000 160.630 135.680 ;
        RECT 4.400 134.280 160.630 135.000 ;
        RECT 4.400 133.600 164.155 134.280 ;
        RECT 4.000 132.280 164.155 133.600 ;
        RECT 4.000 130.920 160.630 132.280 ;
        RECT 4.400 130.880 160.630 130.920 ;
        RECT 4.400 129.520 164.155 130.880 ;
        RECT 4.000 128.880 164.155 129.520 ;
        RECT 4.000 127.480 160.630 128.880 ;
        RECT 4.000 126.840 164.155 127.480 ;
        RECT 4.400 125.480 164.155 126.840 ;
        RECT 4.400 125.440 160.630 125.480 ;
        RECT 4.000 124.080 160.630 125.440 ;
        RECT 4.000 122.760 164.155 124.080 ;
        RECT 4.400 122.080 164.155 122.760 ;
        RECT 4.400 121.360 160.630 122.080 ;
        RECT 4.000 120.680 160.630 121.360 ;
        RECT 4.000 118.680 164.155 120.680 ;
        RECT 4.400 117.280 160.630 118.680 ;
        RECT 4.000 115.280 164.155 117.280 ;
        RECT 4.000 114.600 160.630 115.280 ;
        RECT 4.400 113.880 160.630 114.600 ;
        RECT 4.400 113.200 164.155 113.880 ;
        RECT 4.000 111.880 164.155 113.200 ;
        RECT 4.000 110.520 160.630 111.880 ;
        RECT 4.400 110.480 160.630 110.520 ;
        RECT 4.400 109.120 164.155 110.480 ;
        RECT 4.000 108.480 164.155 109.120 ;
        RECT 4.000 107.080 160.630 108.480 ;
        RECT 4.000 106.440 164.155 107.080 ;
        RECT 4.400 105.080 164.155 106.440 ;
        RECT 4.400 105.040 160.630 105.080 ;
        RECT 4.000 103.680 160.630 105.040 ;
        RECT 4.000 102.360 164.155 103.680 ;
        RECT 4.400 101.680 164.155 102.360 ;
        RECT 4.400 100.960 160.630 101.680 ;
        RECT 4.000 100.280 160.630 100.960 ;
        RECT 4.000 98.280 164.155 100.280 ;
        RECT 4.400 96.880 160.630 98.280 ;
        RECT 4.000 94.880 164.155 96.880 ;
        RECT 4.000 94.200 160.630 94.880 ;
        RECT 4.400 93.480 160.630 94.200 ;
        RECT 4.400 92.800 164.155 93.480 ;
        RECT 4.000 91.480 164.155 92.800 ;
        RECT 4.000 90.120 160.630 91.480 ;
        RECT 4.400 90.080 160.630 90.120 ;
        RECT 4.400 88.720 164.155 90.080 ;
        RECT 4.000 88.080 164.155 88.720 ;
        RECT 4.000 86.680 160.630 88.080 ;
        RECT 4.000 86.040 164.155 86.680 ;
        RECT 4.400 84.680 164.155 86.040 ;
        RECT 4.400 84.640 160.630 84.680 ;
        RECT 4.000 83.280 160.630 84.640 ;
        RECT 4.000 81.960 164.155 83.280 ;
        RECT 4.400 81.280 164.155 81.960 ;
        RECT 4.400 80.560 160.630 81.280 ;
        RECT 4.000 79.880 160.630 80.560 ;
        RECT 4.000 77.880 164.155 79.880 ;
        RECT 4.400 76.480 160.630 77.880 ;
        RECT 4.000 74.480 164.155 76.480 ;
        RECT 4.000 73.800 160.630 74.480 ;
        RECT 4.400 73.080 160.630 73.800 ;
        RECT 4.400 72.400 164.155 73.080 ;
        RECT 4.000 71.080 164.155 72.400 ;
        RECT 4.000 69.720 160.630 71.080 ;
        RECT 4.400 69.680 160.630 69.720 ;
        RECT 4.400 68.320 164.155 69.680 ;
        RECT 4.000 67.680 164.155 68.320 ;
        RECT 4.000 66.280 160.630 67.680 ;
        RECT 4.000 65.640 164.155 66.280 ;
        RECT 4.400 64.280 164.155 65.640 ;
        RECT 4.400 64.240 160.630 64.280 ;
        RECT 4.000 62.880 160.630 64.240 ;
        RECT 4.000 61.560 164.155 62.880 ;
        RECT 4.400 60.880 164.155 61.560 ;
        RECT 4.400 60.160 160.630 60.880 ;
        RECT 4.000 59.480 160.630 60.160 ;
        RECT 4.000 57.480 164.155 59.480 ;
        RECT 4.400 56.080 160.630 57.480 ;
        RECT 4.000 54.080 164.155 56.080 ;
        RECT 4.000 53.400 160.630 54.080 ;
        RECT 4.400 52.680 160.630 53.400 ;
        RECT 4.400 52.000 164.155 52.680 ;
        RECT 4.000 50.680 164.155 52.000 ;
        RECT 4.000 49.320 160.630 50.680 ;
        RECT 4.400 49.280 160.630 49.320 ;
        RECT 4.400 47.920 164.155 49.280 ;
        RECT 4.000 47.280 164.155 47.920 ;
        RECT 4.000 45.880 160.630 47.280 ;
        RECT 4.000 45.240 164.155 45.880 ;
        RECT 4.400 43.880 164.155 45.240 ;
        RECT 4.400 43.840 160.630 43.880 ;
        RECT 4.000 42.480 160.630 43.840 ;
        RECT 4.000 41.160 164.155 42.480 ;
        RECT 4.400 40.480 164.155 41.160 ;
        RECT 4.400 39.760 160.630 40.480 ;
        RECT 4.000 39.080 160.630 39.760 ;
        RECT 4.000 37.080 164.155 39.080 ;
        RECT 4.400 35.680 160.630 37.080 ;
        RECT 4.000 33.680 164.155 35.680 ;
        RECT 4.000 33.000 160.630 33.680 ;
        RECT 4.400 32.280 160.630 33.000 ;
        RECT 4.400 31.600 164.155 32.280 ;
        RECT 4.000 30.280 164.155 31.600 ;
        RECT 4.000 28.920 160.630 30.280 ;
        RECT 4.400 28.880 160.630 28.920 ;
        RECT 4.400 27.520 164.155 28.880 ;
        RECT 4.000 26.880 164.155 27.520 ;
        RECT 4.000 25.480 160.630 26.880 ;
        RECT 4.000 24.840 164.155 25.480 ;
        RECT 4.400 23.480 164.155 24.840 ;
        RECT 4.400 23.440 160.630 23.480 ;
        RECT 4.000 22.080 160.630 23.440 ;
        RECT 4.000 20.760 164.155 22.080 ;
        RECT 4.400 20.080 164.155 20.760 ;
        RECT 4.400 19.360 160.630 20.080 ;
        RECT 4.000 18.680 160.630 19.360 ;
        RECT 4.000 16.680 164.155 18.680 ;
        RECT 4.400 15.280 160.630 16.680 ;
        RECT 4.000 13.280 164.155 15.280 ;
        RECT 4.000 12.600 160.630 13.280 ;
        RECT 4.400 11.880 160.630 12.600 ;
        RECT 4.400 11.200 164.155 11.880 ;
        RECT 4.000 8.520 164.155 11.200 ;
        RECT 4.400 7.120 164.155 8.520 ;
        RECT 4.000 4.440 164.155 7.120 ;
        RECT 4.400 3.575 164.155 4.440 ;
      LAYER met4 ;
        RECT 26.975 163.840 163.465 174.585 ;
        RECT 26.975 23.295 42.730 163.840 ;
        RECT 45.130 23.295 61.935 163.840 ;
        RECT 64.335 23.295 81.140 163.840 ;
        RECT 83.540 23.295 100.345 163.840 ;
        RECT 102.745 23.295 119.550 163.840 ;
        RECT 121.950 23.295 138.755 163.840 ;
        RECT 141.155 23.295 157.960 163.840 ;
        RECT 160.360 23.295 163.465 163.840 ;
  END
END tiny_user_project
END LIBRARY

