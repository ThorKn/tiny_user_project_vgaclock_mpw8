// This is the unpowered netlist.
module tiny_user_project (io_in,
    io_oeb,
    io_out);
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire net17;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net18;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net19;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net55;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net56;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net57;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire \mod.thorkn_vgaclock.io_b ;
 wire \mod.thorkn_vgaclock.io_g ;
 wire \mod.thorkn_vgaclock.io_h_sync ;
 wire \mod.thorkn_vgaclock.io_r ;
 wire \mod.thorkn_vgaclock.io_v_sync ;
 wire \mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ;
 wire \mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ;
 wire \mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[0] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[10] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[11] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[12] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[13] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[14] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[15] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[16] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[17] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[18] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[19] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[20] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[21] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[22] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[23] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[24] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[4] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[5] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[6] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[7] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[8] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[9] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[0] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[11] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[12] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[13] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[14] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[15] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[17] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[18] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[19] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[21] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[22] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[24] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[4] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[5] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[6] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[7] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[8] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[9] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[0] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[0] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[4] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[5] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[0] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[1] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[2] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[3] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[4] ;
 wire \mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[5] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[0] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[1] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[2] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[3] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[4] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[5] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[6] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[7] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[8] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[9] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[8] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[0] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[1] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[2] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[3] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[4] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[5] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[6] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[7] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[8] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[9] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[2] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[3] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[5] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ;
 wire \mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;

 sky130_fd_sc_hd__clkinv_2 _0438_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[0] ));
 sky130_fd_sc_hd__and2_1 _0439_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ),
    .X(_0061_));
 sky130_fd_sc_hd__nor2_1 _0440_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ),
    .Y(_0062_));
 sky130_fd_sc_hd__nor2_1 _0441_ (.A(_0061_),
    .B(_0062_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[1] ));
 sky130_fd_sc_hd__and3_1 _0442_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ),
    .X(_0063_));
 sky130_fd_sc_hd__nor2_1 _0443_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ),
    .B(_0061_),
    .Y(_0064_));
 sky130_fd_sc_hd__nor2_1 _0444_ (.A(_0063_),
    .B(_0064_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[2] ));
 sky130_fd_sc_hd__and2_1 _0445_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .B(_0063_),
    .X(_0065_));
 sky130_fd_sc_hd__nor2_1 _0446_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .B(_0063_),
    .Y(_0066_));
 sky130_fd_sc_hd__nor2_1 _0447_ (.A(_0065_),
    .B(_0066_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[3] ));
 sky130_fd_sc_hd__and3_1 _0448_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .C(_0063_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2_1 _0449_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .B(_0065_),
    .Y(_0068_));
 sky130_fd_sc_hd__nor2_1 _0450_ (.A(_0067_),
    .B(_0068_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[4] ));
 sky130_fd_sc_hd__and2_1 _0451_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .B(_0067_),
    .X(_0069_));
 sky130_fd_sc_hd__buf_2 _0452_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[8] ),
    .X(_0070_));
 sky130_fd_sc_hd__or2_1 _0453_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ),
    .X(_0071_));
 sky130_fd_sc_hd__nor2_1 _0454_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ),
    .B(_0071_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand4_2 _0455_ (.A(_0070_),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .C(_0067_),
    .D(_0072_),
    .Y(_0073_));
 sky130_fd_sc_hd__o21ai_1 _0456_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .A2(_0067_),
    .B1(_0073_),
    .Y(_0074_));
 sky130_fd_sc_hd__nor2_1 _0457_ (.A(_0069_),
    .B(_0074_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[5] ));
 sky130_fd_sc_hd__and3_1 _0458_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_1 _0459_ (.A(_0065_),
    .B(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__o21a_1 _0460_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ),
    .A2(_0069_),
    .B1(_0076_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[6] ));
 sky130_fd_sc_hd__inv_2 _0461_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ),
    .Y(_0077_));
 sky130_fd_sc_hd__nor2_1 _0462_ (.A(_0077_),
    .B(_0076_),
    .Y(_0078_));
 sky130_fd_sc_hd__and2_1 _0463_ (.A(_0077_),
    .B(_0076_),
    .X(_0079_));
 sky130_fd_sc_hd__nor2_1 _0464_ (.A(_0078_),
    .B(_0079_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[7] ));
 sky130_fd_sc_hd__nand2_1 _0465_ (.A(_0070_),
    .B(_0078_),
    .Y(_0080_));
 sky130_fd_sc_hd__o211a_1 _0466_ (.A1(_0070_),
    .A2(_0078_),
    .B1(_0080_),
    .C1(_0073_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[8] ));
 sky130_fd_sc_hd__inv_2 _0467_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .Y(_0081_));
 sky130_fd_sc_hd__and4_1 _0468_ (.A(_0070_),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .C(_0067_),
    .D(_0072_),
    .X(_0082_));
 sky130_fd_sc_hd__a31o_1 _0469_ (.A1(_0070_),
    .A2(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .A3(_0078_),
    .B1(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__a21oi_1 _0470_ (.A1(_0081_),
    .A2(_0080_),
    .B1(_0083_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[9] ));
 sky130_fd_sc_hd__xnor2_1 _0471_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .B(_0073_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[0] ));
 sky130_fd_sc_hd__a21oi_1 _0472_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .A2(_0082_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .Y(_0084_));
 sky130_fd_sc_hd__and3_1 _0473_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .C(_0082_),
    .X(_0085_));
 sky130_fd_sc_hd__nor2_1 _0474_ (.A(_0084_),
    .B(_0085_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[1] ));
 sky130_fd_sc_hd__clkbuf_2 _0475_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[2] ),
    .X(_0086_));
 sky130_fd_sc_hd__inv_2 _0476_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[2] ),
    .Y(_0087_));
 sky130_fd_sc_hd__and2_1 _0477_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .X(_0088_));
 sky130_fd_sc_hd__or3b_1 _0478_ (.A(_0087_),
    .B(_0073_),
    .C_N(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__buf_2 _0479_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[5] ),
    .X(_0090_));
 sky130_fd_sc_hd__or3_2 _0480_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ),
    .X(_0091_));
 sky130_fd_sc_hd__or2_1 _0481_ (.A(_0090_),
    .B(_0091_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_2 _0482_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[3] ),
    .X(_0093_));
 sky130_fd_sc_hd__and4_1 _0483_ (.A(_0087_),
    .B(_0093_),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ),
    .D(_0088_),
    .X(_0094_));
 sky130_fd_sc_hd__or4b_1 _0484_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .B(_0073_),
    .C(_0092_),
    .D_N(_0094_),
    .X(_0095_));
 sky130_fd_sc_hd__o211a_1 _0485_ (.A1(_0086_),
    .A2(_0085_),
    .B1(_0089_),
    .C1(_0095_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[2] ));
 sky130_fd_sc_hd__a31o_1 _0486_ (.A1(_0086_),
    .A2(_0082_),
    .A3(_0088_),
    .B1(_0093_),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _0487_ (.A(_0086_),
    .B(_0093_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _0488_ (.A(_0085_),
    .B(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__clkinv_2 _0489_ (.A(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__and3_1 _0490_ (.A(_0095_),
    .B(_0096_),
    .C(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0491_ (.A(_0100_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[3] ));
 sky130_fd_sc_hd__xor2_1 _0492_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .B(_0098_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[4] ));
 sky130_fd_sc_hd__a21oi_1 _0493_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .A2(_0098_),
    .B1(_0090_),
    .Y(_0101_));
 sky130_fd_sc_hd__and3_1 _0494_ (.A(_0090_),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .C(_0098_),
    .X(_0102_));
 sky130_fd_sc_hd__nor2_1 _0495_ (.A(_0101_),
    .B(_0102_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[5] ));
 sky130_fd_sc_hd__xor2_1 _0496_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .B(_0102_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[6] ));
 sky130_fd_sc_hd__a21oi_1 _0497_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .A2(_0102_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ),
    .Y(_0103_));
 sky130_fd_sc_hd__and3_1 _0498_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .C(_0102_),
    .X(_0104_));
 sky130_fd_sc_hd__nor2_1 _0499_ (.A(_0103_),
    .B(_0104_),
    .Y(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[7] ));
 sky130_fd_sc_hd__xor2_1 _0500_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ),
    .B(_0104_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[8] ));
 sky130_fd_sc_hd__a21o_1 _0501_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ),
    .A2(_0104_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ),
    .X(_0105_));
 sky130_fd_sc_hd__nand3_1 _0502_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ),
    .C(_0104_),
    .Y(_0106_));
 sky130_fd_sc_hd__and3_1 _0503_ (.A(_0095_),
    .B(_0105_),
    .C(_0106_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0504_ (.A(_0107_),
    .X(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[9] ));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ),
    .Y(_0108_));
 sky130_fd_sc_hd__and4b_1 _0506_ (.A_N(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .D(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_1 _0507_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ),
    .Y(_0110_));
 sky130_fd_sc_hd__and4b_1 _0508_ (.A_N(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .C(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .X(_0111_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__and4_1 _0510_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[0] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[3] ),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[2] ),
    .X(_0113_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0511_ (.A(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__nand3_1 _0512_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[4] ),
    .C(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__nand4_1 _0513_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[19] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[21] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[22] ),
    .Y(_0116_));
 sky130_fd_sc_hd__or4bb_1 _0514_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[15] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[17] ),
    .C_N(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[24] ),
    .D_N(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[14] ),
    .X(_0117_));
 sky130_fd_sc_hd__or4bb_1 _0515_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ),
    .B(_0117_),
    .C_N(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ),
    .D_N(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[18] ),
    .X(_0118_));
 sky130_fd_sc_hd__or3_1 _0516_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[7] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[6] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[9] ),
    .X(_0119_));
 sky130_fd_sc_hd__and4b_1 _0517_ (.A_N(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[11] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[13] ),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[12] ),
    .X(_0120_));
 sky130_fd_sc_hd__or3b_1 _0518_ (.A(_0119_),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[8] ),
    .C_N(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__or4_1 _0519_ (.A(_0115_),
    .B(_0116_),
    .C(_0118_),
    .D(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__nor3_1 _0520_ (.A(_0110_),
    .B(_0112_),
    .C(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__and4_1 _0521_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .C(_0109_),
    .D(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__xnor2_1 _0522_ (.A(_0108_),
    .B(_0124_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[0] ));
 sky130_fd_sc_hd__a21oi_1 _0523_ (.A1(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ),
    .A2(_0124_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ),
    .Y(_0125_));
 sky130_fd_sc_hd__and3_1 _0524_ (.A(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ),
    .C(_0124_),
    .X(_0126_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0525_ (.A(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__nor2_1 _0526_ (.A(_0125_),
    .B(_0127_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[1] ));
 sky130_fd_sc_hd__inv_2 _0527_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .Y(_0128_));
 sky130_fd_sc_hd__a21oi_1 _0528_ (.A1(_0128_),
    .A2(_0127_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ),
    .Y(_0129_));
 sky130_fd_sc_hd__a21oi_1 _0529_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ),
    .A2(_0127_),
    .B1(_0129_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[2] ));
 sky130_fd_sc_hd__a21oi_1 _0530_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ),
    .A2(_0127_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .Y(_0130_));
 sky130_fd_sc_hd__a21oi_1 _0531_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .A2(_0127_),
    .B1(_0130_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[3] ));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .Y(_0131_));
 sky130_fd_sc_hd__xnor2_1 _0533_ (.A(_0131_),
    .B(_0123_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[0] ));
 sky130_fd_sc_hd__a21oi_1 _0534_ (.A1(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .A2(_0123_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_1 _0535_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .B(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .Y(_0133_));
 sky130_fd_sc_hd__or3b_1 _0536_ (.A(_0119_),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[8] ),
    .C_N(_0120_),
    .X(_0134_));
 sky130_fd_sc_hd__or4_1 _0537_ (.A(_0115_),
    .B(_0116_),
    .C(_0118_),
    .D(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_2 _0538_ (.A(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__or3_1 _0539_ (.A(_0110_),
    .B(_0112_),
    .C(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__nor2_1 _0540_ (.A(_0133_),
    .B(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__nor2_1 _0541_ (.A(_0132_),
    .B(_0138_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[1] ));
 sky130_fd_sc_hd__nor3_1 _0542_ (.A(_0110_),
    .B(_0112_),
    .C(_0135_),
    .Y(_0139_));
 sky130_fd_sc_hd__nand4_1 _0543_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .C(_0109_),
    .D(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__or2_1 _0544_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ),
    .B(_0138_),
    .X(_0141_));
 sky130_fd_sc_hd__and4_1 _0545_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .B(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ),
    .D(_0139_),
    .X(_0142_));
 sky130_fd_sc_hd__inv_2 _0546_ (.A(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__and3_1 _0547_ (.A(_0140_),
    .B(_0141_),
    .C(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0548_ (.A(_0144_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[2] ));
 sky130_fd_sc_hd__or2_1 _0549_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .B(_0142_),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_1 _0550_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .B(_0142_),
    .Y(_0146_));
 sky130_fd_sc_hd__and3_1 _0551_ (.A(_0140_),
    .B(_0145_),
    .C(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _0552_ (.A(_0147_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[3] ));
 sky130_fd_sc_hd__xor2_1 _0553_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .X(_0148_));
 sky130_fd_sc_hd__or2_1 _0554_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .B(_0142_),
    .X(_0149_));
 sky130_fd_sc_hd__o211a_1 _0555_ (.A1(_0143_),
    .A2(_0148_),
    .B1(_0149_),
    .C1(_0140_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[4] ));
 sky130_fd_sc_hd__xor2_2 _0556_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .X(_0150_));
 sky130_fd_sc_hd__a21o_1 _0557_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .A2(_0142_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ),
    .X(_0151_));
 sky130_fd_sc_hd__o211a_1 _0558_ (.A1(_0146_),
    .A2(_0150_),
    .B1(_0151_),
    .C1(_0140_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[5] ));
 sky130_fd_sc_hd__clkinv_2 _0559_ (.A(_0135_),
    .Y(_0152_));
 sky130_fd_sc_hd__nor2_1 _0560_ (.A(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__nand2_1 _0561_ (.A(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .B(_0152_),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _0562_ (.A(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor2_1 _0563_ (.A(_0153_),
    .B(_0155_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[0] ));
 sky130_fd_sc_hd__nand2_1 _0564_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .B(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .Y(_0156_));
 sky130_fd_sc_hd__o22a_1 _0565_ (.A1(_0156_),
    .A2(_0136_),
    .B1(_0155_),
    .B2(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[1] ));
 sky130_fd_sc_hd__a31o_1 _0566_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .A2(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .A3(_0152_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ),
    .X(_0157_));
 sky130_fd_sc_hd__and4_1 _0567_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .B(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ),
    .D(_0152_),
    .X(_0158_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__and3_1 _0569_ (.A(_0137_),
    .B(_0157_),
    .C(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _0570_ (.A(_0160_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[2] ));
 sky130_fd_sc_hd__or2_1 _0571_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .B(_0158_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _0572_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .B(_0158_),
    .Y(_0162_));
 sky130_fd_sc_hd__and3_1 _0573_ (.A(_0137_),
    .B(_0161_),
    .C(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_1 _0574_ (.A(_0163_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[3] ));
 sky130_fd_sc_hd__xor2_1 _0575_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ),
    .X(_0164_));
 sky130_fd_sc_hd__or2_1 _0576_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ),
    .B(_0158_),
    .X(_0165_));
 sky130_fd_sc_hd__o211a_1 _0577_ (.A1(_0159_),
    .A2(_0164_),
    .B1(_0165_),
    .C1(_0137_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[4] ));
 sky130_fd_sc_hd__or2_1 _0578_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _0579_ (.A(_0110_),
    .B(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__inv_2 _0580_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2_1 _0581_ (.A(_0168_),
    .B(_0162_),
    .Y(_0169_));
 sky130_fd_sc_hd__o211a_1 _0582_ (.A1(_0162_),
    .A2(_0167_),
    .B1(_0169_),
    .C1(_0137_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[5] ));
 sky130_fd_sc_hd__clkinv_2 _0583_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[0] ),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[0] ));
 sky130_fd_sc_hd__xor2_1 _0584_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[0] ),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[1] ));
 sky130_fd_sc_hd__and3_1 _0585_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[0] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[2] ),
    .X(_0170_));
 sky130_fd_sc_hd__a21oi_1 _0586_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[1] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[0] ),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[2] ),
    .Y(_0171_));
 sky130_fd_sc_hd__nor2_1 _0587_ (.A(_0170_),
    .B(_0171_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[2] ));
 sky130_fd_sc_hd__nor2_1 _0588_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[3] ),
    .B(_0170_),
    .Y(_0172_));
 sky130_fd_sc_hd__nor2_1 _0589_ (.A(_0114_),
    .B(_0172_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[3] ));
 sky130_fd_sc_hd__xor2_1 _0590_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[4] ),
    .B(_0114_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[4] ));
 sky130_fd_sc_hd__and3_1 _0591_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[4] ),
    .C(_0114_),
    .X(_0173_));
 sky130_fd_sc_hd__a21oi_1 _0592_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[4] ),
    .A2(_0114_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[5] ),
    .Y(_0174_));
 sky130_fd_sc_hd__nor2_1 _0593_ (.A(_0173_),
    .B(_0174_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[5] ));
 sky130_fd_sc_hd__nor2_1 _0594_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[6] ),
    .B(_0173_),
    .Y(_0175_));
 sky130_fd_sc_hd__and4_1 _0595_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[5] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[4] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[6] ),
    .D(_0114_),
    .X(_0176_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0596_ (.A(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__nor3_1 _0597_ (.A(_0152_),
    .B(_0175_),
    .C(_0177_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[6] ));
 sky130_fd_sc_hd__xor2_1 _0598_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[7] ),
    .B(_0177_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[7] ));
 sky130_fd_sc_hd__nand2_1 _0599_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[7] ),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__xnor2_1 _0600_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[8] ),
    .B(_0178_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[8] ));
 sky130_fd_sc_hd__and4_1 _0601_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[7] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[9] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[8] ),
    .D(_0177_),
    .X(_0179_));
 sky130_fd_sc_hd__a31o_1 _0602_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[7] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[8] ),
    .A3(_0177_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[9] ),
    .X(_0180_));
 sky130_fd_sc_hd__and2b_1 _0603_ (.A_N(_0179_),
    .B(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _0604_ (.A(_0181_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[9] ));
 sky130_fd_sc_hd__xor2_1 _0605_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ),
    .B(_0179_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[10] ));
 sky130_fd_sc_hd__a21o_1 _0606_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ),
    .A2(_0179_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[11] ),
    .X(_0182_));
 sky130_fd_sc_hd__nand3_1 _0607_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[11] ),
    .C(_0179_),
    .Y(_0183_));
 sky130_fd_sc_hd__and3_1 _0608_ (.A(_0136_),
    .B(_0182_),
    .C(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0609_ (.A(_0184_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[11] ));
 sky130_fd_sc_hd__inv_2 _0610_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[12] ),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_1 _0611_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[11] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[12] ),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _0612_ (.A(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__and3_1 _0613_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ),
    .B(_0187_),
    .C(_0179_),
    .X(_0188_));
 sky130_fd_sc_hd__a211oi_1 _0614_ (.A1(_0185_),
    .A2(_0183_),
    .B1(_0188_),
    .C1(_0152_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[12] ));
 sky130_fd_sc_hd__and4_1 _0615_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[13] ),
    .C(_0187_),
    .D(_0179_),
    .X(_0189_));
 sky130_fd_sc_hd__inv_2 _0616_ (.A(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__o211a_1 _0617_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[13] ),
    .A2(_0188_),
    .B1(_0190_),
    .C1(_0136_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[13] ));
 sky130_fd_sc_hd__nand2_1 _0618_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[14] ),
    .B(_0189_),
    .Y(_0191_));
 sky130_fd_sc_hd__o211a_1 _0619_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[14] ),
    .A2(_0189_),
    .B1(_0191_),
    .C1(_0136_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[14] ));
 sky130_fd_sc_hd__a21oi_1 _0620_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[14] ),
    .A2(_0189_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[15] ),
    .Y(_0192_));
 sky130_fd_sc_hd__and3_1 _0621_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[15] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[14] ),
    .C(_0189_),
    .X(_0193_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0622_ (.A(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__nor2_1 _0623_ (.A(_0192_),
    .B(_0194_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[15] ));
 sky130_fd_sc_hd__nor2_1 _0624_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__a211oi_1 _0625_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ),
    .A2(_0194_),
    .B1(_0195_),
    .C1(_0152_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[16] ));
 sky130_fd_sc_hd__a21oi_1 _0626_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ),
    .A2(_0194_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[17] ),
    .Y(_0196_));
 sky130_fd_sc_hd__and3_1 _0627_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[17] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ),
    .C(_0194_),
    .X(_0197_));
 sky130_fd_sc_hd__nor2_1 _0628_ (.A(_0196_),
    .B(_0197_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[17] ));
 sky130_fd_sc_hd__or2_1 _0629_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[18] ),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__and4_1 _0630_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[17] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[18] ),
    .D(_0194_),
    .X(_0199_));
 sky130_fd_sc_hd__inv_2 _0631_ (.A(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__and3_1 _0632_ (.A(_0136_),
    .B(_0198_),
    .C(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _0633_ (.A(_0201_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[18] ));
 sky130_fd_sc_hd__and2_1 _0634_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[19] ),
    .B(_0199_),
    .X(_0202_));
 sky130_fd_sc_hd__inv_2 _0635_ (.A(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__o211a_1 _0636_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[19] ),
    .A2(_0199_),
    .B1(_0203_),
    .C1(_0136_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[19] ));
 sky130_fd_sc_hd__nand2_1 _0637_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ),
    .B(_0202_),
    .Y(_0204_));
 sky130_fd_sc_hd__o211a_1 _0638_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ),
    .A2(_0202_),
    .B1(_0204_),
    .C1(_0136_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[20] ));
 sky130_fd_sc_hd__a31o_1 _0639_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[19] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ),
    .A3(_0199_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[21] ),
    .X(_0205_));
 sky130_fd_sc_hd__nand3_1 _0640_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[21] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ),
    .C(_0202_),
    .Y(_0206_));
 sky130_fd_sc_hd__and3_1 _0641_ (.A(_0136_),
    .B(_0205_),
    .C(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _0642_ (.A(_0207_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[21] ));
 sky130_fd_sc_hd__a31o_1 _0643_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[21] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ),
    .A3(_0202_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[22] ),
    .X(_0208_));
 sky130_fd_sc_hd__o211a_1 _0644_ (.A1(_0116_),
    .A2(_0200_),
    .B1(_0208_),
    .C1(_0136_),
    .X(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[22] ));
 sky130_fd_sc_hd__and4_1 _0645_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[19] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[21] ),
    .C(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[22] ),
    .X(_0209_));
 sky130_fd_sc_hd__a21oi_1 _0646_ (.A1(_0209_),
    .A2(_0199_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ),
    .Y(_0210_));
 sky130_fd_sc_hd__and3_1 _0647_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ),
    .B(_0209_),
    .C(_0199_),
    .X(_0211_));
 sky130_fd_sc_hd__nor2_1 _0648_ (.A(_0210_),
    .B(_0211_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[23] ));
 sky130_fd_sc_hd__nor2_1 _0649_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[24] ),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__a211oi_1 _0650_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[24] ),
    .A2(_0211_),
    .B1(_0212_),
    .C1(_0152_),
    .Y(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[24] ));
 sky130_fd_sc_hd__or2_1 _0651_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ),
    .X(_0213_));
 sky130_fd_sc_hd__or3_1 _0652_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ),
    .C(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__a2bb2o_1 _0653_ (.A1_N(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .A2_N(_0071_),
    .B1(_0075_),
    .B2(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__or4_1 _0654_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ),
    .B(_0070_),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .D(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _0655_ (.A(_0216_),
    .X(\mod.thorkn_vgaclock.io_h_sync ));
 sky130_fd_sc_hd__nand2_1 _0656_ (.A(_0093_),
    .B(_0088_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _0657_ (.A(_0086_),
    .B(_0093_),
    .Y(_0218_));
 sky130_fd_sc_hd__o22a_1 _0658_ (.A1(_0086_),
    .A2(_0217_),
    .B1(_0218_),
    .B2(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .X(_0219_));
 sky130_fd_sc_hd__or4_1 _0659_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ),
    .C(_0092_),
    .D(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0220_),
    .X(\mod.thorkn_vgaclock.io_v_sync ));
 sky130_fd_sc_hd__inv_2 _0661_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .Y(_0221_));
 sky130_fd_sc_hd__a21o_2 _0662_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[2] ),
    .A2(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[3] ),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .X(_0222_));
 sky130_fd_sc_hd__a211o_1 _0663_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[5] ),
    .A2(_0222_),
    .B1(_0091_),
    .C1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ),
    .X(_0223_));
 sky130_fd_sc_hd__clkbuf_2 _0664_ (.A(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__o21a_2 _0665_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .A2(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ),
    .X(_0225_));
 sky130_fd_sc_hd__or3_1 _0666_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[8] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .C(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_2 _0667_ (.A(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__o211a_1 _0668_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .A2(_0221_),
    .B1(_0224_),
    .C1(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_1 _0669_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ),
    .Y(_0229_));
 sky130_fd_sc_hd__a211oi_4 _0670_ (.A1(_0090_),
    .A2(_0222_),
    .B1(_0091_),
    .C1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ),
    .Y(_0230_));
 sky130_fd_sc_hd__nor3_4 _0671_ (.A(_0070_),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .C(_0225_),
    .Y(_0231_));
 sky130_fd_sc_hd__a211oi_1 _0672_ (.A1(_0071_),
    .A2(_0229_),
    .B1(_0230_),
    .C1(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__o211a_1 _0673_ (.A1(_0213_),
    .A2(_0228_),
    .B1(_0232_),
    .C1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .X(_0233_));
 sky130_fd_sc_hd__o211a_1 _0674_ (.A1(_0070_),
    .A2(_0225_),
    .B1(_0224_),
    .C1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ),
    .X(_0234_));
 sky130_fd_sc_hd__xnor2_1 _0675_ (.A(_0070_),
    .B(_0225_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _0676_ (.A(_0223_),
    .B(_0226_),
    .Y(_0236_));
 sky130_fd_sc_hd__clkbuf_2 _0677_ (.A(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__nor3_1 _0678_ (.A(_0072_),
    .B(_0225_),
    .C(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__or2_1 _0679_ (.A(_0235_),
    .B(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0680_ (.A0(_0233_),
    .A1(_0234_),
    .S(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__nor2_2 _0681_ (.A(_0230_),
    .B(_0231_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand3_1 _0682_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ),
    .C(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__nor2_1 _0683_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__a21o_1 _0684_ (.A1(_0241_),
    .A2(_0235_),
    .B1(_0234_),
    .X(_0244_));
 sky130_fd_sc_hd__a311oi_2 _0685_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ),
    .A2(_0071_),
    .A3(_0229_),
    .B1(_0230_),
    .C1(_0231_),
    .Y(_0245_));
 sky130_fd_sc_hd__a211oi_1 _0686_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .A2(_0243_),
    .B1(_0244_),
    .C1(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__a211o_1 _0687_ (.A1(_0090_),
    .A2(_0222_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .C1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ),
    .X(_0247_));
 sky130_fd_sc_hd__xor2_1 _0688_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ),
    .B(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_1 _0689_ (.A(_0237_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__and2_1 _0690_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ),
    .B(_0227_),
    .X(_0250_));
 sky130_fd_sc_hd__o21a_1 _0691_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ),
    .A2(_0247_),
    .B1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__a21oi_2 _0692_ (.A1(_0090_),
    .A2(_0222_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .Y(_0252_));
 sky130_fd_sc_hd__xnor2_2 _0693_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__or2_1 _0694_ (.A(_0237_),
    .B(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _0695_ (.A(_0090_),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .C(_0222_),
    .X(_0255_));
 sky130_fd_sc_hd__or2_1 _0696_ (.A(_0252_),
    .B(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__or2_1 _0697_ (.A(_0086_),
    .B(_0093_),
    .X(_0257_));
 sky130_fd_sc_hd__and4_1 _0698_ (.A(_0218_),
    .B(_0224_),
    .C(_0227_),
    .D(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__nand4_1 _0699_ (.A(_0086_),
    .B(_0253_),
    .C(_0256_),
    .D(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__o31a_1 _0700_ (.A1(_0254_),
    .A2(_0256_),
    .A3(_0257_),
    .B1(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .Y(_0261_));
 sky130_fd_sc_hd__a21oi_1 _0702_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[2] ),
    .A2(_0093_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .Y(_0262_));
 sky130_fd_sc_hd__and3_1 _0703_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[2] ),
    .B(_0093_),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _0704_ (.A(_0262_),
    .B(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__or3b_2 _0705_ (.A(_0230_),
    .B(_0231_),
    .C_N(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__xnor2_1 _0706_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[5] ),
    .B(_0262_),
    .Y(_0266_));
 sky130_fd_sc_hd__and3_1 _0707_ (.A(_0223_),
    .B(_0226_),
    .C(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__clkbuf_2 _0708_ (.A(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__o41a_1 _0709_ (.A1(_0236_),
    .A2(_0253_),
    .A3(_0256_),
    .A4(_0257_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .X(_0269_));
 sky130_fd_sc_hd__and4_1 _0710_ (.A(_0223_),
    .B(_0226_),
    .C(_0266_),
    .D(_0264_),
    .X(_0270_));
 sky130_fd_sc_hd__or3b_1 _0711_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .C_N(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__o41a_1 _0712_ (.A1(_0261_),
    .A2(_0265_),
    .A3(_0268_),
    .A4(_0269_),
    .B1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__or3_1 _0713_ (.A(_0261_),
    .B(_0230_),
    .C(_0231_),
    .X(_0273_));
 sky130_fd_sc_hd__nand2_1 _0714_ (.A(_0270_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor2_1 _0715_ (.A(_0237_),
    .B(_0253_),
    .Y(_0275_));
 sky130_fd_sc_hd__o211a_1 _0716_ (.A1(_0252_),
    .A2(_0255_),
    .B1(_0227_),
    .C1(_0224_),
    .X(_0276_));
 sky130_fd_sc_hd__and3_1 _0717_ (.A(_0087_),
    .B(_0223_),
    .C(_0226_),
    .X(_0277_));
 sky130_fd_sc_hd__and2_1 _0718_ (.A(_0093_),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__or3b_1 _0719_ (.A(_0275_),
    .B(_0276_),
    .C_N(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__and3_1 _0720_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .B(_0223_),
    .C(_0226_),
    .X(_0280_));
 sky130_fd_sc_hd__and4b_1 _0721_ (.A_N(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .B(_0090_),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ),
    .X(_0281_));
 sky130_fd_sc_hd__and3_1 _0722_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ),
    .B(_0280_),
    .C(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__and4b_1 _0723_ (.A_N(_0253_),
    .B(_0270_),
    .C(_0273_),
    .D(_0276_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _0724_ (.A(_0218_),
    .B(_0241_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _0725_ (.A1(_0282_),
    .A2(_0283_),
    .B1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__o221a_1 _0726_ (.A1(_0260_),
    .A2(_0272_),
    .B1(_0274_),
    .B2(_0279_),
    .C1(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__or2_1 _0727_ (.A(_0237_),
    .B(_0248_),
    .X(_0287_));
 sky130_fd_sc_hd__a2111o_1 _0728_ (.A1(_0261_),
    .A2(_0090_),
    .B1(_0264_),
    .C1(_0287_),
    .D1(_0251_),
    .X(_0288_));
 sky130_fd_sc_hd__a221o_1 _0729_ (.A1(_0088_),
    .A2(_0259_),
    .B1(_0260_),
    .B2(_0279_),
    .C1(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__o21ba_1 _0730_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .A2(_0269_),
    .B1_N(_0090_),
    .X(_0290_));
 sky130_fd_sc_hd__o32a_1 _0731_ (.A1(_0249_),
    .A2(_0251_),
    .A3(_0286_),
    .B1(_0289_),
    .B2(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__nor3_1 _0732_ (.A(_0240_),
    .B(_0246_),
    .C(_0291_),
    .Y(\mod.thorkn_vgaclock.io_r ));
 sky130_fd_sc_hd__or3_1 _0733_ (.A(_0072_),
    .B(_0225_),
    .C(_0237_),
    .X(_0292_));
 sky130_fd_sc_hd__xor2_1 _0734_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .A1(_0133_),
    .S(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__xor2_1 _0736_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .X(_0295_));
 sky130_fd_sc_hd__o21ai_1 _0737_ (.A1(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .Y(_0296_));
 sky130_fd_sc_hd__xnor2_1 _0738_ (.A(_0295_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21a_1 _0739_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_2 _0740_ (.A1(_0109_),
    .A2(_0298_),
    .B1(_0148_),
    .Y(_0299_));
 sky130_fd_sc_hd__or3_1 _0741_ (.A(_0109_),
    .B(_0148_),
    .C(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__o211a_1 _0742_ (.A1(_0294_),
    .A2(_0297_),
    .B1(_0299_),
    .C1(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__nand2_1 _0743_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .Y(_0302_));
 sky130_fd_sc_hd__and3_1 _0744_ (.A(_0302_),
    .B(_0150_),
    .C(_0299_),
    .X(_0303_));
 sky130_fd_sc_hd__a21oi_1 _0745_ (.A1(_0302_),
    .A2(_0299_),
    .B1(_0150_),
    .Y(_0304_));
 sky130_fd_sc_hd__or2_1 _0746_ (.A(_0303_),
    .B(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__xnor2_1 _0747_ (.A(_0301_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(_0268_),
    .Y(_0307_));
 sky130_fd_sc_hd__a211oi_1 _0749_ (.A1(_0299_),
    .A2(_0300_),
    .B1(_0294_),
    .C1(_0297_),
    .Y(_0308_));
 sky130_fd_sc_hd__nor3_1 _0750_ (.A(_0307_),
    .B(_0301_),
    .C(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__and4_1 _0751_ (.A(_0087_),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .C(_0224_),
    .D(_0227_),
    .X(_0310_));
 sky130_fd_sc_hd__xnor2_1 _0752_ (.A(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ),
    .B(_0293_),
    .Y(_0311_));
 sky130_fd_sc_hd__a41o_1 _0753_ (.A1(_0218_),
    .A2(_0224_),
    .A3(_0227_),
    .A4(_0257_),
    .B1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a31o_1 _0754_ (.A1(_0087_),
    .A2(_0224_),
    .A3(_0227_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ),
    .X(_0313_));
 sky130_fd_sc_hd__o311a_1 _0755_ (.A1(_0131_),
    .A2(_0280_),
    .A3(_0310_),
    .B1(_0312_),
    .C1(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__xor2_1 _0756_ (.A(_0294_),
    .B(_0297_),
    .X(_0315_));
 sky130_fd_sc_hd__a2bb2o_1 _0757_ (.A1_N(_0315_),
    .A2_N(_0265_),
    .B1(_0258_),
    .B2(_0311_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_1 _0758_ (.A(_0265_),
    .B(_0315_),
    .Y(_0317_));
 sky130_fd_sc_hd__o21bai_1 _0759_ (.A1(_0301_),
    .A2(_0308_),
    .B1_N(_0268_),
    .Y(_0318_));
 sky130_fd_sc_hd__o211a_1 _0760_ (.A1(_0314_),
    .A2(_0316_),
    .B1(_0317_),
    .C1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a211o_1 _0761_ (.A1(_0276_),
    .A2(_0306_),
    .B1(_0309_),
    .C1(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__or2_1 _0762_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .B(_0299_),
    .X(_0321_));
 sky130_fd_sc_hd__or3b_1 _0763_ (.A(_0298_),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ),
    .C_N(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .X(_0322_));
 sky130_fd_sc_hd__a311o_1 _0764_ (.A1(_0150_),
    .A2(_0321_),
    .A3(_0322_),
    .B1(_0303_),
    .C1(_0304_),
    .X(_0323_));
 sky130_fd_sc_hd__o211a_1 _0765_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ),
    .A2(_0299_),
    .B1(_0322_),
    .C1(_0150_),
    .X(_0324_));
 sky130_fd_sc_hd__o31a_1 _0766_ (.A1(_0301_),
    .A2(_0303_),
    .A3(_0304_),
    .B1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__o21bai_1 _0767_ (.A1(_0301_),
    .A2(_0323_),
    .B1_N(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__o2bb2a_1 _0768_ (.A1_N(_0254_),
    .A2_N(_0326_),
    .B1(_0306_),
    .B2(_0276_),
    .X(_0327_));
 sky130_fd_sc_hd__o21ai_1 _0769_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ),
    .A2(_0325_),
    .B1(_0249_),
    .Y(_0328_));
 sky130_fd_sc_hd__o21ai_1 _0770_ (.A1(_0254_),
    .A2(_0326_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a211o_1 _0771_ (.A1(_0320_),
    .A2(_0327_),
    .B1(_0329_),
    .C1(_0251_),
    .X(_0330_));
 sky130_fd_sc_hd__o2111a_1 _0772_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ),
    .A2(_0241_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .C1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ),
    .D1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ),
    .X(_0331_));
 sky130_fd_sc_hd__or3_1 _0773_ (.A(_0228_),
    .B(_0245_),
    .C(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__and3_1 _0774_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .B(_0221_),
    .C(_0232_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _0775_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ),
    .A2(_0213_),
    .B1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__and3b_1 _0776_ (.A_N(_0234_),
    .B(_0235_),
    .C(_0241_),
    .X(_0335_));
 sky130_fd_sc_hd__or3_1 _0777_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ),
    .B(_0249_),
    .C(_0325_),
    .X(_0336_));
 sky130_fd_sc_hd__and4_1 _0778_ (.A(_0332_),
    .B(_0334_),
    .C(_0335_),
    .D(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__and3_1 _0779_ (.A(_0292_),
    .B(_0330_),
    .C(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ),
    .Y(_0339_));
 sky130_fd_sc_hd__o311a_1 _0781_ (.A1(_0086_),
    .A2(_0339_),
    .A3(_0237_),
    .B1(_0273_),
    .C1(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ),
    .X(_0340_));
 sky130_fd_sc_hd__and2_1 _0782_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_1 _0783_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ),
    .Y(_0342_));
 sky130_fd_sc_hd__nor2_1 _0784_ (.A(_0341_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__nor2_1 _0785_ (.A(_0086_),
    .B(_0093_),
    .Y(_0344_));
 sky130_fd_sc_hd__or4_1 _0786_ (.A(_0097_),
    .B(_0230_),
    .C(_0231_),
    .D(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__a2bb2o_1 _0787_ (.A1_N(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ),
    .A2_N(_0277_),
    .B1(_0343_),
    .B2(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _0788_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .B(_0341_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_1 _0789_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .B(_0341_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _0790_ (.A(_0347_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__and3_1 _0791_ (.A(_0224_),
    .B(_0227_),
    .C(_0264_),
    .X(_0350_));
 sky130_fd_sc_hd__o2bb2a_1 _0792_ (.A1_N(_0349_),
    .A2_N(_0350_),
    .B1(_0345_),
    .B2(_0343_),
    .X(_0351_));
 sky130_fd_sc_hd__o21ai_1 _0793_ (.A1(_0340_),
    .A2(_0346_),
    .B1(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__and2_1 _0794_ (.A(_0108_),
    .B(_0341_),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_1 _0795_ (.A1(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ),
    .A2(_0348_),
    .B1(_0353_),
    .B2(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .X(_0354_));
 sky130_fd_sc_hd__o22a_1 _0796_ (.A1(_0268_),
    .A2(_0354_),
    .B1(_0349_),
    .B2(_0350_),
    .X(_0355_));
 sky130_fd_sc_hd__a31o_1 _0797_ (.A1(_0108_),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ),
    .A3(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .B1(_0339_),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _0798_ (.A1(_0276_),
    .A2(_0356_),
    .B1(_0354_),
    .B2(_0268_),
    .X(_0357_));
 sky130_fd_sc_hd__a21o_1 _0799_ (.A1(_0352_),
    .A2(_0355_),
    .B1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__a31oi_1 _0800_ (.A1(_0108_),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ),
    .A3(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ),
    .B1(_0343_),
    .Y(_0359_));
 sky130_fd_sc_hd__o2bb2a_1 _0801_ (.A1_N(_0254_),
    .A2_N(_0359_),
    .B1(_0276_),
    .B2(_0356_),
    .X(_0360_));
 sky130_fd_sc_hd__a21o_1 _0802_ (.A1(_0347_),
    .A2(_0348_),
    .B1(_0353_),
    .X(_0361_));
 sky130_fd_sc_hd__a2bb2o_1 _0803_ (.A1_N(_0254_),
    .A2_N(_0359_),
    .B1(_0361_),
    .B2(_0249_),
    .X(_0362_));
 sky130_fd_sc_hd__a211o_1 _0804_ (.A1(_0358_),
    .A2(_0360_),
    .B1(_0362_),
    .C1(_0251_),
    .X(_0363_));
 sky130_fd_sc_hd__a21o_1 _0805_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .A2(_0333_),
    .B1(_0238_),
    .X(_0364_));
 sky130_fd_sc_hd__a31o_1 _0806_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ),
    .A2(_0224_),
    .A3(_0227_),
    .B1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ),
    .X(_0365_));
 sky130_fd_sc_hd__o21a_1 _0807_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ),
    .A2(_0365_),
    .B1(_0292_),
    .X(_0366_));
 sky130_fd_sc_hd__or3b_1 _0808_ (.A(_0366_),
    .B(_0242_),
    .C_N(_0075_),
    .X(_0367_));
 sky130_fd_sc_hd__o21ba_1 _0809_ (.A1(_0249_),
    .A2(_0361_),
    .B1_N(_0244_),
    .X(_0368_));
 sky130_fd_sc_hd__o311a_1 _0810_ (.A1(_0077_),
    .A2(_0071_),
    .A3(_0237_),
    .B1(_0367_),
    .C1(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__or4b_1 _0811_ (.A(_0086_),
    .B(_0230_),
    .C(_0231_),
    .D_N(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .X(_0370_));
 sky130_fd_sc_hd__a31oi_1 _0812_ (.A1(_0087_),
    .A2(_0224_),
    .A3(_0227_),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .Y(_0371_));
 sky130_fd_sc_hd__xor2_1 _0813_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ),
    .X(_0372_));
 sky130_fd_sc_hd__xor2_1 _0814_ (.A(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .B(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__o41a_1 _0815_ (.A1(_0097_),
    .A2(_0230_),
    .A3(_0231_),
    .A4(_0344_),
    .B1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__a311o_1 _0816_ (.A1(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .A2(_0273_),
    .A3(_0370_),
    .B1(_0371_),
    .C1(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _0817_ (.A0(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .A1(_0156_),
    .S(_0372_),
    .X(_0376_));
 sky130_fd_sc_hd__xor2_1 _0818_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ),
    .X(_0377_));
 sky130_fd_sc_hd__o21ai_1 _0819_ (.A1(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .Y(_0378_));
 sky130_fd_sc_hd__xnor2_2 _0820_ (.A(_0377_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__xor2_1 _0821_ (.A(_0376_),
    .B(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__o22a_1 _0822_ (.A1(_0345_),
    .A2(_0373_),
    .B1(_0380_),
    .B2(_0265_),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _0823_ (.A(_0265_),
    .B(_0380_),
    .X(_0382_));
 sky130_fd_sc_hd__o21a_1 _0824_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ),
    .A2(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .B1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ),
    .X(_0383_));
 sky130_fd_sc_hd__o21ai_2 _0825_ (.A1(_0111_),
    .A2(_0383_),
    .B1(_0164_),
    .Y(_0384_));
 sky130_fd_sc_hd__or3_1 _0826_ (.A(_0111_),
    .B(_0164_),
    .C(_0383_),
    .X(_0385_));
 sky130_fd_sc_hd__o211ai_1 _0827_ (.A1(_0376_),
    .A2(_0379_),
    .B1(_0384_),
    .C1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a211o_1 _0828_ (.A1(_0384_),
    .A2(_0385_),
    .B1(_0376_),
    .C1(_0379_),
    .X(_0387_));
 sky130_fd_sc_hd__a21oi_1 _0829_ (.A1(_0386_),
    .A2(_0387_),
    .B1(_0268_),
    .Y(_0388_));
 sky130_fd_sc_hd__a211o_1 _0830_ (.A1(_0375_),
    .A2(_0381_),
    .B1(_0382_),
    .C1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__o211a_1 _0831_ (.A1(_0376_),
    .A2(_0379_),
    .B1(_0384_),
    .C1(_0385_),
    .X(_0390_));
 sky130_fd_sc_hd__nand2_1 _0832_ (.A(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ),
    .Y(_0391_));
 sky130_fd_sc_hd__and3_1 _0833_ (.A(_0391_),
    .B(_0167_),
    .C(_0384_),
    .X(_0392_));
 sky130_fd_sc_hd__a21oi_1 _0834_ (.A1(_0391_),
    .A2(_0384_),
    .B1(_0167_),
    .Y(_0393_));
 sky130_fd_sc_hd__or3_1 _0835_ (.A(_0390_),
    .B(_0392_),
    .C(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_1 _0836_ (.A1(_0392_),
    .A2(_0393_),
    .B1(_0390_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_1 _0837_ (.A(_0241_),
    .B(_0256_),
    .Y(_0396_));
 sky130_fd_sc_hd__a21o_1 _0838_ (.A1(_0394_),
    .A2(_0395_),
    .B1(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__or3b_1 _0839_ (.A(_0307_),
    .B(_0390_),
    .C_N(_0387_),
    .X(_0398_));
 sky130_fd_sc_hd__and3_1 _0840_ (.A(_0396_),
    .B(_0394_),
    .C(_0395_),
    .X(_0399_));
 sky130_fd_sc_hd__or3b_1 _0841_ (.A(_0383_),
    .B(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ),
    .C_N(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ),
    .X(_0400_));
 sky130_fd_sc_hd__o211a_1 _0842_ (.A1(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ),
    .A2(_0384_),
    .B1(_0400_),
    .C1(_0167_),
    .X(_0401_));
 sky130_fd_sc_hd__o31ai_2 _0843_ (.A1(_0390_),
    .A2(_0392_),
    .A3(_0393_),
    .B1(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__or4_1 _0844_ (.A(_0390_),
    .B(_0392_),
    .C(_0393_),
    .D(_0401_),
    .X(_0403_));
 sky130_fd_sc_hd__a21oi_1 _0845_ (.A1(_0402_),
    .A2(_0403_),
    .B1(_0275_),
    .Y(_0404_));
 sky130_fd_sc_hd__a311o_1 _0846_ (.A1(_0389_),
    .A2(_0397_),
    .A3(_0398_),
    .B1(_0399_),
    .C1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__a21o_1 _0847_ (.A1(_0168_),
    .A2(_0402_),
    .B1(_0287_),
    .X(_0406_));
 sky130_fd_sc_hd__a31oi_1 _0848_ (.A1(_0275_),
    .A2(_0402_),
    .A3(_0403_),
    .B1(_0251_),
    .Y(_0407_));
 sky130_fd_sc_hd__or4b_1 _0849_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ),
    .B(_0213_),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ),
    .D_N(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ),
    .X(_0408_));
 sky130_fd_sc_hd__o21ai_1 _0850_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ),
    .A2(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ),
    .B1(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__or4b_1 _0851_ (.A(_0225_),
    .B(_0237_),
    .C(_0409_),
    .D_N(_0335_),
    .X(_0410_));
 sky130_fd_sc_hd__a211o_1 _0852_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .A2(_0241_),
    .B1(_0228_),
    .C1(_0245_),
    .X(_0411_));
 sky130_fd_sc_hd__or3b_1 _0853_ (.A(_0411_),
    .B(_0070_),
    .C_N(_0234_),
    .X(_0412_));
 sky130_fd_sc_hd__a32o_1 _0854_ (.A1(_0168_),
    .A2(_0287_),
    .A3(_0402_),
    .B1(_0410_),
    .B2(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__a31oi_1 _0855_ (.A1(_0405_),
    .A2(_0406_),
    .A3(_0407_),
    .B1(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__a31o_1 _0856_ (.A1(_0363_),
    .A2(_0364_),
    .A3(_0369_),
    .B1(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__or3_1 _0857_ (.A(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ),
    .B(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ),
    .C(_0257_),
    .X(_0416_));
 sky130_fd_sc_hd__a31o_1 _0858_ (.A1(_0218_),
    .A2(_0241_),
    .A3(_0416_),
    .B1(_0350_),
    .X(_0417_));
 sky130_fd_sc_hd__a21oi_1 _0859_ (.A1(_0268_),
    .A2(_0417_),
    .B1(_0256_),
    .Y(_0418_));
 sky130_fd_sc_hd__or3_1 _0860_ (.A(_0254_),
    .B(_0248_),
    .C(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__nor2_1 _0861_ (.A(_0249_),
    .B(_0251_),
    .Y(_0420_));
 sky130_fd_sc_hd__and3_1 _0862_ (.A(_0284_),
    .B(_0265_),
    .C(_0307_),
    .X(_0421_));
 sky130_fd_sc_hd__o41a_1 _0863_ (.A1(_0092_),
    .A2(_0265_),
    .A3(_0268_),
    .A4(_0278_),
    .B1(_0250_),
    .X(_0422_));
 sky130_fd_sc_hd__a41o_1 _0864_ (.A1(_0254_),
    .A2(_0396_),
    .A3(_0420_),
    .A4(_0421_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__and3b_1 _0865_ (.A_N(_0064_),
    .B(_0333_),
    .C(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .X(_0424_));
 sky130_fd_sc_hd__and4b_1 _0866_ (.A_N(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ),
    .B(_0061_),
    .C(_0241_),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ),
    .X(_0425_));
 sky130_fd_sc_hd__nand3_1 _0867_ (.A(_0292_),
    .B(_0333_),
    .C(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__o211ai_1 _0868_ (.A1(_0239_),
    .A2(_0424_),
    .B1(_0426_),
    .C1(_0234_),
    .Y(_0427_));
 sky130_fd_sc_hd__a211o_1 _0869_ (.A1(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ),
    .A2(_0241_),
    .B1(_0244_),
    .C1(_0411_),
    .X(_0428_));
 sky130_fd_sc_hd__and3b_1 _0870_ (.A_N(_0423_),
    .B(_0427_),
    .C(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__o31a_1 _0871_ (.A1(_0240_),
    .A2(_0246_),
    .A3(_0291_),
    .B1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__o211a_1 _0872_ (.A1(_0338_),
    .A2(_0415_),
    .B1(_0419_),
    .C1(_0430_),
    .X(\mod.thorkn_vgaclock.io_g ));
 sky130_fd_sc_hd__nor2_1 _0873_ (.A(_0237_),
    .B(_0429_),
    .Y(\mod.thorkn_vgaclock.io_b ));
 sky130_fd_sc_hd__clkbuf_2 _0874_ (.A(net2),
    .X(_0431_));
 sky130_fd_sc_hd__buf_4 _0875_ (.A(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(_0432_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0877_ (.A(_0432_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0878_ (.A(_0432_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0879_ (.A(_0432_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0880_ (.A(_0432_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0881_ (.A(_0432_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0882_ (.A(_0432_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0883_ (.A(_0432_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0884_ (.A(_0432_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0885_ (.A(_0432_),
    .Y(_0009_));
 sky130_fd_sc_hd__buf_4 _0886_ (.A(_0431_),
    .X(_0433_));
 sky130_fd_sc_hd__inv_2 _0887_ (.A(_0433_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(_0433_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0889_ (.A(_0433_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0890_ (.A(_0433_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0891_ (.A(_0433_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0892_ (.A(_0433_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0893_ (.A(_0433_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0894_ (.A(_0433_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0895_ (.A(_0433_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0896_ (.A(_0433_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_4 _0897_ (.A(_0431_),
    .X(_0434_));
 sky130_fd_sc_hd__inv_2 _0898_ (.A(_0434_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0899_ (.A(_0434_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0900_ (.A(_0434_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0901_ (.A(_0434_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0902_ (.A(_0434_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0903_ (.A(_0434_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0904_ (.A(_0434_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0905_ (.A(_0434_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0906_ (.A(_0434_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0907_ (.A(_0434_),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_4 _0908_ (.A(_0431_),
    .X(_0435_));
 sky130_fd_sc_hd__inv_2 _0909_ (.A(_0435_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0910_ (.A(_0435_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0911_ (.A(_0435_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0912_ (.A(_0435_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _0913_ (.A(_0435_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0914_ (.A(_0435_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0915_ (.A(_0435_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0916_ (.A(_0435_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0917_ (.A(_0435_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _0918_ (.A(_0435_),
    .Y(_0039_));
 sky130_fd_sc_hd__buf_4 _0919_ (.A(_0431_),
    .X(_0436_));
 sky130_fd_sc_hd__inv_2 _0920_ (.A(_0436_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0921_ (.A(_0436_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _0922_ (.A(_0436_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0923_ (.A(_0436_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(_0436_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _0925_ (.A(_0436_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _0926_ (.A(_0436_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _0927_ (.A(_0436_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(_0436_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _0929_ (.A(_0436_),
    .Y(_0049_));
 sky130_fd_sc_hd__buf_4 _0930_ (.A(_0431_),
    .X(_0437_));
 sky130_fd_sc_hd__inv_2 _0931_ (.A(_0437_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _0932_ (.A(_0437_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _0933_ (.A(_0437_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(_0437_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _0935_ (.A(_0437_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _0936_ (.A(_0437_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _0937_ (.A(_0437_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _0938_ (.A(_0437_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _0939_ (.A(_0437_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _0940_ (.A(_0437_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _0941_ (.A(_0431_),
    .Y(_0060_));
 sky130_fd_sc_hd__dfrtp_2 _0942_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[0] ),
    .RESET_B(_0000_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0943_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[1] ),
    .RESET_B(_0001_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0944_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[2] ),
    .RESET_B(_0002_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[2] ));
 sky130_fd_sc_hd__dfrtp_2 _0945_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[3] ),
    .RESET_B(_0003_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0946_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[4] ),
    .RESET_B(_0004_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__dfrtp_2 _0947_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[5] ),
    .RESET_B(_0005_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0948_ (.CLK(net15),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[6] ),
    .RESET_B(_0006_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__dfrtp_2 _0949_ (.CLK(net15),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[7] ),
    .RESET_B(_0007_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__dfrtp_1 _0950_ (.CLK(net15),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[8] ),
    .RESET_B(_0008_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[8] ));
 sky130_fd_sc_hd__dfrtp_4 _0951_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext[9] ),
    .RESET_B(_0009_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__dfrtp_2 _0952_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[0] ),
    .RESET_B(_0010_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[0] ));
 sky130_fd_sc_hd__dfrtp_2 _0953_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[1] ),
    .RESET_B(_0011_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0954_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[2] ),
    .RESET_B(_0012_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0955_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[3] ),
    .RESET_B(_0013_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[3] ));
 sky130_fd_sc_hd__dfrtp_2 _0956_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[4] ),
    .RESET_B(_0014_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0957_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[5] ),
    .RESET_B(_0015_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[5] ));
 sky130_fd_sc_hd__dfrtp_2 _0958_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[6] ),
    .RESET_B(_0016_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[6] ));
 sky130_fd_sc_hd__dfrtp_2 _0959_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[7] ),
    .RESET_B(_0017_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ));
 sky130_fd_sc_hd__dfrtp_2 _0960_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[8] ),
    .RESET_B(_0018_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ));
 sky130_fd_sc_hd__dfrtp_2 _0961_ (.CLK(net13),
    .D(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext[9] ),
    .RESET_B(_0019_),
    .Q(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__dfrtp_2 _0962_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[0] ),
    .RESET_B(_0020_),
    .Q(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__dfrtp_2 _0963_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[1] ),
    .RESET_B(_0021_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__dfrtp_2 _0964_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[2] ),
    .RESET_B(_0022_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[2] ));
 sky130_fd_sc_hd__dfrtp_4 _0965_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[3] ),
    .RESET_B(_0023_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[3] ));
 sky130_fd_sc_hd__dfrtp_4 _0966_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[4] ),
    .RESET_B(_0024_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[4] ));
 sky130_fd_sc_hd__dfrtp_2 _0967_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext[5] ),
    .RESET_B(_0025_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[5] ));
 sky130_fd_sc_hd__dfrtp_4 _0968_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[0] ),
    .RESET_B(_0026_),
    .Q(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__dfrtp_4 _0969_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[1] ),
    .RESET_B(_0027_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__dfrtp_2 _0970_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[2] ),
    .RESET_B(_0028_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[2] ));
 sky130_fd_sc_hd__dfrtp_2 _0971_ (.CLK(net14),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[3] ),
    .RESET_B(_0029_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[3] ));
 sky130_fd_sc_hd__dfrtp_2 _0972_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[4] ),
    .RESET_B(_0030_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0973_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext[5] ),
    .RESET_B(_0031_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0974_ (.CLK(net9),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[0] ),
    .RESET_B(_0032_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0975_ (.CLK(net9),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[1] ),
    .RESET_B(_0033_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0976_ (.CLK(net9),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[2] ),
    .RESET_B(_0034_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0977_ (.CLK(net9),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[3] ),
    .RESET_B(_0035_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0978_ (.CLK(net9),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[4] ),
    .RESET_B(_0036_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0979_ (.CLK(net9),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[5] ),
    .RESET_B(_0037_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0980_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[6] ),
    .RESET_B(_0038_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[6] ));
 sky130_fd_sc_hd__dfrtp_1 _0981_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[7] ),
    .RESET_B(_0039_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[7] ));
 sky130_fd_sc_hd__dfrtp_1 _0982_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[8] ),
    .RESET_B(_0040_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[8] ));
 sky130_fd_sc_hd__dfrtp_1 _0983_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[9] ),
    .RESET_B(_0041_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[9] ));
 sky130_fd_sc_hd__dfrtp_1 _0984_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[10] ),
    .RESET_B(_0042_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[10] ));
 sky130_fd_sc_hd__dfrtp_1 _0985_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[11] ),
    .RESET_B(_0043_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[11] ));
 sky130_fd_sc_hd__dfrtp_1 _0986_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[12] ),
    .RESET_B(_0044_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[12] ));
 sky130_fd_sc_hd__dfrtp_1 _0987_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[13] ),
    .RESET_B(_0045_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[13] ));
 sky130_fd_sc_hd__dfrtp_1 _0988_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[14] ),
    .RESET_B(_0046_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[14] ));
 sky130_fd_sc_hd__dfrtp_1 _0989_ (.CLK(net8),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[15] ),
    .RESET_B(_0047_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[15] ));
 sky130_fd_sc_hd__dfrtp_1 _0990_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[16] ),
    .RESET_B(_0048_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[16] ));
 sky130_fd_sc_hd__dfrtp_1 _0991_ (.CLK(net9),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[17] ),
    .RESET_B(_0049_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[17] ));
 sky130_fd_sc_hd__dfrtp_1 _0992_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[18] ),
    .RESET_B(_0050_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[18] ));
 sky130_fd_sc_hd__dfrtp_1 _0993_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[19] ),
    .RESET_B(_0051_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[19] ));
 sky130_fd_sc_hd__dfrtp_1 _0994_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[20] ),
    .RESET_B(_0052_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__dfrtp_1 _0995_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[21] ),
    .RESET_B(_0053_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[21] ));
 sky130_fd_sc_hd__dfrtp_1 _0996_ (.CLK(net11),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[22] ),
    .RESET_B(_0054_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[22] ));
 sky130_fd_sc_hd__dfrtp_1 _0997_ (.CLK(net11),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[23] ),
    .RESET_B(_0055_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ));
 sky130_fd_sc_hd__dfrtp_1 _0998_ (.CLK(net10),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext[24] ),
    .RESET_B(_0056_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[24] ));
 sky130_fd_sc_hd__dfrtp_1 _0999_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[0] ),
    .RESET_B(_0057_),
    .Q(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1000_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[1] ),
    .RESET_B(_0058_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1001_ (.CLK(net11),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[2] ),
    .RESET_B(_0059_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1002_ (.CLK(net12),
    .D(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext[3] ),
    .RESET_B(_0060_),
    .Q(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__conb_1 tiny_user_project_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 tiny_user_project_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 tiny_user_project_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 tiny_user_project_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 tiny_user_project_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 tiny_user_project_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 tiny_user_project_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 tiny_user_project_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 tiny_user_project_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 tiny_user_project_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 tiny_user_project_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 tiny_user_project_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 tiny_user_project_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 tiny_user_project_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 tiny_user_project_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 tiny_user_project_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 tiny_user_project_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 tiny_user_project_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tiny_user_project_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tiny_user_project_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tiny_user_project_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tiny_user_project_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 tiny_user_project_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 tiny_user_project_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 tiny_user_project_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 tiny_user_project_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 tiny_user_project_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 tiny_user_project_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 tiny_user_project_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 tiny_user_project_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 tiny_user_project_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 tiny_user_project_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 tiny_user_project_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 tiny_user_project_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 tiny_user_project_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 tiny_user_project_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 tiny_user_project_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 tiny_user_project_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 tiny_user_project_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tiny_user_project_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tiny_user_project_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tiny_user_project_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tiny_user_project_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tiny_user_project_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tiny_user_project_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tiny_user_project_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tiny_user_project_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tiny_user_project_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tiny_user_project_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tiny_user_project_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tiny_user_project_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tiny_user_project_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tiny_user_project_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 tiny_user_project_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 tiny_user_project_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 tiny_user_project_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 tiny_user_project_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 tiny_user_project_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 tiny_user_project_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 tiny_user_project_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 tiny_user_project_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 tiny_user_project_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 tiny_user_project_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 tiny_user_project_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 tiny_user_project_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 tiny_user_project_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 tiny_user_project_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 tiny_user_project_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 tiny_user_project_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 tiny_user_project_86 (.LO(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__B (.DIODE(_0070_));
 sky130_fd_sc_hd__clkbuf_1 _1074_ (.A(\mod.thorkn_vgaclock.io_h_sync ),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 _1075_ (.A(\mod.thorkn_vgaclock.io_v_sync ),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 _1076_ (.A(\mod.thorkn_vgaclock.io_r ),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 _1077_ (.A(\mod.thorkn_vgaclock.io_g ),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 _1078_ (.A(\mod.thorkn_vgaclock.io_b ),
    .X(net7));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[8]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[9]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(io_out[14]));
 sky130_fd_sc_hd__clkbuf_2 fanout8 (.A(net9),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout9 (.A(net11),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 fanout11 (.A(net15),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout15 (.A(net1),
    .X(net15));
 sky130_fd_sc_hd__conb_1 tiny_user_project_16 (.LO(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A1 (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__B (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0469__A1 (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0468__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0466__A1 (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0465__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0455__A (.DIODE(_0070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A2 (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A2 (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__A1 (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A2_N (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0454__B (.DIODE(_0071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__A (.DIODE(_0072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__A (.DIODE(_0072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0468__D (.DIODE(_0072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0455__D (.DIODE(_0072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0484__B (.DIODE(_0073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0478__B (.DIODE(_0073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0471__B (.DIODE(_0073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0466__C1 (.DIODE(_0073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0456__B1 (.DIODE(_0073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__C_N (.DIODE(_0075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__B1 (.DIODE(_0075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0459__B (.DIODE(_0075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0469__A3 (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0466__A2 (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0465__B (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0464__A (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0488__A (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0485__A2 (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0474__B (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__A (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__A (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__A1 (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__A (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__A (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__A1 (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__A (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0487__A (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0486__A1 (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0485__A1 (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__A1 (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A1 (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__A (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__A (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0483__A (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0478__A (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__B1_N (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__A2 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__B (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__A (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__A (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0493__B1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0481__A (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__B (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__A (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__B (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__A2 (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__B (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__B (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__A (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0487__B (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0486__B1 (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0483__B (.DIODE(_0093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__A1 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A1 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__A (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__A (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0524__C (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__A2 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__B (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__A (.DIODE(_0125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0531__A2 (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__A2 (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0529__A2 (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__A2 (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__B (.DIODE(_0127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__A1 (.DIODE(_0128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__C1 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__C1 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0614__C1 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__A (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__D (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0566__A3 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0561__B (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__B (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0582__A1 (.DIODE(_0162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__B (.DIODE(_0162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__C (.DIODE(_0162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__A1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__A (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__C (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__A2 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__A3 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__A2 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__B (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__A (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__A3 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__C (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__A2 (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__B (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__A (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__A2 (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__B (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__B (.DIODE(_0211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__B (.DIODE(_0223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__B (.DIODE(_0223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__A (.DIODE(_0223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__A (.DIODE(_0223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A (.DIODE(_0223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__A (.DIODE(_0223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__A2 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__A2 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__A (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A2 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__A2 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__C (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__C1 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__B (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__B1 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__B1 (.DIODE(_0224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__A (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__B (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__B (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__B (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A2 (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__C (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__C (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__C (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__C (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__B (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__B (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__B (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__A (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__A3 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__A3 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__B (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A3 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__A3 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__D (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__B1 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__C (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__B (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__C1 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__B1 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__A (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__A2 (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__B (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__B (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__B (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__A (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__B1 (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__A (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__B1 (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__A3 (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__C (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__C (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__C (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__B (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__C1 (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__B (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__C1 (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A3 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__A3 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__C (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__C (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A2 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__C (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A2 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__A2 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__A (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__C (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A2 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__B (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__A1 (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__C (.DIODE(_0241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__C1 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__B (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__C1 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A2 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__B (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__B (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__B (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__A1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__B2 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0777__B (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__A1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__B (.DIODE(_0251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__B1 (.DIODE(_0251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__C1 (.DIODE(_0251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__C1 (.DIODE(_0251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__A2 (.DIODE(_0251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__D1 (.DIODE(_0251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A_N (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__B (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A2 (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__B (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__B (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__A2 (.DIODE(_0255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__B (.DIODE(_0255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__B1 (.DIODE(_0256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__B (.DIODE(_0256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A3 (.DIODE(_0256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A2 (.DIODE(_0256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__C (.DIODE(_0256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__C (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__A4 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A4 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A3 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__D (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__B1 (.DIODE(_0258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__D (.DIODE(_0258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A2 (.DIODE(_0259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__B1 (.DIODE(_0259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__C (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__B1 (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__D (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__C_N (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A2 (.DIODE(_0265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__B (.DIODE(_0265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__A (.DIODE(_0265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__B2 (.DIODE(_0265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__A (.DIODE(_0265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__A2_N (.DIODE(_0265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__A2 (.DIODE(_0265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A3 (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__A1 (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__B1 (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__B2 (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A1 (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__B1_N (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__A3 (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__B (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__A (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__C_N (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__A2 (.DIODE(_0273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__B1 (.DIODE(_0273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__C (.DIODE(_0273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__B (.DIODE(_0273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__B1 (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__B1 (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__A1 (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__B2 (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__A1 (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__D (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__B (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__B (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A2 (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__B1 (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__C1 (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__A1 (.DIODE(_0301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__A1 (.DIODE(_0301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A1 (.DIODE(_0301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__B (.DIODE(_0301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__A (.DIODE(_0301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A2 (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__C (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__B (.DIODE(_0315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__A1_N (.DIODE(_0315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__B (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__B (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__B (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__B1 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__B2 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__B1 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__A4 (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__D (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__A2 (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__A2 (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__B (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__B2 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__A2_N (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__B1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__B1 (.DIODE(_0353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__A2_N (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__A2_N (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__B (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__B1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__C (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__B1 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A1 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__B1 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__C1 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A2 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__C1 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__A (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A1 (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__B (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__B1 (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__A (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__B (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__A1 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__B (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__C (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A3 (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__A2 (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__C (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__B (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A1 (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__C (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__A (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__B1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__A3 (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__A2 (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__A3 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__B1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0930__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0880__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0891__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__A (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0916__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0912__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0925__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0931__A (.DIODE(_0437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__A0 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__A (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__B (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0566__A2 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__B (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0561__A (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__A (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0508__C (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__A (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__A0 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__B (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0535__B (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0532__A (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__D (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__C1 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0524__A (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0505__A (.DIODE(\mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__C (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__A2 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__B (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__A2 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0513__C (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0515__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__A1_N (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0524__B (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__A2 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A2 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__B (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__B (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0529__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__A3 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A3 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__B2 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0531__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0527__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__B (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0535__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__C (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__B1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__D_N (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0566__A1 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0565__B2 (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0508__D (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0580__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0578__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0507__A (.DIODE(\mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0442__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0440__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0439__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0438__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__D (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0448__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0446__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0445__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A1_N (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0458__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0449__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0448__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0458__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0456__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0453__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0451__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A2 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__D_N (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__A2 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0460__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0458__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0453__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0461__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0454__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__C1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__C1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0469__A2 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0468__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0467__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0455__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.h_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__B2 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0477__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0473__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0472__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0493__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0492__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0484__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__C1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0498__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0497__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0480__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__A1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0500__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0480__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__C1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__C1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__B (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__A (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__B1 (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0483__C (.DIODE(\mod.thorkn_vgaclock.vga_sync_gen.v_counter_value[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0944__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0943__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__CLK (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0951__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0964__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__CLK (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__CLK (.DIODE(net14));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_327 ();
 assign io_oeb[0] = net16;
 assign io_oeb[10] = net26;
 assign io_oeb[11] = net27;
 assign io_oeb[12] = net28;
 assign io_oeb[13] = net29;
 assign io_oeb[14] = net30;
 assign io_oeb[15] = net31;
 assign io_oeb[16] = net32;
 assign io_oeb[17] = net33;
 assign io_oeb[18] = net34;
 assign io_oeb[19] = net35;
 assign io_oeb[1] = net17;
 assign io_oeb[20] = net36;
 assign io_oeb[21] = net37;
 assign io_oeb[22] = net38;
 assign io_oeb[23] = net39;
 assign io_oeb[24] = net40;
 assign io_oeb[25] = net41;
 assign io_oeb[26] = net42;
 assign io_oeb[27] = net43;
 assign io_oeb[28] = net44;
 assign io_oeb[29] = net45;
 assign io_oeb[2] = net18;
 assign io_oeb[30] = net46;
 assign io_oeb[31] = net47;
 assign io_oeb[32] = net48;
 assign io_oeb[33] = net49;
 assign io_oeb[34] = net50;
 assign io_oeb[35] = net51;
 assign io_oeb[36] = net52;
 assign io_oeb[37] = net53;
 assign io_oeb[3] = net19;
 assign io_oeb[4] = net20;
 assign io_oeb[5] = net21;
 assign io_oeb[6] = net22;
 assign io_oeb[7] = net23;
 assign io_oeb[8] = net24;
 assign io_oeb[9] = net25;
 assign io_out[0] = net54;
 assign io_out[15] = net64;
 assign io_out[16] = net65;
 assign io_out[17] = net66;
 assign io_out[18] = net67;
 assign io_out[19] = net68;
 assign io_out[1] = net55;
 assign io_out[20] = net69;
 assign io_out[21] = net70;
 assign io_out[22] = net71;
 assign io_out[23] = net72;
 assign io_out[24] = net73;
 assign io_out[25] = net74;
 assign io_out[26] = net75;
 assign io_out[27] = net76;
 assign io_out[28] = net77;
 assign io_out[29] = net78;
 assign io_out[2] = net56;
 assign io_out[30] = net79;
 assign io_out[31] = net80;
 assign io_out[32] = net81;
 assign io_out[33] = net82;
 assign io_out[34] = net83;
 assign io_out[35] = net84;
 assign io_out[36] = net85;
 assign io_out[37] = net86;
 assign io_out[3] = net57;
 assign io_out[4] = net58;
 assign io_out[5] = net59;
 assign io_out[6] = net60;
 assign io_out[7] = net61;
 assign io_out[8] = net62;
 assign io_out[9] = net63;
endmodule

