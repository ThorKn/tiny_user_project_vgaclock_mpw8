magic
tech sky130A
magscale 1 2
timestamp 1672533676
<< viali >>
rect 18245 32521 18279 32555
rect 18797 32521 18831 32555
rect 24593 32521 24627 32555
rect 21465 32453 21499 32487
rect 1593 32385 1627 32419
rect 2237 32385 2271 32419
rect 2881 32385 2915 32419
rect 4629 32385 4663 32419
rect 5825 32385 5859 32419
rect 8217 32385 8251 32419
rect 9413 32385 9447 32419
rect 11805 32385 11839 32419
rect 13001 32385 13035 32419
rect 15393 32385 15427 32419
rect 16865 32385 16899 32419
rect 19441 32385 19475 32419
rect 20177 32385 20211 32419
rect 22569 32385 22603 32419
rect 23765 32385 23799 32419
rect 25329 32385 25363 32419
rect 26157 32385 26191 32419
rect 27353 32385 27387 32419
rect 29745 32385 29779 32419
rect 30941 32385 30975 32419
rect 14933 32249 14967 32283
rect 20821 32249 20855 32283
rect 28365 32249 28399 32283
rect 12449 32181 12483 32215
rect 13645 32181 13679 32215
rect 14381 32181 14415 32215
rect 16221 32181 16255 32215
rect 17785 32181 17819 32215
rect 22017 32181 22051 32215
rect 23305 32181 23339 32215
rect 28917 32181 28951 32215
rect 30481 32181 30515 32215
rect 1593 31977 1627 32011
rect 15485 31977 15519 32011
rect 18797 31977 18831 32011
rect 19901 31977 19935 32011
rect 21189 31977 21223 32011
rect 22017 31977 22051 32011
rect 23121 31977 23155 32011
rect 23857 31977 23891 32011
rect 24685 31977 24719 32011
rect 25237 31977 25271 32011
rect 26525 31977 26559 32011
rect 28181 31977 28215 32011
rect 30573 31977 30607 32011
rect 20637 31909 20671 31943
rect 22569 31909 22603 31943
rect 25881 31909 25915 31943
rect 31217 31909 31251 31943
rect 13737 31841 13771 31875
rect 27629 31841 27663 31875
rect 12081 31773 12115 31807
rect 15025 31773 15059 31807
rect 16681 31773 16715 31807
rect 24593 31773 24627 31807
rect 24777 31773 24811 31807
rect 25237 31773 25271 31807
rect 25421 31773 25455 31807
rect 25881 31773 25915 31807
rect 26065 31773 26099 31807
rect 29745 31773 29779 31807
rect 31033 31773 31067 31807
rect 14473 31705 14507 31739
rect 17693 31705 17727 31739
rect 27077 31705 27111 31739
rect 28733 31705 28767 31739
rect 11529 31637 11563 31671
rect 12541 31637 12575 31671
rect 13185 31637 13219 31671
rect 16129 31637 16163 31671
rect 17233 31637 17267 31671
rect 18245 31637 18279 31671
rect 15209 31433 15243 31467
rect 18429 31433 18463 31467
rect 24961 31433 24995 31467
rect 28273 31433 28307 31467
rect 21189 31365 21223 31399
rect 22109 31365 22143 31399
rect 27721 31365 27755 31399
rect 13553 31297 13587 31331
rect 19073 31297 19107 31331
rect 23489 31297 23523 31331
rect 24133 31297 24167 31331
rect 24317 31297 24351 31331
rect 25145 31297 25179 31331
rect 25789 31297 25823 31331
rect 26249 31297 26283 31331
rect 26341 31297 26375 31331
rect 11897 31161 11931 31195
rect 16313 31161 16347 31195
rect 17877 31161 17911 31195
rect 28825 31161 28859 31195
rect 1593 31093 1627 31127
rect 10517 31093 10551 31127
rect 11161 31093 11195 31127
rect 12449 31093 12483 31127
rect 12909 31093 12943 31127
rect 14013 31093 14047 31127
rect 14657 31093 14691 31127
rect 15669 31093 15703 31127
rect 17325 31093 17359 31127
rect 19717 31093 19751 31127
rect 20637 31093 20671 31127
rect 22845 31093 22879 31127
rect 23581 31093 23615 31127
rect 24317 31093 24351 31127
rect 25697 31093 25731 31127
rect 27261 31093 27295 31127
rect 30021 31093 30055 31127
rect 30665 31093 30699 31127
rect 31309 31093 31343 31127
rect 10333 30889 10367 30923
rect 16129 30889 16163 30923
rect 17693 30889 17727 30923
rect 18337 30889 18371 30923
rect 18797 30889 18831 30923
rect 21833 30889 21867 30923
rect 24777 30889 24811 30923
rect 24961 30889 24995 30923
rect 25605 30889 25639 30923
rect 28825 30889 28859 30923
rect 26433 30821 26467 30855
rect 26525 30821 26559 30855
rect 11437 30753 11471 30787
rect 13185 30753 13219 30787
rect 27077 30753 27111 30787
rect 11989 30685 12023 30719
rect 13737 30685 13771 30719
rect 14473 30685 14507 30719
rect 22477 30685 22511 30719
rect 22661 30685 22695 30719
rect 23121 30685 23155 30719
rect 23305 30685 23339 30719
rect 23765 30685 23799 30719
rect 26525 30685 26559 30719
rect 26985 30685 27019 30719
rect 27629 30685 27663 30719
rect 27813 30685 27847 30719
rect 28365 30685 28399 30719
rect 29929 30685 29963 30719
rect 31309 30685 31343 30719
rect 9873 30617 9907 30651
rect 17141 30617 17175 30651
rect 22569 30617 22603 30651
rect 24593 30617 24627 30651
rect 24793 30617 24827 30651
rect 25421 30617 25455 30651
rect 25621 30617 25655 30651
rect 26249 30617 26283 30651
rect 27721 30617 27755 30651
rect 10977 30549 11011 30583
rect 12541 30549 12575 30583
rect 14933 30549 14967 30583
rect 15577 30549 15611 30583
rect 16589 30549 16623 30583
rect 19533 30549 19567 30583
rect 20361 30549 20395 30583
rect 20913 30549 20947 30583
rect 23213 30549 23247 30583
rect 23949 30549 23983 30583
rect 25789 30549 25823 30583
rect 30113 30549 30147 30583
rect 30573 30549 30607 30583
rect 17785 30345 17819 30379
rect 23841 30345 23875 30379
rect 24711 30345 24745 30379
rect 8953 30277 8987 30311
rect 9965 30277 9999 30311
rect 10609 30277 10643 30311
rect 13553 30277 13587 30311
rect 16313 30277 16347 30311
rect 19717 30277 19751 30311
rect 20453 30277 20487 30311
rect 21005 30277 21039 30311
rect 23029 30277 23063 30311
rect 23213 30277 23247 30311
rect 24041 30277 24075 30311
rect 24501 30277 24535 30311
rect 26433 30277 26467 30311
rect 14657 30209 14691 30243
rect 22293 30209 22327 30243
rect 22477 30209 22511 30243
rect 22937 30209 22971 30243
rect 25513 30209 25547 30243
rect 26249 30209 26283 30243
rect 27169 30209 27203 30243
rect 27353 30209 27387 30243
rect 27813 30209 27847 30243
rect 27997 30209 28031 30243
rect 28457 30209 28491 30243
rect 29101 30209 29135 30243
rect 29745 30209 29779 30243
rect 30389 30209 30423 30243
rect 31033 30209 31067 30243
rect 1593 30141 1627 30175
rect 11161 30141 11195 30175
rect 15117 30141 15151 30175
rect 25329 30141 25363 30175
rect 25697 30141 25731 30175
rect 18245 30073 18279 30107
rect 24869 30073 24903 30107
rect 29285 30073 29319 30107
rect 9505 30005 9539 30039
rect 11805 30005 11839 30039
rect 12449 30005 12483 30039
rect 13001 30005 13035 30039
rect 14105 30005 14139 30039
rect 15761 30005 15795 30039
rect 17233 30005 17267 30039
rect 18889 30005 18923 30039
rect 22477 30005 22511 30039
rect 23121 30005 23155 30039
rect 23673 30005 23707 30039
rect 23857 30005 23891 30039
rect 24685 30005 24719 30039
rect 27261 30005 27295 30039
rect 27813 30005 27847 30039
rect 28641 30005 28675 30039
rect 29929 30005 29963 30039
rect 30573 30005 30607 30039
rect 31217 30005 31251 30039
rect 8585 29801 8619 29835
rect 13185 29801 13219 29835
rect 14841 29801 14875 29835
rect 18153 29801 18187 29835
rect 20177 29801 20211 29835
rect 20913 29801 20947 29835
rect 23673 29801 23707 29835
rect 25697 29801 25731 29835
rect 25881 29801 25915 29835
rect 26617 29801 26651 29835
rect 9873 29733 9907 29767
rect 18705 29733 18739 29767
rect 22201 29733 22235 29767
rect 23213 29733 23247 29767
rect 24041 29733 24075 29767
rect 28089 29733 28123 29767
rect 10977 29665 11011 29699
rect 15945 29665 15979 29699
rect 24961 29665 24995 29699
rect 25145 29665 25179 29699
rect 27353 29665 27387 29699
rect 10333 29597 10367 29631
rect 20821 29597 20855 29631
rect 21465 29597 21499 29631
rect 21649 29597 21683 29631
rect 22109 29597 22143 29631
rect 22385 29597 22419 29631
rect 22937 29597 22971 29631
rect 23029 29597 23063 29631
rect 23673 29597 23707 29631
rect 23857 29597 23891 29631
rect 24869 29597 24903 29631
rect 25237 29597 25271 29631
rect 26525 29597 26559 29631
rect 26617 29597 26651 29631
rect 28089 29597 28123 29631
rect 28273 29597 28307 29631
rect 28825 29597 28859 29631
rect 28917 29597 28951 29631
rect 29929 29597 29963 29631
rect 30389 29597 30423 29631
rect 31309 29597 31343 29631
rect 11529 29529 11563 29563
rect 12633 29529 12667 29563
rect 19441 29529 19475 29563
rect 22293 29529 22327 29563
rect 26065 29529 26099 29563
rect 27537 29529 27571 29563
rect 9229 29461 9263 29495
rect 12081 29461 12115 29495
rect 13737 29461 13771 29495
rect 15393 29461 15427 29495
rect 16497 29461 16531 29495
rect 16957 29461 16991 29495
rect 17601 29461 17635 29495
rect 21465 29461 21499 29495
rect 24869 29461 24903 29495
rect 25865 29461 25899 29495
rect 26893 29461 26927 29495
rect 30573 29461 30607 29495
rect 8401 29257 8435 29291
rect 12449 29257 12483 29291
rect 15209 29257 15243 29291
rect 16957 29257 16991 29291
rect 20637 29257 20671 29291
rect 25421 29257 25455 29291
rect 26617 29257 26651 29291
rect 28917 29257 28951 29291
rect 30205 29257 30239 29291
rect 7849 29189 7883 29223
rect 9505 29189 9539 29223
rect 17509 29189 17543 29223
rect 22477 29189 22511 29223
rect 23581 29189 23615 29223
rect 24409 29189 24443 29223
rect 25605 29189 25639 29223
rect 28089 29189 28123 29223
rect 11805 29121 11839 29155
rect 18061 29121 18095 29155
rect 19073 29121 19107 29155
rect 19901 29121 19935 29155
rect 19993 29121 20027 29155
rect 20085 29121 20119 29155
rect 20545 29121 20579 29155
rect 21189 29121 21223 29155
rect 21373 29131 21407 29165
rect 22661 29121 22695 29155
rect 23305 29121 23339 29155
rect 23673 29121 23707 29155
rect 24593 29121 24627 29155
rect 24685 29121 24719 29155
rect 24869 29121 24903 29155
rect 24961 29121 24995 29155
rect 26433 29121 26467 29155
rect 26617 29121 26651 29155
rect 27169 29121 27203 29155
rect 27997 29121 28031 29155
rect 28273 29121 28307 29155
rect 28733 29121 28767 29155
rect 28917 29121 28951 29155
rect 29377 29121 29411 29155
rect 29561 29121 29595 29155
rect 30021 29121 30055 29155
rect 31033 29121 31067 29155
rect 8953 29053 8987 29087
rect 10517 29053 10551 29087
rect 14657 29053 14691 29087
rect 21281 29053 21315 29087
rect 23489 29053 23523 29087
rect 25973 29053 26007 29087
rect 27261 29053 27295 29087
rect 9965 28985 9999 29019
rect 11161 28985 11195 29019
rect 13001 28985 13035 29019
rect 16221 28985 16255 29019
rect 18521 28985 18555 29019
rect 22845 28985 22879 29019
rect 23305 28985 23339 29019
rect 27537 28985 27571 29019
rect 28273 28985 28307 29019
rect 29469 28985 29503 29019
rect 31217 28985 31251 29019
rect 13553 28917 13587 28951
rect 14105 28917 14139 28951
rect 15761 28917 15795 28951
rect 25605 28917 25639 28951
rect 27353 28917 27387 28951
rect 9873 28713 9907 28747
rect 11989 28713 12023 28747
rect 12541 28713 12575 28747
rect 13737 28713 13771 28747
rect 15853 28713 15887 28747
rect 17141 28713 17175 28747
rect 20361 28713 20395 28747
rect 22845 28713 22879 28747
rect 25789 28713 25823 28747
rect 26985 28713 27019 28747
rect 28365 28713 28399 28747
rect 28733 28713 28767 28747
rect 17601 28645 17635 28679
rect 21281 28645 21315 28679
rect 23949 28645 23983 28679
rect 25145 28645 25179 28679
rect 26617 28645 26651 28679
rect 7481 28577 7515 28611
rect 10885 28577 10919 28611
rect 21097 28577 21131 28611
rect 23765 28577 23799 28611
rect 24685 28577 24719 28611
rect 24869 28577 24903 28611
rect 25881 28577 25915 28611
rect 1593 28509 1627 28543
rect 8033 28509 8067 28543
rect 13185 28509 13219 28543
rect 18705 28509 18739 28543
rect 19901 28509 19935 28543
rect 20545 28509 20579 28543
rect 20637 28509 20671 28543
rect 21373 28509 21407 28543
rect 22201 28509 22235 28543
rect 24041 28509 24075 28543
rect 24777 28509 24811 28543
rect 24961 28509 24995 28543
rect 26157 28509 26191 28543
rect 26801 28509 26835 28543
rect 26893 28509 26927 28543
rect 27077 28509 27111 28543
rect 27537 28509 27571 28543
rect 28370 28509 28404 28543
rect 28549 28509 28583 28543
rect 29929 28509 29963 28543
rect 30389 28509 30423 28543
rect 31033 28509 31067 28543
rect 14749 28441 14783 28475
rect 20361 28441 20395 28475
rect 21097 28441 21131 28475
rect 22017 28441 22051 28475
rect 22661 28441 22695 28475
rect 22861 28441 22895 28475
rect 27721 28441 27755 28475
rect 27905 28441 27939 28475
rect 8493 28373 8527 28407
rect 9321 28373 9355 28407
rect 10425 28373 10459 28407
rect 11529 28373 11563 28407
rect 15209 28373 15243 28407
rect 16589 28373 16623 28407
rect 18153 28373 18187 28407
rect 18797 28373 18831 28407
rect 19809 28373 19843 28407
rect 21833 28373 21867 28407
rect 23029 28373 23063 28407
rect 23581 28373 23615 28407
rect 25605 28373 25639 28407
rect 29837 28373 29871 28407
rect 30481 28373 30515 28407
rect 31217 28373 31251 28407
rect 7297 28169 7331 28203
rect 13921 28169 13955 28203
rect 14749 28169 14783 28203
rect 15301 28169 15335 28203
rect 16221 28169 16255 28203
rect 18429 28169 18463 28203
rect 19073 28169 19107 28203
rect 21373 28169 21407 28203
rect 24041 28169 24075 28203
rect 24133 28169 24167 28203
rect 28181 28169 28215 28203
rect 30205 28169 30239 28203
rect 9505 28101 9539 28135
rect 12817 28101 12851 28135
rect 13277 28101 13311 28135
rect 17233 28101 17267 28135
rect 20453 28101 20487 28135
rect 22017 28101 22051 28135
rect 22201 28101 22235 28135
rect 24409 28101 24443 28135
rect 29285 28101 29319 28135
rect 29469 28101 29503 28135
rect 18325 28033 18359 28067
rect 18521 28033 18555 28067
rect 18981 28033 19015 28067
rect 19165 28033 19199 28067
rect 19717 28033 19751 28067
rect 20361 28033 20395 28067
rect 20637 28033 20671 28067
rect 21097 28033 21131 28067
rect 21281 28033 21315 28067
rect 22845 28033 22879 28067
rect 22937 28033 22971 28067
rect 23048 28033 23082 28067
rect 23213 28033 23247 28067
rect 23397 28033 23431 28067
rect 24225 28033 24259 28067
rect 24869 28033 24903 28067
rect 25237 28033 25271 28067
rect 26061 28033 26095 28067
rect 26157 28033 26191 28067
rect 26342 28033 26376 28067
rect 27261 28033 27295 28067
rect 27353 28033 27387 28067
rect 27445 28033 27479 28067
rect 28365 28033 28399 28067
rect 28457 28033 28491 28067
rect 28641 28033 28675 28067
rect 29101 28033 29135 28067
rect 30205 28033 30239 28067
rect 31033 28033 31067 28067
rect 12173 27965 12207 27999
rect 26249 27965 26283 27999
rect 27537 27965 27571 27999
rect 29929 27965 29963 27999
rect 8861 27897 8895 27931
rect 10609 27897 10643 27931
rect 19901 27897 19935 27931
rect 20637 27897 20671 27931
rect 22385 27897 22419 27931
rect 25881 27897 25915 27931
rect 30113 27897 30147 27931
rect 1593 27829 1627 27863
rect 7849 27829 7883 27863
rect 8401 27829 8435 27863
rect 9965 27829 9999 27863
rect 11161 27829 11195 27863
rect 17785 27829 17819 27863
rect 23857 27829 23891 27863
rect 25237 27829 25271 27863
rect 25421 27829 25455 27863
rect 27721 27829 27755 27863
rect 28457 27829 28491 27863
rect 31217 27829 31251 27863
rect 16865 27625 16899 27659
rect 17509 27625 17543 27659
rect 19901 27625 19935 27659
rect 21189 27625 21223 27659
rect 24777 27625 24811 27659
rect 26065 27625 26099 27659
rect 28917 27625 28951 27659
rect 29745 27625 29779 27659
rect 29929 27625 29963 27659
rect 11529 27557 11563 27591
rect 12633 27557 12667 27591
rect 15669 27557 15703 27591
rect 18061 27557 18095 27591
rect 18797 27557 18831 27591
rect 22293 27557 22327 27591
rect 22845 27557 22879 27591
rect 26249 27557 26283 27591
rect 26709 27557 26743 27591
rect 27261 27557 27295 27591
rect 27997 27557 28031 27591
rect 30665 27557 30699 27591
rect 9321 27489 9355 27523
rect 10333 27489 10367 27523
rect 13737 27489 13771 27523
rect 14565 27489 14599 27523
rect 18889 27489 18923 27523
rect 20729 27489 20763 27523
rect 21281 27489 21315 27523
rect 24961 27489 24995 27523
rect 28089 27489 28123 27523
rect 30573 27489 30607 27523
rect 16221 27421 16255 27455
rect 17325 27421 17359 27455
rect 17509 27421 17543 27455
rect 17969 27421 18003 27455
rect 18613 27421 18647 27455
rect 18705 27421 18739 27455
rect 19625 27421 19659 27455
rect 19901 27421 19935 27455
rect 20545 27421 20579 27455
rect 21189 27421 21223 27455
rect 22569 27421 22603 27455
rect 23305 27421 23339 27455
rect 23397 27421 23431 27455
rect 23581 27421 23615 27455
rect 23673 27421 23707 27455
rect 23857 27421 23891 27455
rect 24777 27421 24811 27455
rect 25237 27421 25271 27455
rect 25697 27421 25731 27455
rect 26065 27421 26099 27455
rect 26985 27421 27019 27455
rect 27917 27421 27951 27455
rect 28193 27421 28227 27455
rect 30757 27421 30791 27455
rect 30849 27421 30883 27455
rect 29883 27387 29917 27421
rect 7389 27353 7423 27387
rect 8033 27353 8067 27387
rect 12081 27353 12115 27387
rect 15025 27353 15059 27387
rect 19717 27353 19751 27387
rect 20361 27353 20395 27387
rect 27721 27353 27755 27387
rect 29101 27353 29135 27387
rect 30113 27353 30147 27387
rect 6377 27285 6411 27319
rect 6929 27285 6963 27319
rect 8585 27285 8619 27319
rect 9873 27285 9907 27319
rect 10885 27285 10919 27319
rect 13185 27285 13219 27319
rect 21557 27285 21591 27319
rect 22477 27285 22511 27319
rect 22661 27285 22695 27319
rect 24593 27285 24627 27319
rect 26893 27285 26927 27319
rect 27077 27285 27111 27319
rect 28733 27285 28767 27319
rect 28901 27285 28935 27319
rect 8401 27081 8435 27115
rect 10057 27081 10091 27115
rect 11161 27081 11195 27115
rect 15209 27081 15243 27115
rect 15669 27081 15703 27115
rect 21097 27081 21131 27115
rect 21465 27081 21499 27115
rect 24041 27081 24075 27115
rect 24409 27081 24443 27115
rect 27353 27081 27387 27115
rect 28181 27081 28215 27115
rect 28365 27081 28399 27115
rect 30481 27081 30515 27115
rect 31309 27081 31343 27115
rect 6745 27013 6779 27047
rect 12449 27013 12483 27047
rect 17969 27013 18003 27047
rect 20545 27013 20579 27047
rect 27169 27013 27203 27047
rect 29193 27013 29227 27047
rect 29653 27013 29687 27047
rect 30113 27013 30147 27047
rect 30941 27013 30975 27047
rect 20315 26979 20349 27013
rect 16221 26945 16255 26979
rect 17233 26945 17267 26979
rect 17417 26945 17451 26979
rect 18153 26945 18187 26979
rect 18889 26945 18923 26979
rect 19349 26945 19383 26979
rect 19533 26945 19567 26979
rect 21005 26945 21039 26979
rect 21281 26945 21315 26979
rect 22017 26945 22051 26979
rect 22569 26945 22603 26979
rect 22661 26945 22695 26979
rect 22845 26945 22879 26979
rect 22937 26945 22971 26979
rect 24225 26945 24259 26979
rect 25053 26945 25087 26979
rect 25362 26945 25396 26979
rect 25513 26945 25547 26979
rect 26203 26945 26237 26979
rect 26341 26945 26375 26979
rect 26433 26945 26467 26979
rect 26617 26945 26651 26979
rect 27445 26945 27479 26979
rect 27537 26945 27571 26979
rect 27721 26945 27755 26979
rect 29561 26945 29595 26979
rect 30297 26945 30331 26979
rect 31125 26945 31159 26979
rect 7849 26877 7883 26911
rect 14105 26877 14139 26911
rect 18613 26877 18647 26911
rect 23765 26877 23799 26911
rect 23857 26877 23891 26911
rect 24133 26877 24167 26911
rect 28733 26877 28767 26911
rect 29285 26877 29319 26911
rect 8953 26809 8987 26843
rect 19717 26809 19751 26843
rect 20177 26809 20211 26843
rect 29377 26809 29411 26843
rect 7297 26741 7331 26775
rect 9505 26741 9539 26775
rect 10517 26741 10551 26775
rect 11805 26741 11839 26775
rect 13001 26741 13035 26775
rect 13461 26741 13495 26775
rect 14565 26741 14599 26775
rect 17417 26741 17451 26775
rect 18705 26741 18739 26775
rect 18797 26741 18831 26775
rect 19441 26741 19475 26775
rect 20361 26741 20395 26775
rect 23121 26741 23155 26775
rect 24869 26741 24903 26775
rect 25973 26741 26007 26775
rect 28343 26741 28377 26775
rect 8585 26537 8619 26571
rect 11529 26537 11563 26571
rect 12541 26537 12575 26571
rect 13093 26537 13127 26571
rect 14657 26537 14691 26571
rect 17141 26537 17175 26571
rect 17233 26537 17267 26571
rect 18889 26537 18923 26571
rect 19993 26537 20027 26571
rect 20913 26537 20947 26571
rect 29745 26537 29779 26571
rect 30941 26537 30975 26571
rect 10885 26469 10919 26503
rect 19809 26469 19843 26503
rect 20729 26469 20763 26503
rect 25789 26469 25823 26503
rect 27997 26469 28031 26503
rect 30665 26469 30699 26503
rect 5825 26401 5859 26435
rect 10425 26401 10459 26435
rect 15853 26401 15887 26435
rect 17325 26401 17359 26435
rect 17785 26401 17819 26435
rect 17969 26401 18003 26435
rect 19901 26401 19935 26435
rect 21005 26401 21039 26435
rect 21833 26401 21867 26435
rect 25329 26401 25363 26435
rect 26065 26401 26099 26435
rect 27537 26401 27571 26435
rect 1593 26333 1627 26367
rect 9321 26333 9355 26367
rect 15761 26333 15795 26367
rect 15945 26333 15979 26367
rect 16405 26333 16439 26367
rect 16589 26333 16623 26367
rect 17050 26333 17084 26367
rect 18061 26333 18095 26367
rect 18613 26333 18647 26367
rect 18705 26333 18739 26367
rect 20085 26333 20119 26367
rect 21281 26333 21315 26367
rect 22003 26333 22037 26367
rect 23121 26333 23155 26367
rect 23213 26333 23247 26367
rect 23581 26333 23615 26367
rect 24869 26333 24903 26367
rect 25053 26333 25087 26367
rect 25237 26333 25271 26367
rect 25973 26333 26007 26367
rect 26157 26333 26191 26367
rect 26249 26333 26283 26367
rect 26433 26333 26467 26367
rect 26893 26333 26927 26367
rect 27077 26333 27111 26367
rect 27172 26333 27206 26367
rect 27307 26333 27341 26367
rect 28181 26333 28215 26367
rect 28273 26333 28307 26367
rect 28365 26333 28399 26367
rect 29009 26333 29043 26367
rect 29101 26333 29135 26367
rect 29929 26333 29963 26367
rect 30205 26333 30239 26367
rect 30849 26333 30883 26367
rect 31033 26333 31067 26367
rect 6377 26265 6411 26299
rect 6929 26265 6963 26299
rect 7941 26265 7975 26299
rect 9781 26265 9815 26299
rect 12081 26265 12115 26299
rect 15209 26265 15243 26299
rect 20269 26265 20303 26299
rect 23397 26265 23431 26299
rect 23489 26265 23523 26299
rect 24593 26265 24627 26299
rect 28549 26265 28583 26299
rect 7481 26197 7515 26231
rect 13645 26197 13679 26231
rect 16589 26197 16623 26231
rect 17785 26197 17819 26231
rect 22293 26197 22327 26231
rect 23765 26197 23799 26231
rect 24961 26197 24995 26231
rect 30113 26197 30147 26231
rect 5457 25993 5491 26027
rect 12173 25993 12207 26027
rect 13829 25993 13863 26027
rect 22109 25993 22143 26027
rect 22293 25993 22327 26027
rect 23305 25993 23339 26027
rect 25789 25993 25823 26027
rect 25881 25993 25915 26027
rect 29285 25993 29319 26027
rect 30757 25993 30791 26027
rect 8953 25925 8987 25959
rect 11161 25925 11195 25959
rect 17509 25925 17543 25959
rect 24777 25925 24811 25959
rect 27813 25925 27847 25959
rect 14841 25857 14875 25891
rect 15025 25857 15059 25891
rect 15485 25857 15519 25891
rect 16129 25857 16163 25891
rect 16313 25857 16347 25891
rect 17325 25857 17359 25891
rect 18153 25857 18187 25891
rect 18337 25857 18371 25891
rect 19165 25857 19199 25891
rect 19453 25857 19487 25891
rect 20085 25857 20119 25891
rect 20177 25857 20211 25891
rect 20269 25857 20303 25891
rect 20913 25857 20947 25891
rect 22290 25857 22324 25891
rect 27169 25857 27203 25891
rect 27353 25857 27387 25891
rect 27445 25857 27479 25891
rect 27537 25857 27571 25891
rect 28641 25857 28675 25891
rect 29469 25857 29503 25891
rect 29561 25857 29595 25891
rect 29837 25857 29871 25891
rect 30297 25857 30331 25891
rect 30389 25857 30423 25891
rect 30573 25857 30607 25891
rect 9505 25789 9539 25823
rect 10057 25789 10091 25823
rect 13185 25789 13219 25823
rect 15577 25789 15611 25823
rect 18981 25789 19015 25823
rect 19901 25789 19935 25823
rect 20361 25789 20395 25823
rect 21189 25789 21223 25823
rect 22747 25789 22781 25823
rect 25053 25789 25087 25823
rect 25697 25789 25731 25823
rect 28733 25789 28767 25823
rect 29745 25789 29779 25823
rect 6009 25721 6043 25755
rect 7849 25721 7883 25755
rect 15025 25721 15059 25755
rect 18521 25721 18555 25755
rect 21465 25721 21499 25755
rect 22661 25721 22695 25755
rect 26249 25721 26283 25755
rect 28273 25721 28307 25755
rect 6745 25653 6779 25687
rect 7297 25653 7331 25687
rect 8401 25653 8435 25687
rect 10609 25653 10643 25687
rect 12725 25653 12759 25687
rect 14289 25653 14323 25687
rect 16221 25653 16255 25687
rect 17693 25653 17727 25687
rect 19349 25653 19383 25687
rect 21281 25653 21315 25687
rect 31217 25653 31251 25687
rect 5273 25449 5307 25483
rect 6285 25449 6319 25483
rect 7389 25449 7423 25483
rect 8033 25449 8067 25483
rect 10333 25449 10367 25483
rect 11897 25449 11931 25483
rect 13645 25449 13679 25483
rect 14749 25449 14783 25483
rect 15301 25449 15335 25483
rect 16129 25449 16163 25483
rect 16773 25449 16807 25483
rect 17141 25449 17175 25483
rect 18889 25449 18923 25483
rect 20361 25449 20395 25483
rect 21189 25449 21223 25483
rect 24041 25449 24075 25483
rect 26893 25449 26927 25483
rect 28457 25449 28491 25483
rect 29929 25449 29963 25483
rect 30941 25449 30975 25483
rect 9781 25381 9815 25415
rect 16313 25381 16347 25415
rect 28641 25381 28675 25415
rect 31309 25381 31343 25415
rect 8585 25313 8619 25347
rect 19644 25313 19678 25347
rect 21465 25313 21499 25347
rect 22569 25313 22603 25347
rect 24869 25313 24903 25347
rect 28273 25313 28307 25347
rect 1593 25245 1627 25279
rect 6929 25245 6963 25279
rect 13553 25245 13587 25279
rect 14657 25245 14691 25279
rect 14841 25245 14875 25279
rect 15289 25245 15323 25279
rect 15485 25245 15519 25279
rect 16773 25245 16807 25279
rect 16957 25245 16991 25279
rect 17601 25245 17635 25279
rect 18429 25245 18463 25279
rect 18547 25245 18581 25279
rect 19441 25245 19475 25279
rect 19533 25245 19567 25279
rect 20361 25245 20395 25279
rect 20729 25245 20763 25279
rect 21373 25245 21407 25279
rect 21557 25245 21591 25279
rect 21649 25245 21683 25279
rect 21833 25245 21867 25279
rect 22293 25245 22327 25279
rect 24593 25245 24627 25279
rect 27031 25245 27065 25279
rect 27169 25245 27203 25279
rect 27261 25245 27295 25279
rect 27389 25245 27423 25279
rect 27537 25245 27571 25279
rect 27997 25245 28031 25279
rect 28457 25245 28491 25279
rect 29929 25245 29963 25279
rect 30297 25245 30331 25279
rect 9229 25177 9263 25211
rect 15945 25177 15979 25211
rect 17785 25177 17819 25211
rect 19717 25177 19751 25211
rect 29193 25177 29227 25211
rect 5825 25109 5859 25143
rect 10793 25109 10827 25143
rect 11437 25109 11471 25143
rect 12449 25109 12483 25143
rect 13093 25109 13127 25143
rect 16145 25109 16179 25143
rect 17969 25109 18003 25143
rect 18705 25109 18739 25143
rect 20177 25109 20211 25143
rect 26341 25109 26375 25143
rect 29745 25109 29779 25143
rect 30757 25109 30791 25143
rect 30941 25109 30975 25143
rect 10057 24905 10091 24939
rect 12081 24905 12115 24939
rect 13185 24905 13219 24939
rect 21189 24905 21223 24939
rect 26617 24905 26651 24939
rect 29745 24905 29779 24939
rect 15117 24837 15151 24871
rect 15945 24837 15979 24871
rect 16161 24837 16195 24871
rect 16957 24837 16991 24871
rect 21373 24837 21407 24871
rect 27418 24837 27452 24871
rect 4905 24769 4939 24803
rect 5457 24769 5491 24803
rect 9413 24769 9447 24803
rect 13093 24769 13127 24803
rect 13277 24769 13311 24803
rect 13737 24769 13771 24803
rect 14381 24769 14415 24803
rect 14473 24769 14507 24803
rect 14667 24769 14701 24803
rect 15301 24769 15335 24803
rect 17141 24769 17175 24803
rect 17969 24769 18003 24803
rect 18981 24769 19015 24803
rect 19165 24769 19199 24803
rect 19993 24769 20027 24803
rect 22017 24769 22051 24803
rect 22201 24769 22235 24803
rect 22293 24769 22327 24803
rect 22385 24769 22419 24803
rect 25605 24769 25639 24803
rect 25881 24769 25915 24803
rect 25973 24769 26007 24803
rect 26341 24769 26375 24803
rect 26617 24769 26651 24803
rect 27322 24769 27356 24803
rect 27813 24769 27847 24803
rect 28549 24769 28583 24803
rect 28641 24769 28675 24803
rect 28733 24769 28767 24803
rect 28917 24769 28951 24803
rect 29653 24769 29687 24803
rect 29862 24769 29896 24803
rect 30481 24769 30515 24803
rect 30665 24769 30699 24803
rect 30757 24769 30791 24803
rect 30941 24769 30975 24803
rect 7297 24701 7331 24735
rect 11069 24701 11103 24735
rect 13829 24701 13863 24735
rect 14584 24701 14618 24735
rect 15485 24701 15519 24735
rect 17877 24701 17911 24735
rect 18889 24701 18923 24735
rect 19073 24701 19107 24735
rect 19901 24701 19935 24735
rect 20821 24701 20855 24735
rect 21005 24701 21039 24735
rect 21097 24701 21131 24735
rect 21465 24701 21499 24735
rect 23305 24701 23339 24735
rect 23581 24701 23615 24735
rect 29377 24701 29411 24735
rect 6009 24633 6043 24667
rect 6745 24633 6779 24667
rect 8401 24633 8435 24667
rect 12541 24633 12575 24667
rect 16313 24633 16347 24667
rect 30849 24633 30883 24667
rect 7757 24565 7791 24599
rect 8953 24565 8987 24599
rect 10609 24565 10643 24599
rect 16129 24565 16163 24599
rect 17325 24565 17359 24599
rect 18245 24565 18279 24599
rect 19349 24565 19383 24599
rect 20269 24565 20303 24599
rect 22661 24565 22695 24599
rect 25053 24565 25087 24599
rect 27169 24565 27203 24599
rect 27721 24565 27755 24599
rect 28273 24565 28307 24599
rect 30021 24565 30055 24599
rect 4169 24361 4203 24395
rect 7941 24361 7975 24395
rect 14749 24361 14783 24395
rect 15117 24361 15151 24395
rect 15761 24361 15795 24395
rect 18337 24361 18371 24395
rect 21575 24361 21609 24395
rect 24041 24361 24075 24395
rect 28641 24361 28675 24395
rect 30389 24361 30423 24395
rect 31033 24361 31067 24395
rect 5825 24293 5859 24327
rect 12909 24293 12943 24327
rect 16497 24293 16531 24327
rect 16865 24293 16899 24327
rect 18705 24293 18739 24327
rect 26341 24293 26375 24327
rect 29193 24293 29227 24327
rect 5273 24225 5307 24259
rect 12357 24225 12391 24259
rect 16405 24225 16439 24259
rect 17601 24225 17635 24259
rect 22293 24225 22327 24259
rect 22569 24225 22603 24259
rect 24869 24225 24903 24259
rect 31033 24225 31067 24259
rect 10149 24157 10183 24191
rect 12265 24157 12299 24191
rect 12449 24157 12483 24191
rect 12909 24157 12943 24191
rect 13093 24157 13127 24191
rect 13553 24157 13587 24191
rect 14749 24157 14783 24191
rect 14841 24157 14875 24191
rect 16681 24157 16715 24191
rect 17509 24157 17543 24191
rect 17693 24157 17727 24191
rect 17785 24157 17819 24191
rect 18521 24157 18555 24191
rect 18613 24157 18647 24191
rect 18797 24157 18831 24191
rect 19441 24157 19475 24191
rect 19625 24157 19659 24191
rect 21833 24157 21867 24191
rect 24593 24157 24627 24191
rect 26893 24157 26927 24191
rect 29745 24157 29779 24191
rect 29929 24157 29963 24191
rect 30021 24157 30055 24191
rect 30113 24157 30147 24191
rect 31125 24157 31159 24191
rect 4721 24089 4755 24123
rect 6929 24089 6963 24123
rect 8493 24089 8527 24123
rect 15577 24089 15611 24123
rect 15777 24089 15811 24123
rect 27169 24089 27203 24123
rect 30849 24089 30883 24123
rect 6285 24021 6319 24055
rect 7481 24021 7515 24055
rect 9505 24021 9539 24055
rect 10701 24021 10735 24055
rect 11253 24021 11287 24055
rect 11805 24021 11839 24055
rect 13645 24021 13679 24055
rect 15945 24021 15979 24055
rect 17325 24021 17359 24055
rect 19441 24021 19475 24055
rect 20085 24021 20119 24055
rect 31309 24021 31343 24055
rect 4353 23817 4387 23851
rect 7297 23817 7331 23851
rect 9505 23817 9539 23851
rect 12173 23817 12207 23851
rect 14397 23817 14431 23851
rect 15393 23817 15427 23851
rect 29561 23817 29595 23851
rect 30665 23817 30699 23851
rect 6745 23749 6779 23783
rect 14197 23749 14231 23783
rect 15025 23749 15059 23783
rect 15241 23749 15275 23783
rect 17785 23749 17819 23783
rect 21005 23749 21039 23783
rect 25237 23749 25271 23783
rect 31217 23749 31251 23783
rect 4905 23681 4939 23715
rect 12173 23681 12207 23715
rect 12357 23681 12391 23715
rect 12817 23681 12851 23715
rect 13461 23681 13495 23715
rect 15853 23681 15887 23715
rect 15945 23681 15979 23715
rect 16129 23681 16163 23715
rect 17233 23681 17267 23715
rect 17325 23681 17359 23715
rect 17509 23681 17543 23715
rect 17601 23681 17635 23715
rect 18429 23681 18463 23715
rect 18613 23681 18647 23715
rect 18797 23681 18831 23715
rect 19441 23681 19475 23715
rect 19533 23681 19567 23715
rect 19716 23681 19750 23715
rect 19905 23703 19939 23737
rect 20361 23681 20395 23715
rect 20524 23681 20558 23715
rect 20624 23684 20658 23718
rect 20749 23681 20783 23715
rect 22017 23681 22051 23715
rect 22201 23681 22235 23715
rect 22477 23681 22511 23715
rect 23213 23681 23247 23715
rect 27169 23681 27203 23715
rect 27353 23681 27387 23715
rect 27629 23681 27663 23715
rect 27905 23681 27939 23715
rect 27997 23681 28031 23715
rect 28641 23681 28675 23715
rect 28733 23681 28767 23715
rect 29745 23681 29779 23715
rect 30021 23681 30055 23715
rect 30205 23681 30239 23715
rect 30941 23681 30975 23715
rect 1593 23613 1627 23647
rect 5457 23613 5491 23647
rect 6009 23613 6043 23647
rect 9965 23613 9999 23647
rect 13737 23613 13771 23647
rect 18705 23613 18739 23647
rect 23489 23613 23523 23647
rect 26249 23613 26283 23647
rect 26525 23613 26559 23647
rect 29009 23613 29043 23647
rect 29101 23613 29135 23647
rect 30849 23613 30883 23647
rect 31309 23613 31343 23647
rect 8401 23545 8435 23579
rect 14565 23545 14599 23579
rect 19625 23545 19659 23579
rect 22293 23545 22327 23579
rect 28457 23545 28491 23579
rect 7849 23477 7883 23511
rect 8861 23477 8895 23511
rect 10609 23477 10643 23511
rect 11069 23477 11103 23511
rect 13001 23477 13035 23511
rect 13553 23477 13587 23511
rect 13645 23477 13679 23511
rect 14381 23477 14415 23511
rect 15209 23477 15243 23511
rect 16313 23477 16347 23511
rect 19257 23477 19291 23511
rect 22385 23477 22419 23511
rect 22753 23477 22787 23511
rect 4169 23273 4203 23307
rect 5825 23273 5859 23307
rect 9229 23273 9263 23307
rect 9689 23273 9723 23307
rect 10333 23273 10367 23307
rect 14657 23273 14691 23307
rect 14841 23273 14875 23307
rect 28365 23273 28399 23307
rect 28641 23273 28675 23307
rect 28825 23273 28859 23307
rect 4721 23205 4755 23239
rect 11345 23205 11379 23239
rect 12633 23205 12667 23239
rect 15485 23205 15519 23239
rect 26985 23205 27019 23239
rect 17785 23137 17819 23171
rect 18245 23137 18279 23171
rect 22293 23137 22327 23171
rect 28733 23137 28767 23171
rect 29745 23137 29779 23171
rect 31309 23137 31343 23171
rect 1593 23069 1627 23103
rect 5273 23069 5307 23103
rect 11345 23069 11379 23103
rect 11529 23069 11563 23103
rect 11989 23069 12023 23103
rect 12633 23069 12667 23103
rect 12817 23069 12851 23103
rect 12909 23069 12943 23103
rect 13553 23069 13587 23103
rect 14473 23069 14507 23103
rect 14657 23069 14691 23103
rect 15393 23069 15427 23103
rect 15669 23069 15703 23103
rect 15761 23069 15795 23103
rect 16221 23069 16255 23103
rect 16313 23069 16347 23103
rect 16497 23069 16531 23103
rect 16589 23069 16623 23103
rect 16773 23069 16807 23103
rect 17233 23069 17267 23103
rect 17325 23069 17359 23103
rect 17509 23069 17543 23103
rect 17601 23069 17635 23103
rect 18429 23069 18463 23103
rect 18521 23069 18555 23103
rect 18613 23069 18647 23103
rect 18751 23069 18785 23103
rect 18889 23069 18923 23103
rect 19901 23069 19935 23103
rect 20085 23069 20119 23103
rect 20177 23069 20211 23103
rect 20269 23069 20303 23103
rect 21097 23069 21131 23103
rect 21281 23069 21315 23103
rect 21557 23069 21591 23103
rect 21833 23069 21867 23103
rect 24041 23069 24075 23103
rect 26341 23069 26375 23103
rect 26893 23069 26927 23103
rect 27077 23069 27111 23103
rect 27629 23069 27663 23103
rect 28917 23069 28951 23103
rect 29101 23069 29135 23103
rect 30021 23069 30055 23103
rect 30110 23069 30144 23103
rect 30205 23069 30239 23103
rect 30389 23069 30423 23103
rect 30849 23069 30883 23103
rect 31125 23069 31159 23103
rect 6377 23001 6411 23035
rect 13369 23001 13403 23035
rect 15301 23001 15335 23035
rect 21005 23001 21039 23035
rect 23765 23001 23799 23035
rect 26065 23001 26099 23035
rect 6837 22933 6871 22967
rect 7389 22933 7423 22967
rect 7941 22933 7975 22967
rect 8585 22933 8619 22967
rect 10885 22933 10919 22967
rect 12081 22933 12115 22967
rect 13737 22933 13771 22967
rect 20545 22933 20579 22967
rect 24593 22933 24627 22967
rect 30941 22933 30975 22967
rect 4353 22729 4387 22763
rect 7113 22729 7147 22763
rect 8217 22729 8251 22763
rect 11161 22729 11195 22763
rect 12449 22729 12483 22763
rect 12536 22729 12570 22763
rect 13277 22729 13311 22763
rect 14381 22729 14415 22763
rect 16313 22729 16347 22763
rect 19901 22729 19935 22763
rect 30941 22729 30975 22763
rect 31033 22729 31067 22763
rect 5365 22661 5399 22695
rect 7665 22661 7699 22695
rect 10425 22661 10459 22695
rect 12633 22661 12667 22695
rect 14013 22661 14047 22695
rect 14933 22661 14967 22695
rect 15301 22661 15335 22695
rect 18521 22661 18555 22695
rect 20361 22661 20395 22695
rect 31125 22661 31159 22695
rect 10333 22593 10367 22627
rect 10517 22593 10551 22627
rect 10977 22593 11011 22627
rect 11161 22593 11195 22627
rect 11713 22593 11747 22627
rect 12725 22593 12759 22627
rect 13185 22593 13219 22627
rect 13411 22593 13445 22627
rect 13553 22593 13587 22627
rect 14197 22593 14231 22627
rect 14841 22593 14875 22627
rect 15117 22593 15151 22627
rect 15945 22593 15979 22627
rect 17325 22593 17359 22627
rect 18337 22593 18371 22627
rect 18429 22593 18463 22627
rect 18705 22593 18739 22627
rect 18797 22593 18831 22627
rect 19625 22593 19659 22627
rect 19742 22593 19776 22627
rect 21373 22593 21407 22627
rect 22201 22593 22235 22627
rect 23765 22593 23799 22627
rect 23949 22593 23983 22627
rect 26341 22593 26375 22627
rect 27237 22593 27271 22627
rect 27629 22593 27663 22627
rect 28365 22593 28399 22627
rect 28641 22593 28675 22627
rect 29101 22593 29135 22627
rect 29561 22593 29595 22627
rect 29745 22593 29779 22627
rect 29929 22593 29963 22627
rect 30113 22593 30147 22627
rect 12357 22525 12391 22559
rect 15853 22525 15887 22559
rect 17233 22525 17267 22559
rect 19257 22525 19291 22559
rect 19533 22525 19567 22559
rect 22477 22525 22511 22559
rect 22937 22525 22971 22559
rect 26065 22525 26099 22559
rect 27445 22525 27479 22559
rect 29837 22525 29871 22559
rect 30757 22525 30791 22559
rect 4905 22457 4939 22491
rect 9229 22457 9263 22491
rect 9873 22457 9907 22491
rect 11805 22457 11839 22491
rect 17693 22457 17727 22491
rect 18153 22457 18187 22491
rect 24593 22457 24627 22491
rect 28733 22457 28767 22491
rect 28825 22457 28859 22491
rect 31309 22457 31343 22491
rect 6009 22389 6043 22423
rect 8769 22389 8803 22423
rect 13553 22389 13587 22423
rect 22017 22389 22051 22423
rect 22385 22389 22419 22423
rect 27353 22389 27387 22423
rect 27537 22389 27571 22423
rect 27905 22389 27939 22423
rect 28917 22389 28951 22423
rect 30297 22389 30331 22423
rect 5825 22185 5859 22219
rect 6377 22185 6411 22219
rect 11989 22185 12023 22219
rect 14289 22185 14323 22219
rect 14473 22185 14507 22219
rect 23409 22185 23443 22219
rect 29101 22185 29135 22219
rect 9689 22117 9723 22151
rect 11069 22117 11103 22151
rect 16681 22117 16715 22151
rect 21925 22117 21959 22151
rect 5273 22049 5307 22083
rect 10885 22049 10919 22083
rect 12817 22049 12851 22083
rect 15393 22049 15427 22083
rect 15669 22049 15703 22083
rect 16221 22049 16255 22083
rect 18889 22049 18923 22083
rect 19625 22049 19659 22083
rect 26157 22049 26191 22083
rect 26893 22049 26927 22083
rect 29101 22049 29135 22083
rect 4721 21981 4755 22015
rect 9597 21981 9631 22015
rect 10241 21981 10275 22015
rect 10333 21981 10367 22015
rect 11161 21981 11195 22015
rect 11621 21981 11655 22015
rect 11805 21981 11839 22015
rect 12449 21981 12483 22015
rect 12633 21981 12667 22015
rect 13461 21981 13495 22015
rect 13737 21981 13771 22015
rect 15301 21981 15335 22015
rect 16313 21981 16347 22015
rect 17417 21981 17451 22015
rect 17509 21981 17543 22015
rect 17601 21981 17635 22015
rect 17785 21981 17819 22015
rect 18245 21981 18279 22015
rect 18429 21981 18463 22015
rect 18521 21981 18555 22015
rect 18613 21981 18647 22015
rect 21373 21981 21407 22015
rect 23666 21981 23700 22015
rect 26433 21981 26467 22015
rect 27261 21981 27295 22015
rect 27997 21981 28031 22015
rect 28733 21981 28767 22015
rect 28825 21981 28859 22015
rect 29009 21981 29043 22015
rect 29745 21981 29779 22015
rect 30113 21981 30147 22015
rect 30205 21981 30239 22015
rect 30849 21981 30883 22015
rect 31033 21981 31067 22015
rect 31309 21981 31343 22015
rect 6929 21913 6963 21947
rect 8033 21913 8067 21947
rect 14457 21913 14491 21947
rect 14657 21913 14691 21947
rect 17141 21913 17175 21947
rect 21097 21913 21131 21947
rect 29837 21913 29871 21947
rect 4169 21845 4203 21879
rect 7481 21845 7515 21879
rect 8493 21845 8527 21879
rect 11161 21845 11195 21879
rect 13277 21845 13311 21879
rect 13645 21845 13679 21879
rect 24685 21845 24719 21879
rect 27654 21845 27688 21879
rect 30389 21845 30423 21879
rect 31125 21845 31159 21879
rect 5457 21641 5491 21675
rect 5917 21641 5951 21675
rect 7941 21641 7975 21675
rect 8493 21641 8527 21675
rect 11161 21641 11195 21675
rect 12265 21641 12299 21675
rect 14289 21641 14323 21675
rect 17233 21641 17267 21675
rect 18521 21641 18555 21675
rect 18613 21641 18647 21675
rect 4905 21573 4939 21607
rect 13001 21573 13035 21607
rect 17601 21573 17635 21607
rect 21465 21573 21499 21607
rect 27445 21573 27479 21607
rect 29653 21573 29687 21607
rect 29745 21573 29779 21607
rect 9781 21505 9815 21539
rect 10241 21505 10275 21539
rect 10885 21505 10919 21539
rect 10977 21505 11011 21539
rect 12173 21505 12207 21539
rect 12541 21505 12575 21539
rect 13185 21505 13219 21539
rect 14105 21505 14139 21539
rect 15117 21505 15151 21539
rect 15945 21505 15979 21539
rect 17417 21505 17451 21539
rect 17509 21505 17543 21539
rect 17785 21505 17819 21539
rect 19441 21505 19475 21539
rect 23857 21505 23891 21539
rect 26617 21505 26651 21539
rect 29377 21505 29411 21539
rect 29469 21505 29503 21539
rect 29837 21505 29871 21539
rect 30481 21505 30515 21539
rect 30665 21505 30699 21539
rect 30757 21505 30791 21539
rect 30849 21505 30883 21539
rect 9689 21437 9723 21471
rect 11161 21437 11195 21471
rect 12357 21437 12391 21471
rect 13829 21437 13863 21471
rect 13921 21437 13955 21471
rect 14749 21437 14783 21471
rect 15209 21437 15243 21471
rect 15853 21437 15887 21471
rect 18429 21437 18463 21471
rect 19717 21437 19751 21471
rect 23581 21437 23615 21471
rect 26341 21437 26375 21471
rect 27169 21437 27203 21471
rect 6929 21369 6963 21403
rect 10425 21369 10459 21403
rect 12541 21369 12575 21403
rect 22109 21369 22143 21403
rect 24869 21369 24903 21403
rect 1593 21301 1627 21335
rect 7481 21301 7515 21335
rect 9045 21301 9079 21335
rect 13369 21301 13403 21335
rect 16313 21301 16347 21335
rect 18981 21301 19015 21335
rect 28917 21301 28951 21335
rect 30021 21301 30055 21335
rect 31125 21301 31159 21335
rect 5273 21097 5307 21131
rect 12541 21097 12575 21131
rect 14473 21097 14507 21131
rect 16589 21097 16623 21131
rect 24777 21097 24811 21131
rect 30849 21097 30883 21131
rect 31309 21097 31343 21131
rect 14289 21029 14323 21063
rect 15117 21029 15151 21063
rect 18889 21029 18923 21063
rect 29745 21029 29779 21063
rect 6929 20961 6963 20995
rect 11253 20961 11287 20995
rect 12725 20961 12759 20995
rect 13737 20961 13771 20995
rect 16405 20961 16439 20995
rect 22017 20961 22051 20995
rect 23581 20961 23615 20995
rect 30113 20961 30147 20995
rect 30941 20961 30975 20995
rect 9689 20893 9723 20927
rect 10333 20893 10367 20927
rect 10517 20893 10551 20927
rect 10977 20893 11011 20927
rect 11069 20893 11103 20927
rect 11713 20893 11747 20927
rect 11897 20893 11931 20927
rect 12081 20893 12115 20927
rect 12541 20893 12575 20927
rect 12909 20893 12943 20927
rect 13362 20893 13396 20927
rect 15393 20893 15427 20927
rect 15485 20893 15519 20927
rect 16313 20893 16347 20927
rect 17129 20893 17163 20927
rect 17325 20893 17359 20927
rect 17417 20893 17451 20927
rect 17509 20893 17543 20927
rect 18245 20893 18279 20927
rect 18429 20893 18463 20927
rect 18521 20893 18555 20927
rect 18613 20893 18647 20927
rect 19993 20893 20027 20927
rect 22753 20893 22787 20927
rect 23213 20893 23247 20927
rect 26525 20893 26559 20927
rect 26974 20893 27008 20927
rect 30389 20893 30423 20927
rect 31125 20893 31159 20927
rect 9137 20825 9171 20859
rect 13461 20825 13495 20859
rect 14657 20825 14691 20859
rect 17785 20825 17819 20859
rect 20276 20825 20310 20859
rect 26249 20825 26283 20859
rect 27261 20825 27295 20859
rect 29904 20825 29938 20859
rect 30849 20825 30883 20859
rect 5825 20757 5859 20791
rect 6377 20757 6411 20791
rect 7389 20757 7423 20791
rect 8033 20757 8067 20791
rect 8585 20757 8619 20791
rect 9781 20757 9815 20791
rect 10425 20757 10459 20791
rect 11253 20757 11287 20791
rect 12817 20757 12851 20791
rect 13553 20757 13587 20791
rect 13737 20757 13771 20791
rect 14457 20757 14491 20791
rect 15301 20757 15335 20791
rect 15669 20757 15703 20791
rect 19533 20757 19567 20791
rect 28733 20757 28767 20791
rect 30021 20757 30055 20791
rect 6929 20553 6963 20587
rect 7941 20553 7975 20587
rect 10425 20553 10459 20587
rect 12449 20553 12483 20587
rect 14121 20553 14155 20587
rect 16313 20553 16347 20587
rect 23765 20553 23799 20587
rect 5917 20485 5951 20519
rect 13093 20485 13127 20519
rect 13293 20485 13327 20519
rect 13921 20485 13955 20519
rect 17509 20485 17543 20519
rect 17877 20485 17911 20519
rect 8585 20417 8619 20451
rect 9597 20417 9631 20451
rect 10241 20417 10275 20451
rect 10425 20417 10459 20451
rect 10885 20417 10919 20451
rect 10977 20417 11011 20451
rect 11161 20417 11195 20451
rect 11713 20417 11747 20451
rect 11897 20417 11931 20451
rect 12357 20417 12391 20451
rect 12633 20417 12667 20451
rect 14933 20417 14967 20451
rect 15761 20417 15795 20451
rect 16865 20417 16899 20451
rect 17693 20417 17727 20451
rect 17785 20417 17819 20451
rect 18521 20417 18555 20451
rect 18705 20417 18739 20451
rect 18797 20417 18831 20451
rect 18889 20417 18923 20451
rect 26525 20417 26559 20451
rect 27169 20417 27203 20451
rect 29837 20417 29871 20451
rect 30665 20417 30699 20451
rect 30757 20417 30791 20451
rect 31033 20417 31067 20451
rect 1593 20349 1627 20383
rect 15025 20349 15059 20383
rect 15301 20349 15335 20383
rect 16037 20349 16071 20383
rect 21189 20349 21223 20383
rect 21465 20349 21499 20383
rect 22017 20349 22051 20383
rect 22293 20349 22327 20383
rect 26249 20349 26283 20383
rect 27445 20349 27479 20383
rect 29929 20349 29963 20383
rect 30941 20349 30975 20383
rect 5457 20281 5491 20315
rect 9689 20281 9723 20315
rect 11805 20281 11839 20315
rect 12633 20281 12667 20315
rect 16957 20281 16991 20315
rect 19165 20281 19199 20315
rect 19717 20281 19751 20315
rect 24777 20281 24811 20315
rect 29469 20281 29503 20315
rect 7389 20213 7423 20247
rect 9045 20213 9079 20247
rect 11161 20213 11195 20247
rect 13277 20213 13311 20247
rect 13461 20213 13495 20247
rect 14105 20213 14139 20247
rect 14289 20213 14323 20247
rect 15853 20213 15887 20247
rect 18061 20213 18095 20247
rect 28917 20213 28951 20247
rect 30481 20213 30515 20247
rect 8493 20009 8527 20043
rect 10609 20009 10643 20043
rect 13737 20009 13771 20043
rect 22569 20009 22603 20043
rect 26893 20009 26927 20043
rect 11437 19941 11471 19975
rect 11897 19941 11931 19975
rect 14473 19941 14507 19975
rect 27445 19941 27479 19975
rect 16221 19873 16255 19907
rect 16681 19873 16715 19907
rect 17509 19873 17543 19907
rect 17785 19873 17819 19907
rect 23213 19873 23247 19907
rect 26341 19873 26375 19907
rect 27261 19873 27295 19907
rect 27353 19873 27387 19907
rect 28641 19873 28675 19907
rect 28733 19873 28767 19907
rect 30205 19873 30239 19907
rect 30757 19873 30791 19907
rect 31217 19873 31251 19907
rect 7481 19805 7515 19839
rect 10517 19805 10551 19839
rect 10701 19805 10735 19839
rect 11161 19805 11195 19839
rect 11437 19805 11471 19839
rect 11897 19805 11931 19839
rect 12081 19805 12115 19839
rect 12173 19805 12207 19839
rect 13553 19805 13587 19839
rect 13737 19805 13771 19839
rect 14841 19805 14875 19839
rect 15485 19805 15519 19839
rect 15761 19805 15795 19839
rect 16589 19805 16623 19839
rect 17417 19805 17451 19839
rect 18245 19805 18279 19839
rect 18429 19805 18463 19839
rect 18521 19805 18555 19839
rect 18613 19805 18647 19839
rect 19441 19805 19475 19839
rect 20085 19805 20119 19839
rect 22753 19805 22787 19839
rect 23489 19805 23523 19839
rect 24593 19805 24627 19839
rect 27169 19805 27203 19839
rect 27629 19805 27663 19839
rect 28270 19805 28304 19839
rect 29929 19805 29963 19839
rect 30021 19805 30055 19839
rect 30297 19805 30331 19839
rect 31125 19805 31159 19839
rect 6377 19737 6411 19771
rect 9505 19737 9539 19771
rect 12725 19737 12759 19771
rect 14657 19737 14691 19771
rect 20361 19737 20395 19771
rect 22109 19737 22143 19771
rect 24869 19737 24903 19771
rect 29745 19737 29779 19771
rect 6929 19669 6963 19703
rect 7941 19669 7975 19703
rect 9965 19669 9999 19703
rect 11253 19669 11287 19703
rect 12817 19669 12851 19703
rect 13369 19669 13403 19703
rect 18889 19669 18923 19703
rect 19625 19669 19659 19703
rect 28089 19669 28123 19703
rect 28273 19669 28307 19703
rect 9965 19465 9999 19499
rect 12810 19465 12844 19499
rect 14473 19465 14507 19499
rect 18061 19465 18095 19499
rect 19165 19465 19199 19499
rect 21373 19465 21407 19499
rect 12081 19397 12115 19431
rect 12909 19397 12943 19431
rect 13369 19397 13403 19431
rect 15761 19397 15795 19431
rect 19006 19397 19040 19431
rect 28273 19397 28307 19431
rect 10977 19329 11011 19363
rect 11069 19329 11103 19363
rect 11989 19329 12023 19363
rect 12633 19329 12667 19363
rect 12725 19329 12759 19363
rect 13645 19329 13679 19363
rect 14289 19329 14323 19363
rect 14933 19329 14967 19363
rect 15853 19329 15887 19363
rect 16129 19329 16163 19363
rect 16313 19329 16347 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17601 19329 17635 19363
rect 17693 19329 17727 19363
rect 17877 19329 17911 19363
rect 18797 19329 18831 19363
rect 22293 19329 22327 19363
rect 26617 19329 26651 19363
rect 27353 19329 27387 19363
rect 27629 19329 27663 19363
rect 27813 19329 27847 19363
rect 28733 19329 28767 19363
rect 29745 19329 29779 19363
rect 30389 19329 30423 19363
rect 30481 19329 30515 19363
rect 30665 19329 30699 19363
rect 30757 19329 30791 19363
rect 7205 19261 7239 19295
rect 14105 19261 14139 19295
rect 15025 19261 15059 19295
rect 16957 19261 16991 19295
rect 17785 19261 17819 19295
rect 18521 19261 18555 19295
rect 18889 19261 18923 19295
rect 19625 19261 19659 19295
rect 19901 19261 19935 19295
rect 22569 19261 22603 19295
rect 27537 19261 27571 19295
rect 28641 19261 28675 19295
rect 29377 19261 29411 19295
rect 29837 19261 29871 19295
rect 8861 19193 8895 19227
rect 13553 19193 13587 19227
rect 15301 19193 15335 19227
rect 24869 19193 24903 19227
rect 27169 19193 27203 19227
rect 27445 19193 27479 19227
rect 6653 19125 6687 19159
rect 7665 19125 7699 19159
rect 8309 19125 8343 19159
rect 9413 19125 9447 19159
rect 10517 19125 10551 19159
rect 13461 19125 13495 19159
rect 14933 19125 14967 19159
rect 24041 19125 24075 19159
rect 26359 19125 26393 19159
rect 28365 19125 28399 19159
rect 28917 19125 28951 19159
rect 30941 19125 30975 19159
rect 14749 18921 14783 18955
rect 16681 18921 16715 18955
rect 17877 18921 17911 18955
rect 19533 18921 19567 18955
rect 23857 18921 23891 18955
rect 27905 18921 27939 18955
rect 29101 18921 29135 18955
rect 31217 18921 31251 18955
rect 10517 18853 10551 18887
rect 13461 18853 13495 18887
rect 16865 18853 16899 18887
rect 17417 18853 17451 18887
rect 18889 18853 18923 18887
rect 22477 18853 22511 18887
rect 23673 18853 23707 18887
rect 27445 18853 27479 18887
rect 29745 18853 29779 18887
rect 9965 18785 9999 18819
rect 15945 18785 15979 18819
rect 18429 18785 18463 18819
rect 20269 18785 20303 18819
rect 23029 18785 23063 18819
rect 26341 18785 26375 18819
rect 26801 18785 26835 18819
rect 27169 18785 27203 18819
rect 28090 18785 28124 18819
rect 28181 18785 28215 18819
rect 28273 18785 28307 18819
rect 28917 18785 28951 18819
rect 30205 18785 30239 18819
rect 1593 18717 1627 18751
rect 11529 18717 11563 18751
rect 12173 18717 12207 18751
rect 12357 18717 12391 18751
rect 12817 18717 12851 18751
rect 13645 18717 13679 18751
rect 13737 18717 13771 18751
rect 16497 18717 16531 18751
rect 16773 18717 16807 18751
rect 17325 18717 17359 18751
rect 17541 18717 17575 18751
rect 17693 18717 17727 18751
rect 18521 18717 18555 18751
rect 19993 18717 20027 18751
rect 22937 18717 22971 18751
rect 28365 18717 28399 18751
rect 29193 18717 29227 18751
rect 30113 18717 30147 18751
rect 30757 18717 30791 18751
rect 31033 18717 31067 18751
rect 7481 18649 7515 18683
rect 13461 18649 13495 18683
rect 14933 18649 14967 18683
rect 15117 18649 15151 18683
rect 15577 18649 15611 18683
rect 15761 18649 15795 18683
rect 16405 18649 16439 18683
rect 22017 18649 22051 18683
rect 22845 18649 22879 18683
rect 23825 18649 23859 18683
rect 24041 18649 24075 18683
rect 26065 18649 26099 18683
rect 27286 18649 27320 18683
rect 28917 18649 28951 18683
rect 30849 18649 30883 18683
rect 7941 18581 7975 18615
rect 8493 18581 8527 18615
rect 9321 18581 9355 18615
rect 10977 18581 11011 18615
rect 11621 18581 11655 18615
rect 12357 18581 12391 18615
rect 12909 18581 12943 18615
rect 24593 18581 24627 18615
rect 27077 18581 27111 18615
rect 10057 18377 10091 18411
rect 12909 18377 12943 18411
rect 15193 18377 15227 18411
rect 15853 18377 15887 18411
rect 17509 18377 17543 18411
rect 21373 18377 21407 18411
rect 25329 18377 25363 18411
rect 27721 18377 27755 18411
rect 31125 18377 31159 18411
rect 8401 18309 8435 18343
rect 12265 18309 12299 18343
rect 14197 18309 14231 18343
rect 15393 18309 15427 18343
rect 16313 18309 16347 18343
rect 17693 18309 17727 18343
rect 17877 18309 17911 18343
rect 19901 18309 19935 18343
rect 22293 18309 22327 18343
rect 25881 18309 25915 18343
rect 27353 18309 27387 18343
rect 29193 18309 29227 18343
rect 14427 18275 14461 18309
rect 12173 18241 12207 18275
rect 12817 18241 12851 18275
rect 13645 18241 13679 18275
rect 16037 18241 16071 18275
rect 17601 18241 17635 18275
rect 18613 18241 18647 18275
rect 19625 18241 19659 18275
rect 24225 18241 24259 18275
rect 24685 18241 24719 18275
rect 25605 18241 25639 18275
rect 26433 18241 26467 18275
rect 26617 18241 26651 18275
rect 27169 18241 27203 18275
rect 27445 18241 27479 18275
rect 27537 18241 27571 18275
rect 28549 18241 28583 18275
rect 29377 18241 29411 18275
rect 29469 18241 29503 18275
rect 29653 18241 29687 18275
rect 29745 18241 29779 18275
rect 30205 18241 30239 18275
rect 31125 18241 31159 18275
rect 31309 18241 31343 18275
rect 16221 18173 16255 18207
rect 18337 18173 18371 18207
rect 22017 18173 22051 18207
rect 24593 18173 24627 18207
rect 25513 18173 25547 18207
rect 25973 18173 26007 18207
rect 28181 18173 28215 18207
rect 28641 18173 28675 18207
rect 30389 18173 30423 18207
rect 8953 18105 8987 18139
rect 13645 18105 13679 18139
rect 14565 18105 14599 18139
rect 26433 18105 26467 18139
rect 1593 18037 1627 18071
rect 9505 18037 9539 18071
rect 10609 18037 10643 18071
rect 11161 18037 11195 18071
rect 14381 18037 14415 18071
rect 15025 18037 15059 18071
rect 15209 18037 15243 18071
rect 16037 18037 16071 18071
rect 17325 18037 17359 18071
rect 23765 18037 23799 18071
rect 24685 18037 24719 18071
rect 24869 18037 24903 18071
rect 9321 17833 9355 17867
rect 12173 17833 12207 17867
rect 14749 17833 14783 17867
rect 15669 17833 15703 17867
rect 23029 17833 23063 17867
rect 28181 17833 28215 17867
rect 22845 17765 22879 17799
rect 25697 17765 25731 17799
rect 15485 17697 15519 17731
rect 18613 17697 18647 17731
rect 18889 17697 18923 17731
rect 22109 17697 22143 17731
rect 22385 17697 22419 17731
rect 23489 17697 23523 17731
rect 27721 17697 27755 17731
rect 29009 17697 29043 17731
rect 30021 17697 30055 17731
rect 8585 17629 8619 17663
rect 10885 17629 10919 17663
rect 11529 17629 11563 17663
rect 12173 17629 12207 17663
rect 12357 17629 12391 17663
rect 12817 17629 12851 17663
rect 15393 17629 15427 17663
rect 16287 17629 16321 17663
rect 16405 17629 16439 17663
rect 16497 17629 16531 17663
rect 16589 17629 16623 17663
rect 19441 17629 19475 17663
rect 19625 17629 19659 17663
rect 19717 17629 19751 17663
rect 19809 17629 19843 17663
rect 23029 17629 23063 17663
rect 23397 17629 23431 17663
rect 24869 17629 24903 17663
rect 24961 17629 24995 17663
rect 25053 17629 25087 17663
rect 25237 17629 25271 17663
rect 26065 17629 26099 17663
rect 26893 17629 26927 17663
rect 27261 17629 27295 17663
rect 28089 17629 28123 17663
rect 29193 17629 29227 17663
rect 30205 17629 30239 17663
rect 30665 17629 30699 17663
rect 30849 17629 30883 17663
rect 10977 17561 11011 17595
rect 13645 17561 13679 17595
rect 14381 17561 14415 17595
rect 14565 17561 14599 17595
rect 15669 17561 15703 17595
rect 25881 17561 25915 17595
rect 26249 17561 26283 17595
rect 26985 17561 27019 17595
rect 27077 17561 27111 17595
rect 9873 17493 9907 17527
rect 10425 17493 10459 17527
rect 11621 17493 11655 17527
rect 13001 17493 13035 17527
rect 13553 17493 13587 17527
rect 15209 17493 15243 17527
rect 16129 17493 16163 17527
rect 17141 17493 17175 17527
rect 20085 17493 20119 17527
rect 20637 17493 20671 17527
rect 24593 17493 24627 17527
rect 25973 17493 26007 17527
rect 26709 17493 26743 17527
rect 27905 17493 27939 17527
rect 31033 17493 31067 17527
rect 9965 17289 9999 17323
rect 14121 17289 14155 17323
rect 14841 17289 14875 17323
rect 16313 17289 16347 17323
rect 17141 17289 17175 17323
rect 21097 17289 21131 17323
rect 27169 17289 27203 17323
rect 28641 17289 28675 17323
rect 30389 17289 30423 17323
rect 12541 17221 12575 17255
rect 13093 17221 13127 17255
rect 13293 17221 13327 17255
rect 13921 17221 13955 17255
rect 20361 17221 20395 17255
rect 21249 17221 21283 17255
rect 21465 17221 21499 17255
rect 23581 17221 23615 17255
rect 28733 17221 28767 17255
rect 29561 17221 29595 17255
rect 30021 17221 30055 17255
rect 31001 17221 31035 17255
rect 31217 17221 31251 17255
rect 29331 17187 29365 17221
rect 10977 17153 11011 17187
rect 11713 17153 11747 17187
rect 12357 17153 12391 17187
rect 12633 17153 12667 17187
rect 14749 17153 14783 17187
rect 15669 17153 15703 17187
rect 15832 17153 15866 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 16865 17153 16899 17187
rect 17141 17153 17175 17187
rect 23857 17153 23891 17187
rect 27537 17153 27571 17187
rect 28457 17153 28491 17187
rect 30205 17153 30239 17187
rect 9413 17085 9447 17119
rect 11805 17085 11839 17119
rect 15117 17085 15151 17119
rect 18153 17085 18187 17119
rect 18383 17085 18417 17119
rect 20637 17085 20671 17119
rect 24317 17085 24351 17119
rect 24593 17085 24627 17119
rect 26065 17085 26099 17119
rect 27445 17085 27479 17119
rect 11069 17017 11103 17051
rect 13461 17017 13495 17051
rect 17049 17017 17083 17051
rect 26525 17017 26559 17051
rect 28273 17017 28307 17051
rect 29193 17017 29227 17051
rect 10517 16949 10551 16983
rect 12357 16949 12391 16983
rect 13277 16949 13311 16983
rect 14105 16949 14139 16983
rect 14289 16949 14323 16983
rect 15025 16949 15059 16983
rect 15209 16949 15243 16983
rect 18889 16949 18923 16983
rect 21281 16949 21315 16983
rect 22109 16949 22143 16983
rect 29377 16949 29411 16983
rect 30849 16949 30883 16983
rect 31033 16949 31067 16983
rect 11069 16745 11103 16779
rect 15301 16745 15335 16779
rect 16681 16745 16715 16779
rect 21189 16745 21223 16779
rect 23949 16745 23983 16779
rect 28917 16745 28951 16779
rect 29929 16745 29963 16779
rect 10425 16677 10459 16711
rect 13001 16677 13035 16711
rect 13737 16677 13771 16711
rect 14565 16677 14599 16711
rect 18889 16677 18923 16711
rect 1593 16609 1627 16643
rect 9965 16609 9999 16643
rect 11621 16609 11655 16643
rect 17417 16609 17451 16643
rect 23121 16609 23155 16643
rect 25697 16609 25731 16643
rect 25881 16609 25915 16643
rect 26065 16609 26099 16643
rect 26157 16609 26191 16643
rect 26709 16609 26743 16643
rect 27261 16609 27295 16643
rect 11529 16541 11563 16575
rect 11707 16541 11741 16575
rect 12357 16541 12391 16575
rect 12817 16541 12851 16575
rect 13001 16541 13035 16575
rect 13461 16541 13495 16575
rect 14289 16541 14323 16575
rect 14381 16541 14415 16575
rect 15025 16541 15059 16575
rect 15301 16541 15335 16575
rect 16037 16541 16071 16575
rect 16221 16541 16255 16575
rect 16313 16541 16347 16575
rect 16405 16541 16439 16575
rect 17141 16541 17175 16575
rect 19441 16541 19475 16575
rect 23397 16541 23431 16575
rect 23857 16541 23891 16575
rect 24869 16541 24903 16575
rect 24961 16541 24995 16575
rect 25053 16541 25087 16575
rect 25237 16541 25271 16575
rect 25973 16541 26007 16575
rect 27077 16541 27111 16575
rect 28181 16541 28215 16575
rect 29009 16541 29043 16575
rect 29101 16541 29135 16575
rect 12265 16473 12299 16507
rect 13737 16473 13771 16507
rect 14565 16473 14599 16507
rect 19717 16473 19751 16507
rect 27905 16473 27939 16507
rect 29897 16473 29931 16507
rect 30113 16473 30147 16507
rect 30757 16473 30791 16507
rect 13553 16405 13587 16439
rect 15577 16405 15611 16439
rect 21649 16405 21683 16439
rect 24593 16405 24627 16439
rect 27077 16405 27111 16439
rect 28733 16405 28767 16439
rect 29745 16405 29779 16439
rect 30665 16405 30699 16439
rect 11069 16201 11103 16235
rect 12173 16201 12207 16235
rect 16313 16201 16347 16235
rect 20545 16201 20579 16235
rect 23765 16201 23799 16235
rect 28273 16201 28307 16235
rect 29285 16201 29319 16235
rect 31217 16201 31251 16235
rect 10609 16133 10643 16167
rect 12725 16133 12759 16167
rect 16957 16133 16991 16167
rect 21465 16133 21499 16167
rect 22293 16133 22327 16167
rect 24501 16133 24535 16167
rect 30021 16133 30055 16167
rect 30573 16133 30607 16167
rect 12633 16065 12667 16099
rect 13277 16065 13311 16099
rect 13461 16065 13495 16099
rect 13921 16065 13955 16099
rect 14197 16065 14231 16099
rect 14841 16065 14875 16099
rect 14933 16065 14967 16099
rect 15025 16065 15059 16099
rect 16037 16065 16071 16099
rect 16154 16065 16188 16099
rect 17785 16065 17819 16099
rect 18153 16065 18187 16099
rect 18245 16065 18279 16099
rect 21005 16065 21039 16099
rect 21097 16065 21131 16099
rect 21281 16065 21315 16099
rect 22017 16065 22051 16099
rect 26433 16065 26467 16099
rect 27169 16065 27203 16099
rect 28089 16065 28123 16099
rect 28181 16065 28215 16099
rect 29101 16065 29135 16099
rect 29745 16065 29779 16099
rect 29837 16065 29871 16099
rect 15669 15997 15703 16031
rect 15945 15997 15979 16031
rect 17141 15997 17175 16031
rect 18797 15997 18831 16031
rect 19073 15997 19107 16031
rect 21373 15997 21407 16031
rect 24225 15997 24259 16031
rect 27353 15997 27387 16031
rect 28457 15997 28491 16031
rect 28917 15997 28951 16031
rect 14105 15929 14139 15963
rect 14197 15929 14231 15963
rect 15209 15929 15243 15963
rect 17601 15929 17635 15963
rect 26525 15929 26559 15963
rect 28181 15929 28215 15963
rect 30757 15929 30791 15963
rect 13369 15861 13403 15895
rect 14657 15861 14691 15895
rect 17877 15861 17911 15895
rect 25973 15861 26007 15895
rect 29745 15861 29779 15895
rect 11345 15657 11379 15691
rect 11805 15657 11839 15691
rect 14841 15657 14875 15691
rect 15301 15657 15335 15691
rect 15485 15657 15519 15691
rect 16497 15657 16531 15691
rect 16681 15657 16715 15691
rect 21189 15657 21223 15691
rect 27905 15657 27939 15691
rect 28089 15657 28123 15691
rect 30573 15657 30607 15691
rect 12357 15589 12391 15623
rect 13645 15589 13679 15623
rect 23949 15589 23983 15623
rect 29929 15589 29963 15623
rect 16405 15521 16439 15555
rect 21925 15521 21959 15555
rect 28549 15521 28583 15555
rect 1593 15453 1627 15487
rect 12909 15453 12943 15487
rect 13553 15453 13587 15487
rect 14749 15453 14783 15487
rect 14841 15453 14875 15487
rect 16129 15453 16163 15487
rect 18889 15453 18923 15487
rect 19441 15453 19475 15487
rect 21649 15453 21683 15487
rect 23857 15453 23891 15487
rect 24593 15453 24627 15487
rect 26985 15453 27019 15487
rect 27169 15453 27203 15487
rect 27261 15453 27295 15487
rect 29745 15453 29779 15487
rect 14565 15385 14599 15419
rect 15669 15385 15703 15419
rect 18613 15385 18647 15419
rect 19717 15385 19751 15419
rect 24869 15385 24903 15419
rect 27721 15385 27755 15419
rect 28733 15385 28767 15419
rect 28917 15385 28951 15419
rect 30665 15385 30699 15419
rect 13001 15317 13035 15351
rect 15469 15317 15503 15351
rect 17141 15317 17175 15351
rect 23397 15317 23431 15351
rect 26341 15317 26375 15351
rect 26801 15317 26835 15351
rect 27931 15317 27965 15351
rect 31217 15317 31251 15351
rect 11989 15113 12023 15147
rect 26525 15113 26559 15147
rect 27537 15113 27571 15147
rect 13001 15045 13035 15079
rect 15117 15045 15151 15079
rect 23489 15045 23523 15079
rect 30849 15045 30883 15079
rect 13829 14977 13863 15011
rect 14473 14977 14507 15011
rect 15301 14977 15335 15011
rect 15393 14977 15427 15011
rect 16957 14977 16991 15011
rect 17601 14977 17635 15011
rect 21189 14977 21223 15011
rect 26433 14977 26467 15011
rect 26617 14977 26651 15011
rect 27353 14977 27387 15011
rect 28089 14977 28123 15011
rect 28825 14977 28859 15011
rect 29653 14977 29687 15011
rect 30297 14977 30331 15011
rect 30757 14977 30791 15011
rect 15853 14909 15887 14943
rect 16313 14909 16347 14943
rect 17693 14909 17727 14943
rect 19901 14909 19935 14943
rect 20177 14909 20211 14943
rect 21465 14909 21499 14943
rect 22017 14909 22051 14943
rect 23765 14909 23799 14943
rect 24225 14909 24259 14943
rect 24501 14909 24535 14943
rect 27169 14909 27203 14943
rect 29561 14909 29595 14943
rect 30205 14909 30239 14943
rect 14565 14841 14599 14875
rect 16037 14841 16071 14875
rect 17969 14841 18003 14875
rect 14013 14773 14047 14807
rect 15117 14773 15151 14807
rect 18429 14773 18463 14807
rect 25973 14773 26007 14807
rect 28089 14773 28123 14807
rect 28917 14773 28951 14807
rect 14657 14569 14691 14603
rect 17325 14569 17359 14603
rect 24593 14569 24627 14603
rect 26801 14569 26835 14603
rect 28825 14569 28859 14603
rect 30481 14569 30515 14603
rect 31309 14569 31343 14603
rect 13645 14501 13679 14535
rect 15945 14501 15979 14535
rect 18889 14501 18923 14535
rect 25145 14501 25179 14535
rect 27721 14501 27755 14535
rect 13093 14433 13127 14467
rect 17601 14433 17635 14467
rect 17693 14433 17727 14467
rect 18429 14433 18463 14467
rect 19993 14433 20027 14467
rect 21925 14433 21959 14467
rect 26157 14433 26191 14467
rect 14473 14365 14507 14399
rect 14657 14365 14691 14399
rect 15117 14365 15151 14399
rect 15761 14365 15795 14399
rect 15945 14365 15979 14399
rect 16405 14365 16439 14399
rect 16681 14365 16715 14399
rect 17509 14365 17543 14399
rect 17785 14365 17819 14399
rect 18521 14365 18555 14399
rect 19441 14365 19475 14399
rect 19717 14365 19751 14399
rect 22201 14365 22235 14399
rect 23213 14365 23247 14399
rect 23489 14365 23523 14399
rect 25605 14365 25639 14399
rect 25973 14365 26007 14399
rect 27445 14365 27479 14399
rect 27537 14365 27571 14399
rect 27721 14365 27755 14399
rect 28181 14365 28215 14399
rect 28365 14365 28399 14399
rect 29009 14365 29043 14399
rect 29745 14365 29779 14399
rect 30665 14365 30699 14399
rect 15209 14297 15243 14331
rect 16497 14297 16531 14331
rect 19809 14297 19843 14331
rect 24961 14297 24995 14331
rect 25881 14297 25915 14331
rect 26785 14297 26819 14331
rect 26985 14297 27019 14331
rect 28273 14297 28307 14331
rect 16865 14229 16899 14263
rect 19625 14229 19659 14263
rect 20453 14229 20487 14263
rect 23949 14229 23983 14263
rect 24777 14229 24811 14263
rect 24869 14229 24903 14263
rect 25789 14229 25823 14263
rect 26617 14229 26651 14263
rect 29837 14229 29871 14263
rect 13829 14025 13863 14059
rect 15577 14025 15611 14059
rect 16221 14025 16255 14059
rect 17141 14025 17175 14059
rect 21097 14025 21131 14059
rect 23765 14025 23799 14059
rect 25447 14025 25481 14059
rect 27905 14025 27939 14059
rect 14381 13957 14415 13991
rect 17233 13957 17267 13991
rect 21249 13957 21283 13991
rect 21465 13957 21499 13991
rect 25237 13957 25271 13991
rect 26065 13957 26099 13991
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 16129 13889 16163 13923
rect 17141 13889 17175 13923
rect 17417 13889 17451 13923
rect 18061 13889 18095 13923
rect 18889 13889 18923 13923
rect 22017 13889 22051 13923
rect 24593 13889 24627 13923
rect 26249 13889 26283 13923
rect 27169 13889 27203 13923
rect 27353 13889 27387 13923
rect 27813 13889 27847 13923
rect 27997 13889 28031 13923
rect 28457 13889 28491 13923
rect 28641 13889 28675 13923
rect 29285 13889 29319 13923
rect 30665 13889 30699 13923
rect 31309 13889 31343 13923
rect 1593 13821 1627 13855
rect 13277 13821 13311 13855
rect 14933 13821 14967 13855
rect 18153 13821 18187 13855
rect 18429 13821 18463 13855
rect 19165 13821 19199 13855
rect 20637 13821 20671 13855
rect 24225 13821 24259 13855
rect 24501 13821 24535 13855
rect 27261 13821 27295 13855
rect 30021 13821 30055 13855
rect 25605 13753 25639 13787
rect 21281 13685 21315 13719
rect 22274 13685 22308 13719
rect 25421 13685 25455 13719
rect 28457 13685 28491 13719
rect 29193 13685 29227 13719
rect 15209 13481 15243 13515
rect 17877 13481 17911 13515
rect 25053 13481 25087 13515
rect 27353 13481 27387 13515
rect 27905 13481 27939 13515
rect 28549 13481 28583 13515
rect 30021 13481 30055 13515
rect 31125 13481 31159 13515
rect 16497 13413 16531 13447
rect 25237 13413 25271 13447
rect 26433 13413 26467 13447
rect 15853 13345 15887 13379
rect 18429 13345 18463 13379
rect 18889 13345 18923 13379
rect 19441 13345 19475 13379
rect 21649 13345 21683 13379
rect 23397 13345 23431 13379
rect 25769 13345 25803 13379
rect 30665 13345 30699 13379
rect 1593 13277 1627 13311
rect 15761 13277 15795 13311
rect 15939 13277 15973 13311
rect 16405 13277 16439 13311
rect 17049 13277 17083 13311
rect 17693 13277 17727 13311
rect 17877 13277 17911 13311
rect 18521 13277 18555 13311
rect 21189 13277 21223 13311
rect 24041 13277 24075 13311
rect 25973 13277 26007 13311
rect 27169 13277 27203 13311
rect 27353 13277 27387 13311
rect 27813 13277 27847 13311
rect 28641 13277 28675 13311
rect 31309 13277 31343 13311
rect 20913 13209 20947 13243
rect 21925 13209 21959 13243
rect 24869 13209 24903 13243
rect 25085 13209 25119 13243
rect 25697 13209 25731 13243
rect 26617 13209 26651 13243
rect 17141 13141 17175 13175
rect 23857 13141 23891 13175
rect 25881 13141 25915 13175
rect 29101 13141 29135 13175
rect 24317 12937 24351 12971
rect 25789 12937 25823 12971
rect 26433 12937 26467 12971
rect 27261 12937 27295 12971
rect 16221 12869 16255 12903
rect 19057 12869 19091 12903
rect 19257 12869 19291 12903
rect 19993 12869 20027 12903
rect 22293 12869 22327 12903
rect 16957 12801 16991 12835
rect 17601 12801 17635 12835
rect 17785 12801 17819 12835
rect 18245 12801 18279 12835
rect 22017 12801 22051 12835
rect 24225 12801 24259 12835
rect 24961 12801 24995 12835
rect 25053 12801 25087 12835
rect 25237 12801 25271 12835
rect 25881 12801 25915 12835
rect 26341 12801 26375 12835
rect 27169 12801 27203 12835
rect 31309 12801 31343 12835
rect 17049 12733 17083 12767
rect 19717 12733 19751 12767
rect 23765 12733 23799 12767
rect 27813 12733 27847 12767
rect 18429 12665 18463 12699
rect 25237 12665 25271 12699
rect 28917 12665 28951 12699
rect 30021 12665 30055 12699
rect 17693 12597 17727 12631
rect 18889 12597 18923 12631
rect 19073 12597 19107 12631
rect 21465 12597 21499 12631
rect 28457 12597 28491 12631
rect 29469 12597 29503 12631
rect 30573 12597 30607 12631
rect 18153 12393 18187 12427
rect 19993 12393 20027 12427
rect 22845 12393 22879 12427
rect 24685 12393 24719 12427
rect 26617 12393 26651 12427
rect 27721 12393 27755 12427
rect 31309 12393 31343 12427
rect 18797 12325 18831 12359
rect 23673 12325 23707 12359
rect 26065 12325 26099 12359
rect 20913 12257 20947 12291
rect 17049 12189 17083 12223
rect 18061 12189 18095 12223
rect 18245 12189 18279 12223
rect 18889 12189 18923 12223
rect 19993 12189 20027 12223
rect 20177 12189 20211 12223
rect 20637 12189 20671 12223
rect 22845 12189 22879 12223
rect 23121 12189 23155 12223
rect 23581 12189 23615 12223
rect 24777 12189 24811 12223
rect 25237 12189 25271 12223
rect 25421 12189 25455 12223
rect 25881 12189 25915 12223
rect 26709 12189 26743 12223
rect 17601 12053 17635 12087
rect 19809 12053 19843 12087
rect 22385 12053 22419 12087
rect 23029 12053 23063 12087
rect 25329 12053 25363 12087
rect 27169 12053 27203 12087
rect 28273 12053 28307 12087
rect 28825 12053 28859 12087
rect 29837 12053 29871 12087
rect 30389 12053 30423 12087
rect 19533 11849 19567 11883
rect 22017 11849 22051 11883
rect 22185 11849 22219 11883
rect 22937 11849 22971 11883
rect 23581 11849 23615 11883
rect 24225 11849 24259 11883
rect 24869 11849 24903 11883
rect 26249 11849 26283 11883
rect 28825 11849 28859 11883
rect 17325 11781 17359 11815
rect 22385 11781 22419 11815
rect 29929 11781 29963 11815
rect 18337 11713 18371 11747
rect 18981 11713 19015 11747
rect 19441 11713 19475 11747
rect 20361 11713 20395 11747
rect 21005 11713 21039 11747
rect 23029 11713 23063 11747
rect 23673 11713 23707 11747
rect 24317 11713 24351 11747
rect 24961 11713 24995 11747
rect 25697 11713 25731 11747
rect 26341 11713 26375 11747
rect 31309 11713 31343 11747
rect 18889 11645 18923 11679
rect 21189 11645 21223 11679
rect 25605 11645 25639 11679
rect 20361 11577 20395 11611
rect 27169 11577 27203 11611
rect 28273 11577 28307 11611
rect 1593 11509 1627 11543
rect 20821 11509 20855 11543
rect 22201 11509 22235 11543
rect 27721 11509 27755 11543
rect 29377 11509 29411 11543
rect 30481 11509 30515 11543
rect 20729 11305 20763 11339
rect 21649 11305 21683 11339
rect 22201 11305 22235 11339
rect 22845 11305 22879 11339
rect 23489 11305 23523 11339
rect 26801 11305 26835 11339
rect 28549 11305 28583 11339
rect 31309 11305 31343 11339
rect 19809 11237 19843 11271
rect 30389 11169 30423 11203
rect 19717 11101 19751 11135
rect 20729 11101 20763 11135
rect 20821 11101 20855 11135
rect 21465 11101 21499 11135
rect 22109 11101 22143 11135
rect 22753 11101 22787 11135
rect 23581 11101 23615 11135
rect 27445 11101 27479 11135
rect 18889 11033 18923 11067
rect 21005 11033 21039 11067
rect 24685 11033 24719 11067
rect 25697 11033 25731 11067
rect 25237 10965 25271 10999
rect 26341 10965 26375 10999
rect 27905 10965 27939 10999
rect 29009 10965 29043 10999
rect 29745 10965 29779 10999
rect 19625 10761 19659 10795
rect 20177 10761 20211 10795
rect 20913 10761 20947 10795
rect 22109 10761 22143 10795
rect 22753 10761 22787 10795
rect 29377 10761 29411 10795
rect 31033 10761 31067 10795
rect 23397 10693 23431 10727
rect 28825 10693 28859 10727
rect 30481 10693 30515 10727
rect 20085 10625 20119 10659
rect 20269 10625 20303 10659
rect 20729 10625 20763 10659
rect 20913 10625 20947 10659
rect 22017 10625 22051 10659
rect 22661 10625 22695 10659
rect 23489 10625 23523 10659
rect 24593 10625 24627 10659
rect 1593 10557 1627 10591
rect 29929 10557 29963 10591
rect 26249 10489 26283 10523
rect 28273 10489 28307 10523
rect 21465 10421 21499 10455
rect 24041 10421 24075 10455
rect 25329 10421 25363 10455
rect 27169 10421 27203 10455
rect 27721 10421 27755 10455
rect 21005 10217 21039 10251
rect 22845 10217 22879 10251
rect 23765 10217 23799 10251
rect 24593 10217 24627 10251
rect 25513 10217 25547 10251
rect 29745 10217 29779 10251
rect 30297 10217 30331 10251
rect 22293 10149 22327 10183
rect 20453 10081 20487 10115
rect 21649 10081 21683 10115
rect 21097 10013 21131 10047
rect 21557 10013 21591 10047
rect 22201 10013 22235 10047
rect 27445 10013 27479 10047
rect 31309 10013 31343 10047
rect 26617 9877 26651 9911
rect 27905 9877 27939 9911
rect 28825 9877 28859 9911
rect 21097 9673 21131 9707
rect 22109 9673 22143 9707
rect 22661 9673 22695 9707
rect 23121 9673 23155 9707
rect 23857 9673 23891 9707
rect 24869 9673 24903 9707
rect 29653 9673 29687 9707
rect 25421 9605 25455 9639
rect 28457 9605 28491 9639
rect 27353 9469 27387 9503
rect 25881 9401 25915 9435
rect 26433 9333 26467 9367
rect 29009 9333 29043 9367
rect 30113 9333 30147 9367
rect 31309 9333 31343 9367
rect 23121 9129 23155 9163
rect 30205 9129 30239 9163
rect 24869 9061 24903 9095
rect 26065 9061 26099 9095
rect 28089 9061 28123 9095
rect 23765 8993 23799 9027
rect 28549 8993 28583 9027
rect 30849 8993 30883 9027
rect 1593 8925 1627 8959
rect 26709 8925 26743 8959
rect 27445 8857 27479 8891
rect 21925 8789 21959 8823
rect 22569 8789 22603 8823
rect 25329 8789 25363 8823
rect 29101 8789 29135 8823
rect 23673 8585 23707 8619
rect 24317 8585 24351 8619
rect 24869 8585 24903 8619
rect 25513 8585 25547 8619
rect 26525 8585 26559 8619
rect 27169 8585 27203 8619
rect 29193 8585 29227 8619
rect 29745 8585 29779 8619
rect 28641 8517 28675 8551
rect 22569 8381 22603 8415
rect 23213 8381 23247 8415
rect 1593 8313 1627 8347
rect 27721 8313 27755 8347
rect 30389 8313 30423 8347
rect 31309 8313 31343 8347
rect 25881 8041 25915 8075
rect 26525 8041 26559 8075
rect 27261 8041 27295 8075
rect 28365 8041 28399 8075
rect 28825 8041 28859 8075
rect 29745 8041 29779 8075
rect 30481 8041 30515 8075
rect 31033 8041 31067 8075
rect 27813 7905 27847 7939
rect 24869 7701 24903 7735
rect 25421 7701 25455 7735
rect 28273 7497 28307 7531
rect 28917 7497 28951 7531
rect 26065 7429 26099 7463
rect 26617 7429 26651 7463
rect 27629 7429 27663 7463
rect 29377 7429 29411 7463
rect 30481 7429 30515 7463
rect 29929 7293 29963 7327
rect 31309 7225 31343 7259
rect 24961 7157 24995 7191
rect 25513 7157 25547 7191
rect 28181 6817 28215 6851
rect 29101 6817 29135 6851
rect 30021 6817 30055 6851
rect 1593 6749 1627 6783
rect 31033 6749 31067 6783
rect 27353 6681 27387 6715
rect 30481 6681 30515 6715
rect 25697 6613 25731 6647
rect 26249 6613 26283 6647
rect 26801 6613 26835 6647
rect 29745 6409 29779 6443
rect 26617 6205 26651 6239
rect 28733 6205 28767 6239
rect 30389 6205 30423 6239
rect 28181 6137 28215 6171
rect 27721 6069 27755 6103
rect 31309 6069 31343 6103
rect 28641 5865 28675 5899
rect 29193 5865 29227 5899
rect 29745 5797 29779 5831
rect 30297 5729 30331 5763
rect 1593 5661 1627 5695
rect 31309 5661 31343 5695
rect 27537 5525 27571 5559
rect 28089 5525 28123 5559
rect 27813 5321 27847 5355
rect 30941 5185 30975 5219
rect 29377 5117 29411 5151
rect 30389 5049 30423 5083
rect 28365 4981 28399 5015
rect 28917 4981 28951 5015
rect 29101 4777 29135 4811
rect 29929 4709 29963 4743
rect 30481 4641 30515 4675
rect 31033 4573 31067 4607
rect 29929 4097 29963 4131
rect 1593 4029 1627 4063
rect 30481 3893 30515 3927
rect 31309 3893 31343 3927
rect 30573 3689 30607 3723
rect 1593 3485 1627 3519
rect 31309 3485 31343 3519
rect 1593 2805 1627 2839
rect 1593 2397 1627 2431
<< metal1 >>
rect 9122 33464 9128 33516
rect 9180 33504 9186 33516
rect 27522 33504 27528 33516
rect 9180 33476 27528 33504
rect 9180 33464 9186 33476
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 10134 33328 10140 33380
rect 10192 33368 10198 33380
rect 24578 33368 24584 33380
rect 10192 33340 24584 33368
rect 10192 33328 10198 33340
rect 24578 33328 24584 33340
rect 24636 33328 24642 33380
rect 12894 33260 12900 33312
rect 12952 33300 12958 33312
rect 27614 33300 27620 33312
rect 12952 33272 27620 33300
rect 12952 33260 12958 33272
rect 27614 33260 27620 33272
rect 27672 33260 27678 33312
rect 13170 33192 13176 33244
rect 13228 33232 13234 33244
rect 25406 33232 25412 33244
rect 13228 33204 25412 33232
rect 13228 33192 13234 33204
rect 25406 33192 25412 33204
rect 25464 33192 25470 33244
rect 12802 33124 12808 33176
rect 12860 33164 12866 33176
rect 25682 33164 25688 33176
rect 12860 33136 25688 33164
rect 12860 33124 12866 33136
rect 25682 33124 25688 33136
rect 25740 33124 25746 33176
rect 10502 32920 10508 32972
rect 10560 32960 10566 32972
rect 22094 32960 22100 32972
rect 10560 32932 22100 32960
rect 10560 32920 10566 32932
rect 22094 32920 22100 32932
rect 22152 32920 22158 32972
rect 13630 32784 13636 32836
rect 13688 32824 13694 32836
rect 18230 32824 18236 32836
rect 13688 32796 18236 32824
rect 13688 32784 13694 32796
rect 18230 32784 18236 32796
rect 18288 32784 18294 32836
rect 19886 32784 19892 32836
rect 19944 32824 19950 32836
rect 25222 32824 25228 32836
rect 19944 32796 25228 32824
rect 19944 32784 19950 32796
rect 25222 32784 25228 32796
rect 25280 32784 25286 32836
rect 9582 32716 9588 32768
rect 9640 32756 9646 32768
rect 21634 32756 21640 32768
rect 9640 32728 21640 32756
rect 9640 32716 9646 32728
rect 21634 32716 21640 32728
rect 21692 32716 21698 32768
rect 1104 32666 31992 32688
rect 1104 32614 8632 32666
rect 8684 32614 8696 32666
rect 8748 32614 8760 32666
rect 8812 32614 8824 32666
rect 8876 32614 8888 32666
rect 8940 32614 16314 32666
rect 16366 32614 16378 32666
rect 16430 32614 16442 32666
rect 16494 32614 16506 32666
rect 16558 32614 16570 32666
rect 16622 32614 23996 32666
rect 24048 32614 24060 32666
rect 24112 32614 24124 32666
rect 24176 32614 24188 32666
rect 24240 32614 24252 32666
rect 24304 32614 31678 32666
rect 31730 32614 31742 32666
rect 31794 32614 31806 32666
rect 31858 32614 31870 32666
rect 31922 32614 31934 32666
rect 31986 32614 31992 32666
rect 1104 32592 31992 32614
rect 18230 32552 18236 32564
rect 18191 32524 18236 32552
rect 18230 32512 18236 32524
rect 18288 32552 18294 32564
rect 18785 32555 18843 32561
rect 18785 32552 18797 32555
rect 18288 32524 18797 32552
rect 18288 32512 18294 32524
rect 18785 32521 18797 32524
rect 18831 32552 18843 32555
rect 21266 32552 21272 32564
rect 18831 32524 21272 32552
rect 18831 32521 18843 32524
rect 18785 32515 18843 32521
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 24578 32552 24584 32564
rect 24539 32524 24584 32552
rect 24578 32512 24584 32524
rect 24636 32512 24642 32564
rect 21450 32484 21456 32496
rect 21363 32456 21456 32484
rect 21450 32444 21456 32456
rect 21508 32484 21514 32496
rect 24854 32484 24860 32496
rect 21508 32456 24860 32484
rect 21508 32444 21514 32456
rect 24854 32444 24860 32456
rect 24912 32444 24918 32496
rect 25130 32444 25136 32496
rect 25188 32484 25194 32496
rect 28166 32484 28172 32496
rect 25188 32456 28172 32484
rect 25188 32444 25194 32456
rect 28166 32444 28172 32456
rect 28224 32444 28230 32496
rect 934 32376 940 32428
rect 992 32416 998 32428
rect 1581 32419 1639 32425
rect 1581 32416 1593 32419
rect 992 32388 1593 32416
rect 992 32376 998 32388
rect 1581 32385 1593 32388
rect 1627 32385 1639 32419
rect 2222 32416 2228 32428
rect 2183 32388 2228 32416
rect 1581 32379 1639 32385
rect 2222 32376 2228 32388
rect 2280 32376 2286 32428
rect 2866 32416 2872 32428
rect 2827 32388 2872 32416
rect 2866 32376 2872 32388
rect 2924 32376 2930 32428
rect 4614 32416 4620 32428
rect 4575 32388 4620 32416
rect 4614 32376 4620 32388
rect 4672 32376 4678 32428
rect 5810 32416 5816 32428
rect 5771 32388 5816 32416
rect 5810 32376 5816 32388
rect 5868 32376 5874 32428
rect 8202 32416 8208 32428
rect 8163 32388 8208 32416
rect 8202 32376 8208 32388
rect 8260 32376 8266 32428
rect 9398 32416 9404 32428
rect 9359 32388 9404 32416
rect 9398 32376 9404 32388
rect 9456 32376 9462 32428
rect 11790 32416 11796 32428
rect 11751 32388 11796 32416
rect 11790 32376 11796 32388
rect 11848 32376 11854 32428
rect 12986 32416 12992 32428
rect 12947 32388 12992 32416
rect 12986 32376 12992 32388
rect 13044 32376 13050 32428
rect 15378 32416 15384 32428
rect 15339 32388 15384 32416
rect 15378 32376 15384 32388
rect 15436 32376 15442 32428
rect 16666 32376 16672 32428
rect 16724 32416 16730 32428
rect 16853 32419 16911 32425
rect 16853 32416 16865 32419
rect 16724 32388 16865 32416
rect 16724 32376 16730 32388
rect 16853 32385 16865 32388
rect 16899 32385 16911 32419
rect 16853 32379 16911 32385
rect 18874 32376 18880 32428
rect 18932 32416 18938 32428
rect 19429 32419 19487 32425
rect 19429 32416 19441 32419
rect 18932 32388 19441 32416
rect 18932 32376 18938 32388
rect 19429 32385 19441 32388
rect 19475 32385 19487 32419
rect 19429 32379 19487 32385
rect 20070 32376 20076 32428
rect 20128 32416 20134 32428
rect 20165 32419 20223 32425
rect 20165 32416 20177 32419
rect 20128 32388 20177 32416
rect 20128 32376 20134 32388
rect 20165 32385 20177 32388
rect 20211 32385 20223 32419
rect 20165 32379 20223 32385
rect 22462 32376 22468 32428
rect 22520 32416 22526 32428
rect 22557 32419 22615 32425
rect 22557 32416 22569 32419
rect 22520 32388 22569 32416
rect 22520 32376 22526 32388
rect 22557 32385 22569 32388
rect 22603 32385 22615 32419
rect 22557 32379 22615 32385
rect 23658 32376 23664 32428
rect 23716 32416 23722 32428
rect 23753 32419 23811 32425
rect 23753 32416 23765 32419
rect 23716 32388 23765 32416
rect 23716 32376 23722 32388
rect 23753 32385 23765 32388
rect 23799 32385 23811 32419
rect 23753 32379 23811 32385
rect 23842 32376 23848 32428
rect 23900 32416 23906 32428
rect 25314 32416 25320 32428
rect 23900 32388 25320 32416
rect 23900 32376 23906 32388
rect 25314 32376 25320 32388
rect 25372 32376 25378 32428
rect 26050 32376 26056 32428
rect 26108 32416 26114 32428
rect 26145 32419 26203 32425
rect 26145 32416 26157 32419
rect 26108 32388 26157 32416
rect 26108 32376 26114 32388
rect 26145 32385 26157 32388
rect 26191 32385 26203 32419
rect 26145 32379 26203 32385
rect 27246 32376 27252 32428
rect 27304 32416 27310 32428
rect 27341 32419 27399 32425
rect 27341 32416 27353 32419
rect 27304 32388 27353 32416
rect 27304 32376 27310 32388
rect 27341 32385 27353 32388
rect 27387 32385 27399 32419
rect 27341 32379 27399 32385
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 29733 32419 29791 32425
rect 29733 32416 29745 32419
rect 29696 32388 29745 32416
rect 29696 32376 29702 32388
rect 29733 32385 29745 32388
rect 29779 32385 29791 32419
rect 30926 32416 30932 32428
rect 30887 32388 30932 32416
rect 29733 32379 29791 32385
rect 30926 32376 30932 32388
rect 30984 32376 30990 32428
rect 13538 32308 13544 32360
rect 13596 32348 13602 32360
rect 20622 32348 20628 32360
rect 13596 32320 20628 32348
rect 13596 32308 13602 32320
rect 20622 32308 20628 32320
rect 20680 32308 20686 32360
rect 21174 32308 21180 32360
rect 21232 32348 21238 32360
rect 26510 32348 26516 32360
rect 21232 32320 26516 32348
rect 21232 32308 21238 32320
rect 26510 32308 26516 32320
rect 26568 32308 26574 32360
rect 27522 32308 27528 32360
rect 27580 32348 27586 32360
rect 32214 32348 32220 32360
rect 27580 32320 32220 32348
rect 27580 32308 27586 32320
rect 32214 32308 32220 32320
rect 32272 32308 32278 32360
rect 11606 32240 11612 32292
rect 11664 32280 11670 32292
rect 14826 32280 14832 32292
rect 11664 32252 14832 32280
rect 11664 32240 11670 32252
rect 14826 32240 14832 32252
rect 14884 32240 14890 32292
rect 14918 32240 14924 32292
rect 14976 32280 14982 32292
rect 16942 32280 16948 32292
rect 14976 32252 16948 32280
rect 14976 32240 14982 32252
rect 16942 32240 16948 32252
rect 17000 32240 17006 32292
rect 19058 32240 19064 32292
rect 19116 32280 19122 32292
rect 20809 32283 20867 32289
rect 20809 32280 20821 32283
rect 19116 32252 20821 32280
rect 19116 32240 19122 32252
rect 20809 32249 20821 32252
rect 20855 32280 20867 32283
rect 21542 32280 21548 32292
rect 20855 32252 21548 32280
rect 20855 32249 20867 32252
rect 20809 32243 20867 32249
rect 21542 32240 21548 32252
rect 21600 32240 21606 32292
rect 23106 32240 23112 32292
rect 23164 32280 23170 32292
rect 26878 32280 26884 32292
rect 23164 32252 26884 32280
rect 23164 32240 23170 32252
rect 26878 32240 26884 32252
rect 26936 32240 26942 32292
rect 28350 32280 28356 32292
rect 28311 32252 28356 32280
rect 28350 32240 28356 32252
rect 28408 32240 28414 32292
rect 12342 32172 12348 32224
rect 12400 32212 12406 32224
rect 12437 32215 12495 32221
rect 12437 32212 12449 32215
rect 12400 32184 12449 32212
rect 12400 32172 12406 32184
rect 12437 32181 12449 32184
rect 12483 32181 12495 32215
rect 12437 32175 12495 32181
rect 13078 32172 13084 32224
rect 13136 32212 13142 32224
rect 13633 32215 13691 32221
rect 13633 32212 13645 32215
rect 13136 32184 13645 32212
rect 13136 32172 13142 32184
rect 13633 32181 13645 32184
rect 13679 32181 13691 32215
rect 13633 32175 13691 32181
rect 14369 32215 14427 32221
rect 14369 32181 14381 32215
rect 14415 32212 14427 32215
rect 15102 32212 15108 32224
rect 14415 32184 15108 32212
rect 14415 32181 14427 32184
rect 14369 32175 14427 32181
rect 15102 32172 15108 32184
rect 15160 32172 15166 32224
rect 16022 32172 16028 32224
rect 16080 32212 16086 32224
rect 16209 32215 16267 32221
rect 16209 32212 16221 32215
rect 16080 32184 16221 32212
rect 16080 32172 16086 32184
rect 16209 32181 16221 32184
rect 16255 32181 16267 32215
rect 17770 32212 17776 32224
rect 17731 32184 17776 32212
rect 16209 32175 16267 32181
rect 17770 32172 17776 32184
rect 17828 32172 17834 32224
rect 18782 32172 18788 32224
rect 18840 32212 18846 32224
rect 21082 32212 21088 32224
rect 18840 32184 21088 32212
rect 18840 32172 18846 32184
rect 21082 32172 21088 32184
rect 21140 32212 21146 32224
rect 22005 32215 22063 32221
rect 22005 32212 22017 32215
rect 21140 32184 22017 32212
rect 21140 32172 21146 32184
rect 22005 32181 22017 32184
rect 22051 32181 22063 32215
rect 22005 32175 22063 32181
rect 22370 32172 22376 32224
rect 22428 32212 22434 32224
rect 23290 32212 23296 32224
rect 22428 32184 23296 32212
rect 22428 32172 22434 32184
rect 23290 32172 23296 32184
rect 23348 32172 23354 32224
rect 23566 32172 23572 32224
rect 23624 32212 23630 32224
rect 25038 32212 25044 32224
rect 23624 32184 25044 32212
rect 23624 32172 23630 32184
rect 25038 32172 25044 32184
rect 25096 32172 25102 32224
rect 25222 32172 25228 32224
rect 25280 32212 25286 32224
rect 28905 32215 28963 32221
rect 28905 32212 28917 32215
rect 25280 32184 28917 32212
rect 25280 32172 25286 32184
rect 28905 32181 28917 32184
rect 28951 32212 28963 32215
rect 30282 32212 30288 32224
rect 28951 32184 30288 32212
rect 28951 32181 28963 32184
rect 28905 32175 28963 32181
rect 30282 32172 30288 32184
rect 30340 32172 30346 32224
rect 30469 32215 30527 32221
rect 30469 32181 30481 32215
rect 30515 32212 30527 32215
rect 30834 32212 30840 32224
rect 30515 32184 30840 32212
rect 30515 32181 30527 32184
rect 30469 32175 30527 32181
rect 30834 32172 30840 32184
rect 30892 32172 30898 32224
rect 1104 32122 31832 32144
rect 1104 32070 4791 32122
rect 4843 32070 4855 32122
rect 4907 32070 4919 32122
rect 4971 32070 4983 32122
rect 5035 32070 5047 32122
rect 5099 32070 12473 32122
rect 12525 32070 12537 32122
rect 12589 32070 12601 32122
rect 12653 32070 12665 32122
rect 12717 32070 12729 32122
rect 12781 32070 20155 32122
rect 20207 32070 20219 32122
rect 20271 32070 20283 32122
rect 20335 32070 20347 32122
rect 20399 32070 20411 32122
rect 20463 32070 27837 32122
rect 27889 32070 27901 32122
rect 27953 32070 27965 32122
rect 28017 32070 28029 32122
rect 28081 32070 28093 32122
rect 28145 32070 31832 32122
rect 1104 32048 31832 32070
rect 1578 32008 1584 32020
rect 1539 31980 1584 32008
rect 1578 31968 1584 31980
rect 1636 31968 1642 32020
rect 14826 31968 14832 32020
rect 14884 32008 14890 32020
rect 15473 32011 15531 32017
rect 15473 32008 15485 32011
rect 14884 31980 15485 32008
rect 14884 31968 14890 31980
rect 15473 31977 15485 31980
rect 15519 31977 15531 32011
rect 15473 31971 15531 31977
rect 18230 31968 18236 32020
rect 18288 32008 18294 32020
rect 18782 32008 18788 32020
rect 18288 31980 18788 32008
rect 18288 31968 18294 31980
rect 18782 31968 18788 31980
rect 18840 31968 18846 32020
rect 19886 32008 19892 32020
rect 19847 31980 19892 32008
rect 19886 31968 19892 31980
rect 19944 31968 19950 32020
rect 19978 31968 19984 32020
rect 20036 32008 20042 32020
rect 21174 32008 21180 32020
rect 20036 31980 20668 32008
rect 21135 31980 21180 32008
rect 20036 31968 20042 31980
rect 11882 31900 11888 31952
rect 11940 31940 11946 31952
rect 20070 31940 20076 31952
rect 11940 31912 20076 31940
rect 11940 31900 11946 31912
rect 20070 31900 20076 31912
rect 20128 31900 20134 31952
rect 20640 31949 20668 31980
rect 21174 31968 21180 31980
rect 21232 31968 21238 32020
rect 22005 32011 22063 32017
rect 22005 31977 22017 32011
rect 22051 32008 22063 32011
rect 22738 32008 22744 32020
rect 22051 31980 22744 32008
rect 22051 31977 22063 31980
rect 22005 31971 22063 31977
rect 22738 31968 22744 31980
rect 22796 31968 22802 32020
rect 23106 32008 23112 32020
rect 23067 31980 23112 32008
rect 23106 31968 23112 31980
rect 23164 31968 23170 32020
rect 23842 32008 23848 32020
rect 23803 31980 23848 32008
rect 23842 31968 23848 31980
rect 23900 31968 23906 32020
rect 24486 31968 24492 32020
rect 24544 32008 24550 32020
rect 24673 32011 24731 32017
rect 24673 32008 24685 32011
rect 24544 31980 24685 32008
rect 24544 31968 24550 31980
rect 24673 31977 24685 31980
rect 24719 31977 24731 32011
rect 25222 32008 25228 32020
rect 25183 31980 25228 32008
rect 24673 31971 24731 31977
rect 25222 31968 25228 31980
rect 25280 31968 25286 32020
rect 26326 32008 26332 32020
rect 25792 31980 26332 32008
rect 20625 31943 20683 31949
rect 20625 31909 20637 31943
rect 20671 31940 20683 31943
rect 22557 31943 22615 31949
rect 22557 31940 22569 31943
rect 20671 31912 22569 31940
rect 20671 31909 20683 31912
rect 20625 31903 20683 31909
rect 22557 31909 22569 31912
rect 22603 31940 22615 31943
rect 24578 31940 24584 31952
rect 22603 31912 24584 31940
rect 22603 31909 22615 31912
rect 22557 31903 22615 31909
rect 24578 31900 24584 31912
rect 24636 31900 24642 31952
rect 24762 31900 24768 31952
rect 24820 31940 24826 31952
rect 25792 31940 25820 31980
rect 26326 31968 26332 31980
rect 26384 31968 26390 32020
rect 26510 32008 26516 32020
rect 26471 31980 26516 32008
rect 26510 31968 26516 31980
rect 26568 32008 26574 32020
rect 27522 32008 27528 32020
rect 26568 31980 27528 32008
rect 26568 31968 26574 31980
rect 27522 31968 27528 31980
rect 27580 32008 27586 32020
rect 28169 32011 28227 32017
rect 28169 32008 28181 32011
rect 27580 31980 28181 32008
rect 27580 31968 27586 31980
rect 28169 31977 28181 31980
rect 28215 31977 28227 32011
rect 30558 32008 30564 32020
rect 30519 31980 30564 32008
rect 28169 31971 28227 31977
rect 30558 31968 30564 31980
rect 30616 31968 30622 32020
rect 24820 31912 25820 31940
rect 25869 31943 25927 31949
rect 24820 31900 24826 31912
rect 25869 31909 25881 31943
rect 25915 31940 25927 31943
rect 29270 31940 29276 31952
rect 25915 31912 29276 31940
rect 25915 31909 25927 31912
rect 25869 31903 25927 31909
rect 29270 31900 29276 31912
rect 29328 31900 29334 31952
rect 31202 31940 31208 31952
rect 31163 31912 31208 31940
rect 31202 31900 31208 31912
rect 31260 31900 31266 31952
rect 13725 31875 13783 31881
rect 13725 31841 13737 31875
rect 13771 31872 13783 31875
rect 15930 31872 15936 31884
rect 13771 31844 15936 31872
rect 13771 31841 13783 31844
rect 13725 31835 13783 31841
rect 15930 31832 15936 31844
rect 15988 31872 15994 31884
rect 24394 31872 24400 31884
rect 15988 31844 24400 31872
rect 15988 31832 15994 31844
rect 24394 31832 24400 31844
rect 24452 31832 24458 31884
rect 27617 31875 27675 31881
rect 27617 31872 27629 31875
rect 24504 31844 27629 31872
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31804 12127 31807
rect 14734 31804 14740 31816
rect 12115 31776 14740 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 14734 31764 14740 31776
rect 14792 31764 14798 31816
rect 15013 31807 15071 31813
rect 15013 31773 15025 31807
rect 15059 31804 15071 31807
rect 15838 31804 15844 31816
rect 15059 31776 15844 31804
rect 15059 31773 15071 31776
rect 15013 31767 15071 31773
rect 15838 31764 15844 31776
rect 15896 31764 15902 31816
rect 16666 31804 16672 31816
rect 16579 31776 16672 31804
rect 16666 31764 16672 31776
rect 16724 31804 16730 31816
rect 20806 31804 20812 31816
rect 16724 31776 20812 31804
rect 16724 31764 16730 31776
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 21174 31764 21180 31816
rect 21232 31804 21238 31816
rect 24504 31804 24532 31844
rect 21232 31776 24532 31804
rect 24581 31807 24639 31813
rect 21232 31764 21238 31776
rect 24581 31773 24593 31807
rect 24627 31804 24639 31807
rect 24670 31804 24676 31816
rect 24627 31776 24676 31804
rect 24627 31773 24639 31776
rect 24581 31767 24639 31773
rect 10318 31696 10324 31748
rect 10376 31736 10382 31748
rect 14458 31736 14464 31748
rect 10376 31708 14464 31736
rect 10376 31696 10382 31708
rect 14458 31696 14464 31708
rect 14516 31696 14522 31748
rect 15654 31696 15660 31748
rect 15712 31736 15718 31748
rect 17681 31739 17739 31745
rect 17681 31736 17693 31739
rect 15712 31708 17693 31736
rect 15712 31696 15718 31708
rect 17681 31705 17693 31708
rect 17727 31705 17739 31739
rect 17681 31699 17739 31705
rect 18322 31696 18328 31748
rect 18380 31736 18386 31748
rect 24596 31736 24624 31767
rect 24670 31764 24676 31776
rect 24728 31764 24734 31816
rect 24762 31764 24768 31816
rect 24820 31804 24826 31816
rect 25240 31813 25268 31844
rect 27617 31841 27629 31844
rect 27663 31841 27675 31875
rect 27617 31835 27675 31841
rect 27706 31832 27712 31884
rect 27764 31872 27770 31884
rect 32490 31872 32496 31884
rect 27764 31844 32496 31872
rect 27764 31832 27770 31844
rect 32490 31832 32496 31844
rect 32548 31832 32554 31884
rect 25225 31807 25283 31813
rect 24820 31776 24865 31804
rect 24820 31764 24826 31776
rect 25225 31773 25237 31807
rect 25271 31773 25283 31807
rect 25225 31767 25283 31773
rect 25409 31807 25467 31813
rect 25409 31773 25421 31807
rect 25455 31773 25467 31807
rect 25409 31767 25467 31773
rect 18380 31708 24624 31736
rect 18380 31696 18386 31708
rect 11514 31668 11520 31680
rect 11475 31640 11520 31668
rect 11514 31628 11520 31640
rect 11572 31668 11578 31680
rect 12342 31668 12348 31680
rect 11572 31640 12348 31668
rect 11572 31628 11578 31640
rect 12342 31628 12348 31640
rect 12400 31668 12406 31680
rect 12529 31671 12587 31677
rect 12529 31668 12541 31671
rect 12400 31640 12541 31668
rect 12400 31628 12406 31640
rect 12529 31637 12541 31640
rect 12575 31637 12587 31671
rect 12529 31631 12587 31637
rect 13173 31671 13231 31677
rect 13173 31637 13185 31671
rect 13219 31668 13231 31671
rect 14642 31668 14648 31680
rect 13219 31640 14648 31668
rect 13219 31637 13231 31640
rect 13173 31631 13231 31637
rect 14642 31628 14648 31640
rect 14700 31628 14706 31680
rect 16117 31671 16175 31677
rect 16117 31637 16129 31671
rect 16163 31668 16175 31671
rect 16206 31668 16212 31680
rect 16163 31640 16212 31668
rect 16163 31637 16175 31640
rect 16117 31631 16175 31637
rect 16206 31628 16212 31640
rect 16264 31628 16270 31680
rect 17221 31671 17279 31677
rect 17221 31637 17233 31671
rect 17267 31668 17279 31671
rect 17402 31668 17408 31680
rect 17267 31640 17408 31668
rect 17267 31637 17279 31640
rect 17221 31631 17279 31637
rect 17402 31628 17408 31640
rect 17460 31628 17466 31680
rect 18233 31671 18291 31677
rect 18233 31637 18245 31671
rect 18279 31668 18291 31671
rect 19886 31668 19892 31680
rect 18279 31640 19892 31668
rect 18279 31637 18291 31640
rect 18233 31631 18291 31637
rect 19886 31628 19892 31640
rect 19944 31628 19950 31680
rect 21818 31628 21824 31680
rect 21876 31668 21882 31680
rect 23106 31668 23112 31680
rect 21876 31640 23112 31668
rect 21876 31628 21882 31640
rect 23106 31628 23112 31640
rect 23164 31628 23170 31680
rect 23842 31628 23848 31680
rect 23900 31668 23906 31680
rect 25424 31668 25452 31767
rect 25774 31764 25780 31816
rect 25832 31804 25838 31816
rect 25869 31807 25927 31813
rect 25869 31804 25881 31807
rect 25832 31776 25881 31804
rect 25832 31764 25838 31776
rect 25869 31773 25881 31776
rect 25915 31773 25927 31807
rect 25869 31767 25927 31773
rect 26053 31807 26111 31813
rect 26053 31773 26065 31807
rect 26099 31804 26111 31807
rect 26142 31804 26148 31816
rect 26099 31776 26148 31804
rect 26099 31773 26111 31776
rect 26053 31767 26111 31773
rect 26142 31764 26148 31776
rect 26200 31764 26206 31816
rect 29730 31804 29736 31816
rect 29691 31776 29736 31804
rect 29730 31764 29736 31776
rect 29788 31764 29794 31816
rect 29822 31764 29828 31816
rect 29880 31804 29886 31816
rect 31021 31807 31079 31813
rect 31021 31804 31033 31807
rect 29880 31776 31033 31804
rect 29880 31764 29886 31776
rect 31021 31773 31033 31776
rect 31067 31773 31079 31807
rect 31021 31767 31079 31773
rect 26970 31696 26976 31748
rect 27028 31736 27034 31748
rect 27065 31739 27123 31745
rect 27065 31736 27077 31739
rect 27028 31708 27077 31736
rect 27028 31696 27034 31708
rect 27065 31705 27077 31708
rect 27111 31705 27123 31739
rect 27065 31699 27123 31705
rect 27706 31696 27712 31748
rect 27764 31736 27770 31748
rect 28718 31736 28724 31748
rect 27764 31708 28724 31736
rect 27764 31696 27770 31708
rect 28718 31696 28724 31708
rect 28776 31696 28782 31748
rect 28810 31668 28816 31680
rect 23900 31640 28816 31668
rect 23900 31628 23906 31640
rect 28810 31628 28816 31640
rect 28868 31628 28874 31680
rect 1104 31578 31992 31600
rect 1104 31526 8632 31578
rect 8684 31526 8696 31578
rect 8748 31526 8760 31578
rect 8812 31526 8824 31578
rect 8876 31526 8888 31578
rect 8940 31526 16314 31578
rect 16366 31526 16378 31578
rect 16430 31526 16442 31578
rect 16494 31526 16506 31578
rect 16558 31526 16570 31578
rect 16622 31526 23996 31578
rect 24048 31526 24060 31578
rect 24112 31526 24124 31578
rect 24176 31526 24188 31578
rect 24240 31526 24252 31578
rect 24304 31526 31678 31578
rect 31730 31526 31742 31578
rect 31794 31526 31806 31578
rect 31858 31526 31870 31578
rect 31922 31526 31934 31578
rect 31986 31526 31992 31578
rect 1104 31504 31992 31526
rect 15197 31467 15255 31473
rect 15197 31433 15209 31467
rect 15243 31464 15255 31467
rect 16758 31464 16764 31476
rect 15243 31436 16764 31464
rect 15243 31433 15255 31436
rect 15197 31427 15255 31433
rect 16758 31424 16764 31436
rect 16816 31424 16822 31476
rect 16942 31424 16948 31476
rect 17000 31464 17006 31476
rect 18417 31467 18475 31473
rect 18417 31464 18429 31467
rect 17000 31436 18429 31464
rect 17000 31424 17006 31436
rect 18417 31433 18429 31436
rect 18463 31464 18475 31467
rect 19150 31464 19156 31476
rect 18463 31436 19156 31464
rect 18463 31433 18475 31436
rect 18417 31427 18475 31433
rect 19150 31424 19156 31436
rect 19208 31464 19214 31476
rect 21450 31464 21456 31476
rect 19208 31436 21456 31464
rect 19208 31424 19214 31436
rect 21450 31424 21456 31436
rect 21508 31424 21514 31476
rect 22738 31424 22744 31476
rect 22796 31464 22802 31476
rect 23750 31464 23756 31476
rect 22796 31436 23756 31464
rect 22796 31424 22802 31436
rect 23750 31424 23756 31436
rect 23808 31424 23814 31476
rect 23842 31424 23848 31476
rect 23900 31464 23906 31476
rect 24486 31464 24492 31476
rect 23900 31436 24492 31464
rect 23900 31424 23906 31436
rect 24486 31424 24492 31436
rect 24544 31424 24550 31476
rect 24578 31424 24584 31476
rect 24636 31464 24642 31476
rect 24949 31467 25007 31473
rect 24949 31464 24961 31467
rect 24636 31436 24961 31464
rect 24636 31424 24642 31436
rect 24949 31433 24961 31436
rect 24995 31464 25007 31467
rect 28258 31464 28264 31476
rect 24995 31436 28264 31464
rect 24995 31433 25007 31436
rect 24949 31427 25007 31433
rect 28258 31424 28264 31436
rect 28316 31424 28322 31476
rect 14734 31356 14740 31408
rect 14792 31396 14798 31408
rect 17034 31396 17040 31408
rect 14792 31368 17040 31396
rect 14792 31356 14798 31368
rect 17034 31356 17040 31368
rect 17092 31396 17098 31408
rect 21174 31396 21180 31408
rect 17092 31368 21180 31396
rect 17092 31356 17098 31368
rect 21174 31356 21180 31368
rect 21232 31356 21238 31408
rect 22094 31356 22100 31408
rect 22152 31396 22158 31408
rect 27709 31399 27767 31405
rect 27709 31396 27721 31399
rect 22152 31368 27721 31396
rect 22152 31356 22158 31368
rect 27709 31365 27721 31368
rect 27755 31365 27767 31399
rect 27709 31359 27767 31365
rect 13538 31328 13544 31340
rect 13499 31300 13544 31328
rect 13538 31288 13544 31300
rect 13596 31288 13602 31340
rect 14826 31288 14832 31340
rect 14884 31328 14890 31340
rect 14884 31300 16574 31328
rect 14884 31288 14890 31300
rect 16546 31260 16574 31300
rect 18414 31288 18420 31340
rect 18472 31328 18478 31340
rect 19061 31331 19119 31337
rect 19061 31328 19073 31331
rect 18472 31300 19073 31328
rect 18472 31288 18478 31300
rect 19061 31297 19073 31300
rect 19107 31328 19119 31331
rect 20530 31328 20536 31340
rect 19107 31300 20536 31328
rect 19107 31297 19119 31300
rect 19061 31291 19119 31297
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 23477 31331 23535 31337
rect 23477 31297 23489 31331
rect 23523 31328 23535 31331
rect 23566 31328 23572 31340
rect 23523 31300 23572 31328
rect 23523 31297 23535 31300
rect 23477 31291 23535 31297
rect 22094 31260 22100 31272
rect 16546 31232 22100 31260
rect 22094 31220 22100 31232
rect 22152 31220 22158 31272
rect 22186 31220 22192 31272
rect 22244 31260 22250 31272
rect 23492 31260 23520 31291
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 23750 31288 23756 31340
rect 23808 31328 23814 31340
rect 24121 31331 24179 31337
rect 24121 31328 24133 31331
rect 23808 31300 24133 31328
rect 23808 31288 23814 31300
rect 24121 31297 24133 31300
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 24305 31331 24363 31337
rect 24305 31297 24317 31331
rect 24351 31328 24363 31331
rect 24486 31328 24492 31340
rect 24351 31300 24492 31328
rect 24351 31297 24363 31300
rect 24305 31291 24363 31297
rect 24486 31288 24492 31300
rect 24544 31288 24550 31340
rect 25133 31331 25191 31337
rect 25133 31328 25145 31331
rect 24826 31300 25145 31328
rect 22244 31232 23520 31260
rect 22244 31220 22250 31232
rect 23658 31220 23664 31272
rect 23716 31260 23722 31272
rect 23842 31260 23848 31272
rect 23716 31232 23848 31260
rect 23716 31220 23722 31232
rect 23842 31220 23848 31232
rect 23900 31220 23906 31272
rect 11885 31195 11943 31201
rect 11885 31161 11897 31195
rect 11931 31192 11943 31195
rect 12342 31192 12348 31204
rect 11931 31164 12348 31192
rect 11931 31161 11943 31164
rect 11885 31155 11943 31161
rect 12342 31152 12348 31164
rect 12400 31152 12406 31204
rect 16206 31152 16212 31204
rect 16264 31192 16270 31204
rect 16301 31195 16359 31201
rect 16301 31192 16313 31195
rect 16264 31164 16313 31192
rect 16264 31152 16270 31164
rect 16301 31161 16313 31164
rect 16347 31192 16359 31195
rect 17865 31195 17923 31201
rect 17865 31192 17877 31195
rect 16347 31164 17877 31192
rect 16347 31161 16359 31164
rect 16301 31155 16359 31161
rect 17865 31161 17877 31164
rect 17911 31192 17923 31195
rect 18046 31192 18052 31204
rect 17911 31164 18052 31192
rect 17911 31161 17923 31164
rect 17865 31155 17923 31161
rect 18046 31152 18052 31164
rect 18104 31152 18110 31204
rect 18138 31152 18144 31204
rect 18196 31192 18202 31204
rect 22370 31192 22376 31204
rect 18196 31164 22376 31192
rect 18196 31152 18202 31164
rect 22370 31152 22376 31164
rect 22428 31152 22434 31204
rect 22462 31152 22468 31204
rect 22520 31192 22526 31204
rect 24826 31192 24854 31300
rect 25133 31297 25145 31300
rect 25179 31297 25191 31331
rect 25133 31291 25191 31297
rect 25777 31331 25835 31337
rect 25777 31297 25789 31331
rect 25823 31328 25835 31331
rect 25866 31328 25872 31340
rect 25823 31300 25872 31328
rect 25823 31297 25835 31300
rect 25777 31291 25835 31297
rect 25148 31260 25176 31291
rect 25866 31288 25872 31300
rect 25924 31288 25930 31340
rect 26142 31288 26148 31340
rect 26200 31328 26206 31340
rect 26237 31331 26295 31337
rect 26237 31328 26249 31331
rect 26200 31300 26249 31328
rect 26200 31288 26206 31300
rect 26237 31297 26249 31300
rect 26283 31297 26295 31331
rect 26237 31291 26295 31297
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31328 26387 31331
rect 27154 31328 27160 31340
rect 26375 31300 27160 31328
rect 26375 31297 26387 31300
rect 26329 31291 26387 31297
rect 27154 31288 27160 31300
rect 27212 31328 27218 31340
rect 30742 31328 30748 31340
rect 27212 31300 30748 31328
rect 27212 31288 27218 31300
rect 30742 31288 30748 31300
rect 30800 31288 30806 31340
rect 26694 31260 26700 31272
rect 25148 31232 26700 31260
rect 26694 31220 26700 31232
rect 26752 31220 26758 31272
rect 32122 31260 32128 31272
rect 26804 31232 32128 31260
rect 22520 31164 24854 31192
rect 22520 31152 22526 31164
rect 25038 31152 25044 31204
rect 25096 31192 25102 31204
rect 26602 31192 26608 31204
rect 25096 31164 26608 31192
rect 25096 31152 25102 31164
rect 26602 31152 26608 31164
rect 26660 31152 26666 31204
rect 1578 31124 1584 31136
rect 1539 31096 1584 31124
rect 1578 31084 1584 31096
rect 1636 31084 1642 31136
rect 10502 31124 10508 31136
rect 10463 31096 10508 31124
rect 10502 31084 10508 31096
rect 10560 31084 10566 31136
rect 11149 31127 11207 31133
rect 11149 31093 11161 31127
rect 11195 31124 11207 31127
rect 11790 31124 11796 31136
rect 11195 31096 11796 31124
rect 11195 31093 11207 31096
rect 11149 31087 11207 31093
rect 11790 31084 11796 31096
rect 11848 31084 11854 31136
rect 12158 31084 12164 31136
rect 12216 31124 12222 31136
rect 12437 31127 12495 31133
rect 12437 31124 12449 31127
rect 12216 31096 12449 31124
rect 12216 31084 12222 31096
rect 12437 31093 12449 31096
rect 12483 31093 12495 31127
rect 12437 31087 12495 31093
rect 12802 31084 12808 31136
rect 12860 31124 12866 31136
rect 12897 31127 12955 31133
rect 12897 31124 12909 31127
rect 12860 31096 12909 31124
rect 12860 31084 12866 31096
rect 12897 31093 12909 31096
rect 12943 31093 12955 31127
rect 13998 31124 14004 31136
rect 13959 31096 14004 31124
rect 12897 31087 12955 31093
rect 13998 31084 14004 31096
rect 14056 31084 14062 31136
rect 14645 31127 14703 31133
rect 14645 31093 14657 31127
rect 14691 31124 14703 31127
rect 14734 31124 14740 31136
rect 14691 31096 14740 31124
rect 14691 31093 14703 31096
rect 14645 31087 14703 31093
rect 14734 31084 14740 31096
rect 14792 31084 14798 31136
rect 15562 31084 15568 31136
rect 15620 31124 15626 31136
rect 15657 31127 15715 31133
rect 15657 31124 15669 31127
rect 15620 31096 15669 31124
rect 15620 31084 15626 31096
rect 15657 31093 15669 31096
rect 15703 31093 15715 31127
rect 15657 31087 15715 31093
rect 17218 31084 17224 31136
rect 17276 31124 17282 31136
rect 17313 31127 17371 31133
rect 17313 31124 17325 31127
rect 17276 31096 17325 31124
rect 17276 31084 17282 31096
rect 17313 31093 17325 31096
rect 17359 31093 17371 31127
rect 17313 31087 17371 31093
rect 17770 31084 17776 31136
rect 17828 31124 17834 31136
rect 18966 31124 18972 31136
rect 17828 31096 18972 31124
rect 17828 31084 17834 31096
rect 18966 31084 18972 31096
rect 19024 31124 19030 31136
rect 19705 31127 19763 31133
rect 19705 31124 19717 31127
rect 19024 31096 19717 31124
rect 19024 31084 19030 31096
rect 19705 31093 19717 31096
rect 19751 31093 19763 31127
rect 19705 31087 19763 31093
rect 19794 31084 19800 31136
rect 19852 31124 19858 31136
rect 20625 31127 20683 31133
rect 20625 31124 20637 31127
rect 19852 31096 20637 31124
rect 19852 31084 19858 31096
rect 20625 31093 20637 31096
rect 20671 31093 20683 31127
rect 20625 31087 20683 31093
rect 22002 31084 22008 31136
rect 22060 31124 22066 31136
rect 22833 31127 22891 31133
rect 22833 31124 22845 31127
rect 22060 31096 22845 31124
rect 22060 31084 22066 31096
rect 22833 31093 22845 31096
rect 22879 31093 22891 31127
rect 22833 31087 22891 31093
rect 23569 31127 23627 31133
rect 23569 31093 23581 31127
rect 23615 31124 23627 31127
rect 23750 31124 23756 31136
rect 23615 31096 23756 31124
rect 23615 31093 23627 31096
rect 23569 31087 23627 31093
rect 23750 31084 23756 31096
rect 23808 31084 23814 31136
rect 23842 31084 23848 31136
rect 23900 31124 23906 31136
rect 24302 31124 24308 31136
rect 23900 31096 24308 31124
rect 23900 31084 23906 31096
rect 24302 31084 24308 31096
rect 24360 31084 24366 31136
rect 24578 31084 24584 31136
rect 24636 31124 24642 31136
rect 24762 31124 24768 31136
rect 24636 31096 24768 31124
rect 24636 31084 24642 31096
rect 24762 31084 24768 31096
rect 24820 31084 24826 31136
rect 24854 31084 24860 31136
rect 24912 31124 24918 31136
rect 25498 31124 25504 31136
rect 24912 31096 25504 31124
rect 24912 31084 24918 31096
rect 25498 31084 25504 31096
rect 25556 31084 25562 31136
rect 25685 31127 25743 31133
rect 25685 31093 25697 31127
rect 25731 31124 25743 31127
rect 26804 31124 26832 31232
rect 32122 31220 32128 31232
rect 32180 31220 32186 31272
rect 26878 31152 26884 31204
rect 26936 31192 26942 31204
rect 28813 31195 28871 31201
rect 28813 31192 28825 31195
rect 26936 31164 28825 31192
rect 26936 31152 26942 31164
rect 28813 31161 28825 31164
rect 28859 31161 28871 31195
rect 28813 31155 28871 31161
rect 27246 31124 27252 31136
rect 25731 31096 26832 31124
rect 27207 31096 27252 31124
rect 25731 31093 25743 31096
rect 25685 31087 25743 31093
rect 27246 31084 27252 31096
rect 27304 31084 27310 31136
rect 27338 31084 27344 31136
rect 27396 31124 27402 31136
rect 29362 31124 29368 31136
rect 27396 31096 29368 31124
rect 27396 31084 27402 31096
rect 29362 31084 29368 31096
rect 29420 31084 29426 31136
rect 30006 31124 30012 31136
rect 29967 31096 30012 31124
rect 30006 31084 30012 31096
rect 30064 31084 30070 31136
rect 30650 31124 30656 31136
rect 30611 31096 30656 31124
rect 30650 31084 30656 31096
rect 30708 31084 30714 31136
rect 31297 31127 31355 31133
rect 31297 31093 31309 31127
rect 31343 31124 31355 31127
rect 32030 31124 32036 31136
rect 31343 31096 32036 31124
rect 31343 31093 31355 31096
rect 31297 31087 31355 31093
rect 32030 31084 32036 31096
rect 32088 31084 32094 31136
rect 1104 31034 31832 31056
rect 1104 30982 4791 31034
rect 4843 30982 4855 31034
rect 4907 30982 4919 31034
rect 4971 30982 4983 31034
rect 5035 30982 5047 31034
rect 5099 30982 12473 31034
rect 12525 30982 12537 31034
rect 12589 30982 12601 31034
rect 12653 30982 12665 31034
rect 12717 30982 12729 31034
rect 12781 30982 20155 31034
rect 20207 30982 20219 31034
rect 20271 30982 20283 31034
rect 20335 30982 20347 31034
rect 20399 30982 20411 31034
rect 20463 30982 27837 31034
rect 27889 30982 27901 31034
rect 27953 30982 27965 31034
rect 28017 30982 28029 31034
rect 28081 30982 28093 31034
rect 28145 30982 31832 31034
rect 1104 30960 31832 30982
rect 9030 30880 9036 30932
rect 9088 30920 9094 30932
rect 10318 30920 10324 30932
rect 9088 30892 10324 30920
rect 9088 30880 9094 30892
rect 10318 30880 10324 30892
rect 10376 30880 10382 30932
rect 13998 30920 14004 30932
rect 10520 30892 14004 30920
rect 4062 30812 4068 30864
rect 4120 30852 4126 30864
rect 10520 30852 10548 30892
rect 13998 30880 14004 30892
rect 14056 30880 14062 30932
rect 16114 30920 16120 30932
rect 16075 30892 16120 30920
rect 16114 30880 16120 30892
rect 16172 30880 16178 30932
rect 17218 30880 17224 30932
rect 17276 30920 17282 30932
rect 17678 30920 17684 30932
rect 17276 30892 17684 30920
rect 17276 30880 17282 30892
rect 17678 30880 17684 30892
rect 17736 30880 17742 30932
rect 18322 30920 18328 30932
rect 18283 30892 18328 30920
rect 18322 30880 18328 30892
rect 18380 30880 18386 30932
rect 18690 30880 18696 30932
rect 18748 30920 18754 30932
rect 18785 30923 18843 30929
rect 18785 30920 18797 30923
rect 18748 30892 18797 30920
rect 18748 30880 18754 30892
rect 18785 30889 18797 30892
rect 18831 30889 18843 30923
rect 18785 30883 18843 30889
rect 19334 30880 19340 30932
rect 19392 30920 19398 30932
rect 21821 30923 21879 30929
rect 21821 30920 21833 30923
rect 19392 30892 21833 30920
rect 19392 30880 19398 30892
rect 21821 30889 21833 30892
rect 21867 30889 21879 30923
rect 21821 30883 21879 30889
rect 23014 30880 23020 30932
rect 23072 30920 23078 30932
rect 24578 30920 24584 30932
rect 23072 30892 24584 30920
rect 23072 30880 23078 30892
rect 24578 30880 24584 30892
rect 24636 30880 24642 30932
rect 24762 30920 24768 30932
rect 24723 30892 24768 30920
rect 24762 30880 24768 30892
rect 24820 30880 24826 30932
rect 24946 30920 24952 30932
rect 24907 30892 24952 30920
rect 24946 30880 24952 30892
rect 25004 30880 25010 30932
rect 25222 30880 25228 30932
rect 25280 30920 25286 30932
rect 25593 30923 25651 30929
rect 25593 30920 25605 30923
rect 25280 30892 25605 30920
rect 25280 30880 25286 30892
rect 25593 30889 25605 30892
rect 25639 30889 25651 30923
rect 28718 30920 28724 30932
rect 25593 30883 25651 30889
rect 26436 30892 28724 30920
rect 4120 30824 10548 30852
rect 4120 30812 4126 30824
rect 11882 30812 11888 30864
rect 11940 30852 11946 30864
rect 21358 30852 21364 30864
rect 11940 30824 21364 30852
rect 11940 30812 11946 30824
rect 21358 30812 21364 30824
rect 21416 30812 21422 30864
rect 21450 30812 21456 30864
rect 21508 30852 21514 30864
rect 21508 30824 23152 30852
rect 21508 30812 21514 30824
rect 11422 30784 11428 30796
rect 11383 30756 11428 30784
rect 11422 30744 11428 30756
rect 11480 30744 11486 30796
rect 11790 30744 11796 30796
rect 11848 30784 11854 30796
rect 13078 30784 13084 30796
rect 11848 30756 13084 30784
rect 11848 30744 11854 30756
rect 13078 30744 13084 30756
rect 13136 30784 13142 30796
rect 13173 30787 13231 30793
rect 13173 30784 13185 30787
rect 13136 30756 13185 30784
rect 13136 30744 13142 30756
rect 13173 30753 13185 30756
rect 13219 30784 13231 30787
rect 13219 30756 17254 30784
rect 13219 30753 13231 30756
rect 13173 30747 13231 30753
rect 11054 30676 11060 30728
rect 11112 30716 11118 30728
rect 11514 30716 11520 30728
rect 11112 30688 11520 30716
rect 11112 30676 11118 30688
rect 11514 30676 11520 30688
rect 11572 30716 11578 30728
rect 11977 30719 12035 30725
rect 11977 30716 11989 30719
rect 11572 30688 11989 30716
rect 11572 30676 11578 30688
rect 11977 30685 11989 30688
rect 12023 30716 12035 30719
rect 12066 30716 12072 30728
rect 12023 30688 12072 30716
rect 12023 30685 12035 30688
rect 11977 30679 12035 30685
rect 12066 30676 12072 30688
rect 12124 30676 12130 30728
rect 12250 30676 12256 30728
rect 12308 30716 12314 30728
rect 13725 30719 13783 30725
rect 13725 30716 13737 30719
rect 12308 30688 13737 30716
rect 12308 30676 12314 30688
rect 13725 30685 13737 30688
rect 13771 30716 13783 30719
rect 14461 30719 14519 30725
rect 14461 30716 14473 30719
rect 13771 30688 14473 30716
rect 13771 30685 13783 30688
rect 13725 30679 13783 30685
rect 14461 30685 14473 30688
rect 14507 30716 14519 30719
rect 15562 30716 15568 30728
rect 14507 30688 15568 30716
rect 14507 30685 14519 30688
rect 14461 30679 14519 30685
rect 15562 30676 15568 30688
rect 15620 30676 15626 30728
rect 9861 30651 9919 30657
rect 9861 30617 9873 30651
rect 9907 30648 9919 30651
rect 13354 30648 13360 30660
rect 9907 30620 13360 30648
rect 9907 30617 9919 30620
rect 9861 30611 9919 30617
rect 13354 30608 13360 30620
rect 13412 30608 13418 30660
rect 17126 30648 17132 30660
rect 17087 30620 17132 30648
rect 17126 30608 17132 30620
rect 17184 30608 17190 30660
rect 17226 30648 17254 30756
rect 17494 30744 17500 30796
rect 17552 30784 17558 30796
rect 17552 30756 22508 30784
rect 17552 30744 17558 30756
rect 17862 30676 17868 30728
rect 17920 30716 17926 30728
rect 22370 30716 22376 30728
rect 17920 30688 22376 30716
rect 17920 30676 17926 30688
rect 22370 30676 22376 30688
rect 22428 30676 22434 30728
rect 22480 30725 22508 30756
rect 22465 30719 22523 30725
rect 22465 30685 22477 30719
rect 22511 30685 22523 30719
rect 22465 30679 22523 30685
rect 22649 30719 22707 30725
rect 22649 30685 22661 30719
rect 22695 30716 22707 30719
rect 22830 30716 22836 30728
rect 22695 30688 22836 30716
rect 22695 30685 22707 30688
rect 22649 30679 22707 30685
rect 22830 30676 22836 30688
rect 22888 30676 22894 30728
rect 23124 30725 23152 30824
rect 23198 30812 23204 30864
rect 23256 30852 23262 30864
rect 26234 30852 26240 30864
rect 23256 30824 26240 30852
rect 23256 30812 23262 30824
rect 26234 30812 26240 30824
rect 26292 30812 26298 30864
rect 26436 30861 26464 30892
rect 28718 30880 28724 30892
rect 28776 30880 28782 30932
rect 28810 30880 28816 30932
rect 28868 30920 28874 30932
rect 28868 30892 28913 30920
rect 28868 30880 28874 30892
rect 26421 30855 26479 30861
rect 26421 30821 26433 30855
rect 26467 30821 26479 30855
rect 26421 30815 26479 30821
rect 26513 30855 26571 30861
rect 26513 30821 26525 30855
rect 26559 30852 26571 30855
rect 29730 30852 29736 30864
rect 26559 30824 29736 30852
rect 26559 30821 26571 30824
rect 26513 30815 26571 30821
rect 29730 30812 29736 30824
rect 29788 30812 29794 30864
rect 23382 30744 23388 30796
rect 23440 30784 23446 30796
rect 27065 30787 27123 30793
rect 23440 30756 25652 30784
rect 23440 30744 23446 30756
rect 23109 30719 23167 30725
rect 23109 30685 23121 30719
rect 23155 30685 23167 30719
rect 23290 30716 23296 30728
rect 23251 30688 23296 30716
rect 23109 30679 23167 30685
rect 23290 30676 23296 30688
rect 23348 30676 23354 30728
rect 23566 30676 23572 30728
rect 23624 30716 23630 30728
rect 23753 30719 23811 30725
rect 23753 30716 23765 30719
rect 23624 30688 23765 30716
rect 23624 30676 23630 30688
rect 23753 30685 23765 30688
rect 23799 30685 23811 30719
rect 23753 30679 23811 30685
rect 24320 30716 24532 30718
rect 24320 30690 25452 30716
rect 18046 30648 18052 30660
rect 17226 30620 18052 30648
rect 18046 30608 18052 30620
rect 18104 30648 18110 30660
rect 18104 30620 21036 30648
rect 18104 30608 18110 30620
rect 10965 30583 11023 30589
rect 10965 30549 10977 30583
rect 11011 30580 11023 30583
rect 11238 30580 11244 30592
rect 11011 30552 11244 30580
rect 11011 30549 11023 30552
rect 10965 30543 11023 30549
rect 11238 30540 11244 30552
rect 11296 30540 11302 30592
rect 12342 30540 12348 30592
rect 12400 30580 12406 30592
rect 12529 30583 12587 30589
rect 12529 30580 12541 30583
rect 12400 30552 12541 30580
rect 12400 30540 12406 30552
rect 12529 30549 12541 30552
rect 12575 30549 12587 30583
rect 12529 30543 12587 30549
rect 14642 30540 14648 30592
rect 14700 30580 14706 30592
rect 14921 30583 14979 30589
rect 14921 30580 14933 30583
rect 14700 30552 14933 30580
rect 14700 30540 14706 30552
rect 14921 30549 14933 30552
rect 14967 30549 14979 30583
rect 14921 30543 14979 30549
rect 15565 30583 15623 30589
rect 15565 30549 15577 30583
rect 15611 30580 15623 30583
rect 15654 30580 15660 30592
rect 15611 30552 15660 30580
rect 15611 30549 15623 30552
rect 15565 30543 15623 30549
rect 15654 30540 15660 30552
rect 15712 30540 15718 30592
rect 15746 30540 15752 30592
rect 15804 30580 15810 30592
rect 16577 30583 16635 30589
rect 16577 30580 16589 30583
rect 15804 30552 16589 30580
rect 15804 30540 15810 30552
rect 16577 30549 16589 30552
rect 16623 30549 16635 30583
rect 16577 30543 16635 30549
rect 17678 30540 17684 30592
rect 17736 30580 17742 30592
rect 18966 30580 18972 30592
rect 17736 30552 18972 30580
rect 17736 30540 17742 30552
rect 18966 30540 18972 30552
rect 19024 30540 19030 30592
rect 19518 30580 19524 30592
rect 19479 30552 19524 30580
rect 19518 30540 19524 30552
rect 19576 30540 19582 30592
rect 20346 30580 20352 30592
rect 20307 30552 20352 30580
rect 20346 30540 20352 30552
rect 20404 30540 20410 30592
rect 20898 30580 20904 30592
rect 20859 30552 20904 30580
rect 20898 30540 20904 30552
rect 20956 30540 20962 30592
rect 21008 30580 21036 30620
rect 21726 30608 21732 30660
rect 21784 30648 21790 30660
rect 22557 30651 22615 30657
rect 22557 30648 22569 30651
rect 21784 30620 22569 30648
rect 21784 30608 21790 30620
rect 22557 30617 22569 30620
rect 22603 30617 22615 30651
rect 22557 30611 22615 30617
rect 22922 30608 22928 30660
rect 22980 30648 22986 30660
rect 24320 30648 24348 30690
rect 24504 30688 25452 30690
rect 22980 30620 24348 30648
rect 22980 30608 22986 30620
rect 24486 30608 24492 30660
rect 24544 30648 24550 30660
rect 24581 30651 24639 30657
rect 24581 30648 24593 30651
rect 24544 30620 24593 30648
rect 24544 30608 24550 30620
rect 24581 30617 24593 30620
rect 24627 30617 24639 30651
rect 24581 30611 24639 30617
rect 24670 30608 24676 30660
rect 24728 30648 24734 30660
rect 25424 30657 25452 30688
rect 25624 30657 25652 30756
rect 27065 30753 27077 30787
rect 27111 30784 27123 30787
rect 28442 30784 28448 30796
rect 27111 30756 28448 30784
rect 27111 30753 27123 30756
rect 27065 30747 27123 30753
rect 28442 30744 28448 30756
rect 28500 30744 28506 30796
rect 26513 30719 26571 30725
rect 26513 30716 26525 30719
rect 25700 30688 26525 30716
rect 24781 30651 24839 30657
rect 24781 30648 24793 30651
rect 24728 30620 24793 30648
rect 24728 30608 24734 30620
rect 24781 30617 24793 30620
rect 24827 30617 24839 30651
rect 24781 30611 24839 30617
rect 25409 30651 25467 30657
rect 25409 30617 25421 30651
rect 25455 30617 25467 30651
rect 25409 30611 25467 30617
rect 25609 30651 25667 30657
rect 25609 30617 25621 30651
rect 25655 30617 25667 30651
rect 25609 30611 25667 30617
rect 23014 30580 23020 30592
rect 21008 30552 23020 30580
rect 23014 30540 23020 30552
rect 23072 30540 23078 30592
rect 23201 30583 23259 30589
rect 23201 30549 23213 30583
rect 23247 30580 23259 30583
rect 23842 30580 23848 30592
rect 23247 30552 23848 30580
rect 23247 30549 23259 30552
rect 23201 30543 23259 30549
rect 23842 30540 23848 30552
rect 23900 30540 23906 30592
rect 23937 30583 23995 30589
rect 23937 30549 23949 30583
rect 23983 30580 23995 30583
rect 25222 30580 25228 30592
rect 23983 30552 25228 30580
rect 23983 30549 23995 30552
rect 23937 30543 23995 30549
rect 25222 30540 25228 30552
rect 25280 30540 25286 30592
rect 25498 30540 25504 30592
rect 25556 30580 25562 30592
rect 25700 30580 25728 30688
rect 26513 30685 26525 30688
rect 26559 30685 26571 30719
rect 26513 30679 26571 30685
rect 26602 30676 26608 30728
rect 26660 30716 26666 30728
rect 26973 30719 27031 30725
rect 26973 30716 26985 30719
rect 26660 30688 26985 30716
rect 26660 30676 26666 30688
rect 26973 30685 26985 30688
rect 27019 30685 27031 30719
rect 26973 30679 27031 30685
rect 26237 30651 26295 30657
rect 26237 30617 26249 30651
rect 26283 30648 26295 30651
rect 26418 30648 26424 30660
rect 26283 30620 26424 30648
rect 26283 30617 26295 30620
rect 26237 30611 26295 30617
rect 26418 30608 26424 30620
rect 26476 30608 26482 30660
rect 25556 30552 25728 30580
rect 25777 30583 25835 30589
rect 25556 30540 25562 30552
rect 25777 30549 25789 30583
rect 25823 30580 25835 30583
rect 25958 30580 25964 30592
rect 25823 30552 25964 30580
rect 25823 30549 25835 30552
rect 25777 30543 25835 30549
rect 25958 30540 25964 30552
rect 26016 30540 26022 30592
rect 26988 30580 27016 30679
rect 27430 30676 27436 30728
rect 27488 30716 27494 30728
rect 27617 30719 27675 30725
rect 27617 30716 27629 30719
rect 27488 30688 27629 30716
rect 27488 30676 27494 30688
rect 27617 30685 27629 30688
rect 27663 30685 27675 30719
rect 27617 30679 27675 30685
rect 27801 30719 27859 30725
rect 27801 30685 27813 30719
rect 27847 30716 27859 30719
rect 28166 30716 28172 30728
rect 27847 30688 28172 30716
rect 27847 30685 27859 30688
rect 27801 30679 27859 30685
rect 28166 30676 28172 30688
rect 28224 30676 28230 30728
rect 28350 30716 28356 30728
rect 28311 30688 28356 30716
rect 28350 30676 28356 30688
rect 28408 30676 28414 30728
rect 29917 30719 29975 30725
rect 29917 30685 29929 30719
rect 29963 30716 29975 30719
rect 30466 30716 30472 30728
rect 29963 30688 30472 30716
rect 29963 30685 29975 30688
rect 29917 30679 29975 30685
rect 30466 30676 30472 30688
rect 30524 30676 30530 30728
rect 31297 30719 31355 30725
rect 31297 30685 31309 30719
rect 31343 30716 31355 30719
rect 31570 30716 31576 30728
rect 31343 30688 31576 30716
rect 31343 30685 31355 30688
rect 31297 30679 31355 30685
rect 31570 30676 31576 30688
rect 31628 30676 31634 30728
rect 27709 30651 27767 30657
rect 27709 30617 27721 30651
rect 27755 30648 27767 30651
rect 28902 30648 28908 30660
rect 27755 30620 28908 30648
rect 27755 30617 27767 30620
rect 27709 30611 27767 30617
rect 28902 30608 28908 30620
rect 28960 30608 28966 30660
rect 28994 30580 29000 30592
rect 26988 30552 29000 30580
rect 28994 30540 29000 30552
rect 29052 30540 29058 30592
rect 30098 30580 30104 30592
rect 30059 30552 30104 30580
rect 30098 30540 30104 30552
rect 30156 30540 30162 30592
rect 30558 30580 30564 30592
rect 30519 30552 30564 30580
rect 30558 30540 30564 30552
rect 30616 30540 30622 30592
rect 1104 30490 31992 30512
rect 1104 30438 8632 30490
rect 8684 30438 8696 30490
rect 8748 30438 8760 30490
rect 8812 30438 8824 30490
rect 8876 30438 8888 30490
rect 8940 30438 16314 30490
rect 16366 30438 16378 30490
rect 16430 30438 16442 30490
rect 16494 30438 16506 30490
rect 16558 30438 16570 30490
rect 16622 30438 23996 30490
rect 24048 30438 24060 30490
rect 24112 30438 24124 30490
rect 24176 30438 24188 30490
rect 24240 30438 24252 30490
rect 24304 30438 31678 30490
rect 31730 30438 31742 30490
rect 31794 30438 31806 30490
rect 31858 30438 31870 30490
rect 31922 30438 31934 30490
rect 31986 30438 31992 30490
rect 1104 30416 31992 30438
rect 2682 30336 2688 30388
rect 2740 30376 2746 30388
rect 10042 30376 10048 30388
rect 2740 30348 10048 30376
rect 2740 30336 2746 30348
rect 8941 30311 8999 30317
rect 8941 30277 8953 30311
rect 8987 30308 8999 30311
rect 9030 30308 9036 30320
rect 8987 30280 9036 30308
rect 8987 30277 8999 30280
rect 8941 30271 8999 30277
rect 9030 30268 9036 30280
rect 9088 30268 9094 30320
rect 9968 30317 9996 30348
rect 10042 30336 10048 30348
rect 10100 30336 10106 30388
rect 11146 30336 11152 30388
rect 11204 30376 11210 30388
rect 14642 30376 14648 30388
rect 11204 30348 14648 30376
rect 11204 30336 11210 30348
rect 14642 30336 14648 30348
rect 14700 30336 14706 30388
rect 14918 30336 14924 30388
rect 14976 30376 14982 30388
rect 17773 30379 17831 30385
rect 17773 30376 17785 30379
rect 14976 30348 17785 30376
rect 14976 30336 14982 30348
rect 17773 30345 17785 30348
rect 17819 30376 17831 30379
rect 19242 30376 19248 30388
rect 17819 30348 19248 30376
rect 17819 30345 17831 30348
rect 17773 30339 17831 30345
rect 19242 30336 19248 30348
rect 19300 30336 19306 30388
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 19484 30348 21128 30376
rect 19484 30336 19490 30348
rect 9953 30311 10011 30317
rect 9953 30277 9965 30311
rect 9999 30277 10011 30311
rect 9953 30271 10011 30277
rect 10597 30311 10655 30317
rect 10597 30277 10609 30311
rect 10643 30308 10655 30311
rect 12342 30308 12348 30320
rect 10643 30280 12348 30308
rect 10643 30277 10655 30280
rect 10597 30271 10655 30277
rect 9858 30200 9864 30252
rect 9916 30240 9922 30252
rect 10612 30240 10640 30271
rect 12342 30268 12348 30280
rect 12400 30268 12406 30320
rect 13541 30311 13599 30317
rect 13541 30277 13553 30311
rect 13587 30308 13599 30311
rect 13630 30308 13636 30320
rect 13587 30280 13636 30308
rect 13587 30277 13599 30280
rect 13541 30271 13599 30277
rect 13630 30268 13636 30280
rect 13688 30268 13694 30320
rect 16114 30268 16120 30320
rect 16172 30308 16178 30320
rect 16301 30311 16359 30317
rect 16301 30308 16313 30311
rect 16172 30280 16313 30308
rect 16172 30268 16178 30280
rect 16301 30277 16313 30280
rect 16347 30308 16359 30311
rect 19334 30308 19340 30320
rect 16347 30280 19340 30308
rect 16347 30277 16359 30280
rect 16301 30271 16359 30277
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 19705 30311 19763 30317
rect 19705 30277 19717 30311
rect 19751 30308 19763 30311
rect 19794 30308 19800 30320
rect 19751 30280 19800 30308
rect 19751 30277 19763 30280
rect 19705 30271 19763 30277
rect 19794 30268 19800 30280
rect 19852 30268 19858 30320
rect 20438 30308 20444 30320
rect 20399 30280 20444 30308
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 20622 30268 20628 30320
rect 20680 30308 20686 30320
rect 20993 30311 21051 30317
rect 20993 30308 21005 30311
rect 20680 30280 21005 30308
rect 20680 30268 20686 30280
rect 20993 30277 21005 30280
rect 21039 30277 21051 30311
rect 21100 30308 21128 30348
rect 21358 30336 21364 30388
rect 21416 30376 21422 30388
rect 23106 30376 23112 30388
rect 21416 30348 23112 30376
rect 21416 30336 21422 30348
rect 23106 30336 23112 30348
rect 23164 30336 23170 30388
rect 23829 30379 23887 30385
rect 23829 30376 23841 30379
rect 23296 30348 23841 30376
rect 21100 30280 22610 30308
rect 20993 30271 21051 30277
rect 9916 30212 10640 30240
rect 9916 30200 9922 30212
rect 12066 30200 12072 30252
rect 12124 30240 12130 30252
rect 14645 30243 14703 30249
rect 14645 30240 14657 30243
rect 12124 30212 14657 30240
rect 12124 30200 12130 30212
rect 14645 30209 14657 30212
rect 14691 30240 14703 30243
rect 18322 30240 18328 30252
rect 14691 30212 18328 30240
rect 14691 30209 14703 30212
rect 14645 30203 14703 30209
rect 18322 30200 18328 30212
rect 18380 30200 18386 30252
rect 18598 30200 18604 30252
rect 18656 30240 18662 30252
rect 22281 30243 22339 30249
rect 22281 30240 22293 30243
rect 18656 30212 22293 30240
rect 18656 30200 18662 30212
rect 22281 30209 22293 30212
rect 22327 30209 22339 30243
rect 22281 30203 22339 30209
rect 22370 30200 22376 30252
rect 22428 30240 22434 30252
rect 22465 30243 22523 30249
rect 22465 30240 22477 30243
rect 22428 30212 22477 30240
rect 22428 30200 22434 30212
rect 22465 30209 22477 30212
rect 22511 30209 22523 30243
rect 22582 30240 22610 30280
rect 22646 30268 22652 30320
rect 22704 30308 22710 30320
rect 23017 30311 23075 30317
rect 23017 30308 23029 30311
rect 22704 30280 23029 30308
rect 22704 30268 22710 30280
rect 23017 30277 23029 30280
rect 23063 30277 23075 30311
rect 23198 30308 23204 30320
rect 23159 30280 23204 30308
rect 23017 30271 23075 30277
rect 23198 30268 23204 30280
rect 23256 30268 23262 30320
rect 22922 30240 22928 30252
rect 22582 30212 22928 30240
rect 22465 30203 22523 30209
rect 22922 30200 22928 30212
rect 22980 30200 22986 30252
rect 23296 30240 23324 30348
rect 23829 30345 23841 30348
rect 23875 30376 23887 30379
rect 24699 30379 24757 30385
rect 23875 30348 24616 30376
rect 23875 30345 23887 30348
rect 23829 30339 23887 30345
rect 24029 30311 24087 30317
rect 24029 30277 24041 30311
rect 24075 30308 24087 30311
rect 24210 30308 24216 30320
rect 24075 30280 24216 30308
rect 24075 30277 24087 30280
rect 23032 30212 23324 30240
rect 23750 30224 23756 30276
rect 23808 30240 23814 30276
rect 24029 30271 24087 30277
rect 24210 30268 24216 30280
rect 24268 30268 24274 30320
rect 24489 30311 24547 30317
rect 24489 30277 24501 30311
rect 24535 30277 24547 30311
rect 24588 30308 24616 30348
rect 24699 30345 24711 30379
rect 24745 30376 24757 30379
rect 24946 30376 24952 30388
rect 24745 30348 24952 30376
rect 24745 30345 24757 30348
rect 24699 30339 24757 30345
rect 24946 30336 24952 30348
rect 25004 30336 25010 30388
rect 25038 30336 25044 30388
rect 25096 30376 25102 30388
rect 25314 30376 25320 30388
rect 25096 30348 25320 30376
rect 25096 30336 25102 30348
rect 25314 30336 25320 30348
rect 25372 30336 25378 30388
rect 25498 30336 25504 30388
rect 25556 30376 25562 30388
rect 25866 30376 25872 30388
rect 25556 30348 25872 30376
rect 25556 30336 25562 30348
rect 25866 30336 25872 30348
rect 25924 30336 25930 30388
rect 26234 30336 26240 30388
rect 26292 30376 26298 30388
rect 26878 30376 26884 30388
rect 26292 30348 26884 30376
rect 26292 30336 26298 30348
rect 26878 30336 26884 30348
rect 26936 30336 26942 30388
rect 27982 30376 27988 30388
rect 26977 30348 27988 30376
rect 26421 30311 26479 30317
rect 24588 30280 26353 30308
rect 24489 30271 24547 30277
rect 24504 30240 24532 30271
rect 24670 30240 24676 30252
rect 23808 30224 23872 30240
rect 23768 30212 23872 30224
rect 24504 30212 24676 30240
rect 23032 30184 23060 30212
rect 1578 30172 1584 30184
rect 1539 30144 1584 30172
rect 1578 30132 1584 30144
rect 1636 30132 1642 30184
rect 11149 30175 11207 30181
rect 11149 30141 11161 30175
rect 11195 30172 11207 30175
rect 14090 30172 14096 30184
rect 11195 30144 14096 30172
rect 11195 30141 11207 30144
rect 11149 30135 11207 30141
rect 14090 30132 14096 30144
rect 14148 30132 14154 30184
rect 14182 30132 14188 30184
rect 14240 30172 14246 30184
rect 15102 30172 15108 30184
rect 14240 30144 15108 30172
rect 14240 30132 14246 30144
rect 15102 30132 15108 30144
rect 15160 30132 15166 30184
rect 15470 30132 15476 30184
rect 15528 30172 15534 30184
rect 17402 30172 17408 30184
rect 15528 30144 17408 30172
rect 15528 30132 15534 30144
rect 17402 30132 17408 30144
rect 17460 30172 17466 30184
rect 20070 30172 20076 30184
rect 17460 30144 20076 30172
rect 17460 30132 17466 30144
rect 20070 30132 20076 30144
rect 20128 30172 20134 30184
rect 21174 30172 21180 30184
rect 20128 30144 21180 30172
rect 20128 30132 20134 30144
rect 21174 30132 21180 30144
rect 21232 30132 21238 30184
rect 23014 30132 23020 30184
rect 23072 30132 23078 30184
rect 23106 30132 23112 30184
rect 23164 30172 23170 30184
rect 23750 30172 23756 30184
rect 23164 30144 23756 30172
rect 23164 30132 23170 30144
rect 23750 30132 23756 30144
rect 23808 30132 23814 30184
rect 23844 30172 23872 30212
rect 24670 30200 24676 30212
rect 24728 30200 24734 30252
rect 24946 30200 24952 30252
rect 25004 30240 25010 30252
rect 25498 30240 25504 30252
rect 25004 30212 25504 30240
rect 25004 30200 25010 30212
rect 25498 30200 25504 30212
rect 25556 30200 25562 30252
rect 26237 30243 26295 30249
rect 26237 30240 26249 30243
rect 25608 30212 26249 30240
rect 25222 30172 25228 30184
rect 23844 30144 25228 30172
rect 25222 30132 25228 30144
rect 25280 30132 25286 30184
rect 25317 30175 25375 30181
rect 25317 30141 25329 30175
rect 25363 30172 25375 30175
rect 25406 30172 25412 30184
rect 25363 30144 25412 30172
rect 25363 30141 25375 30144
rect 25317 30135 25375 30141
rect 25406 30132 25412 30144
rect 25464 30132 25470 30184
rect 18138 30104 18144 30116
rect 11808 30076 18144 30104
rect 9490 30036 9496 30048
rect 9451 30008 9496 30036
rect 9490 29996 9496 30008
rect 9548 29996 9554 30048
rect 10410 29996 10416 30048
rect 10468 30036 10474 30048
rect 11808 30045 11836 30076
rect 18138 30064 18144 30076
rect 18196 30104 18202 30116
rect 18233 30107 18291 30113
rect 18233 30104 18245 30107
rect 18196 30076 18245 30104
rect 18196 30064 18202 30076
rect 18233 30073 18245 30076
rect 18279 30104 18291 30107
rect 18279 30076 19012 30104
rect 18279 30073 18291 30076
rect 18233 30067 18291 30073
rect 11793 30039 11851 30045
rect 11793 30036 11805 30039
rect 10468 30008 11805 30036
rect 10468 29996 10474 30008
rect 11793 30005 11805 30008
rect 11839 30005 11851 30039
rect 11793 29999 11851 30005
rect 12437 30039 12495 30045
rect 12437 30005 12449 30039
rect 12483 30036 12495 30039
rect 12802 30036 12808 30048
rect 12483 30008 12808 30036
rect 12483 30005 12495 30008
rect 12437 29999 12495 30005
rect 12802 29996 12808 30008
rect 12860 29996 12866 30048
rect 12986 30036 12992 30048
rect 12947 30008 12992 30036
rect 12986 29996 12992 30008
rect 13044 30036 13050 30048
rect 13262 30036 13268 30048
rect 13044 30008 13268 30036
rect 13044 29996 13050 30008
rect 13262 29996 13268 30008
rect 13320 29996 13326 30048
rect 14093 30039 14151 30045
rect 14093 30005 14105 30039
rect 14139 30036 14151 30039
rect 14366 30036 14372 30048
rect 14139 30008 14372 30036
rect 14139 30005 14151 30008
rect 14093 29999 14151 30005
rect 14366 29996 14372 30008
rect 14424 29996 14430 30048
rect 14458 29996 14464 30048
rect 14516 30036 14522 30048
rect 15749 30039 15807 30045
rect 15749 30036 15761 30039
rect 14516 30008 15761 30036
rect 14516 29996 14522 30008
rect 15749 30005 15761 30008
rect 15795 30036 15807 30039
rect 16022 30036 16028 30048
rect 15795 30008 16028 30036
rect 15795 30005 15807 30008
rect 15749 29999 15807 30005
rect 16022 29996 16028 30008
rect 16080 29996 16086 30048
rect 17221 30039 17279 30045
rect 17221 30005 17233 30039
rect 17267 30036 17279 30039
rect 17402 30036 17408 30048
rect 17267 30008 17408 30036
rect 17267 30005 17279 30008
rect 17221 29999 17279 30005
rect 17402 29996 17408 30008
rect 17460 29996 17466 30048
rect 17954 29996 17960 30048
rect 18012 30036 18018 30048
rect 18598 30036 18604 30048
rect 18012 30008 18604 30036
rect 18012 29996 18018 30008
rect 18598 29996 18604 30008
rect 18656 29996 18662 30048
rect 18874 30036 18880 30048
rect 18835 30008 18880 30036
rect 18874 29996 18880 30008
rect 18932 29996 18938 30048
rect 18984 30036 19012 30076
rect 19242 30064 19248 30116
rect 19300 30104 19306 30116
rect 21542 30104 21548 30116
rect 19300 30076 21548 30104
rect 19300 30064 19306 30076
rect 21542 30064 21548 30076
rect 21600 30064 21606 30116
rect 21910 30064 21916 30116
rect 21968 30104 21974 30116
rect 22922 30104 22928 30116
rect 21968 30076 22928 30104
rect 21968 30064 21974 30076
rect 22922 30064 22928 30076
rect 22980 30064 22986 30116
rect 23566 30064 23572 30116
rect 23624 30104 23630 30116
rect 23624 30076 23888 30104
rect 23624 30064 23630 30076
rect 22186 30036 22192 30048
rect 18984 30008 22192 30036
rect 22186 29996 22192 30008
rect 22244 29996 22250 30048
rect 22465 30039 22523 30045
rect 22465 30005 22477 30039
rect 22511 30036 22523 30039
rect 22646 30036 22652 30048
rect 22511 30008 22652 30036
rect 22511 30005 22523 30008
rect 22465 29999 22523 30005
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 23106 30036 23112 30048
rect 23067 30008 23112 30036
rect 23106 29996 23112 30008
rect 23164 29996 23170 30048
rect 23198 29996 23204 30048
rect 23256 30036 23262 30048
rect 23860 30045 23888 30076
rect 24118 30064 24124 30116
rect 24176 30104 24182 30116
rect 24762 30104 24768 30116
rect 24176 30076 24768 30104
rect 24176 30064 24182 30076
rect 24762 30064 24768 30076
rect 24820 30064 24826 30116
rect 24857 30107 24915 30113
rect 24857 30073 24869 30107
rect 24903 30104 24915 30107
rect 25608 30104 25636 30212
rect 26237 30209 26249 30212
rect 26283 30209 26295 30243
rect 26325 30240 26353 30280
rect 26421 30277 26433 30311
rect 26467 30308 26479 30311
rect 26786 30308 26792 30320
rect 26467 30280 26792 30308
rect 26467 30277 26479 30280
rect 26421 30271 26479 30277
rect 26786 30268 26792 30280
rect 26844 30268 26850 30320
rect 26977 30240 27005 30348
rect 27982 30336 27988 30348
rect 28040 30336 28046 30388
rect 30006 30308 30012 30320
rect 27264 30280 30012 30308
rect 26325 30212 27005 30240
rect 26237 30203 26295 30209
rect 27062 30200 27068 30252
rect 27120 30240 27126 30252
rect 27157 30243 27215 30249
rect 27157 30240 27169 30243
rect 27120 30212 27169 30240
rect 27120 30200 27126 30212
rect 27157 30209 27169 30212
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 25685 30175 25743 30181
rect 25685 30141 25697 30175
rect 25731 30141 25743 30175
rect 25685 30135 25743 30141
rect 24903 30076 25636 30104
rect 25700 30104 25728 30135
rect 26050 30132 26056 30184
rect 26108 30172 26114 30184
rect 27264 30172 27292 30280
rect 27816 30249 27844 30280
rect 30006 30268 30012 30280
rect 30064 30268 30070 30320
rect 30098 30268 30104 30320
rect 30156 30308 30162 30320
rect 30156 30280 31064 30308
rect 30156 30268 30162 30280
rect 27341 30243 27399 30249
rect 27341 30209 27353 30243
rect 27387 30209 27399 30243
rect 27341 30203 27399 30209
rect 27801 30243 27859 30249
rect 27801 30209 27813 30243
rect 27847 30209 27859 30243
rect 27801 30203 27859 30209
rect 26108 30144 27292 30172
rect 26108 30132 26114 30144
rect 26234 30104 26240 30116
rect 25700 30076 26240 30104
rect 24903 30073 24915 30076
rect 24857 30067 24915 30073
rect 26234 30064 26240 30076
rect 26292 30064 26298 30116
rect 26786 30064 26792 30116
rect 26844 30104 26850 30116
rect 27356 30104 27384 30203
rect 27982 30200 27988 30252
rect 28040 30240 28046 30252
rect 28445 30243 28503 30249
rect 28040 30212 28133 30240
rect 28040 30200 28046 30212
rect 28445 30209 28457 30243
rect 28491 30240 28503 30243
rect 28534 30240 28540 30252
rect 28491 30212 28540 30240
rect 28491 30209 28503 30212
rect 28445 30203 28503 30209
rect 28534 30200 28540 30212
rect 28592 30200 28598 30252
rect 28902 30200 28908 30252
rect 28960 30240 28966 30252
rect 29089 30243 29147 30249
rect 29089 30240 29101 30243
rect 28960 30212 29101 30240
rect 28960 30200 28966 30212
rect 29089 30209 29101 30212
rect 29135 30209 29147 30243
rect 29730 30240 29736 30252
rect 29691 30212 29736 30240
rect 29089 30203 29147 30209
rect 29730 30200 29736 30212
rect 29788 30200 29794 30252
rect 30190 30200 30196 30252
rect 30248 30240 30254 30252
rect 31036 30249 31064 30280
rect 30377 30243 30435 30249
rect 30377 30240 30389 30243
rect 30248 30212 30389 30240
rect 30248 30200 30254 30212
rect 30377 30209 30389 30212
rect 30423 30209 30435 30243
rect 30377 30203 30435 30209
rect 31021 30243 31079 30249
rect 31021 30209 31033 30243
rect 31067 30209 31079 30243
rect 31021 30203 31079 30209
rect 27430 30132 27436 30184
rect 27488 30172 27494 30184
rect 27890 30172 27896 30184
rect 27488 30144 27896 30172
rect 27488 30132 27494 30144
rect 27890 30132 27896 30144
rect 27948 30132 27954 30184
rect 28000 30172 28028 30200
rect 29546 30172 29552 30184
rect 28000 30144 29552 30172
rect 29546 30132 29552 30144
rect 29604 30132 29610 30184
rect 29273 30107 29331 30113
rect 26844 30076 28764 30104
rect 26844 30064 26850 30076
rect 23661 30039 23719 30045
rect 23661 30036 23673 30039
rect 23256 30008 23673 30036
rect 23256 29996 23262 30008
rect 23661 30005 23673 30008
rect 23707 30005 23719 30039
rect 23661 29999 23719 30005
rect 23845 30039 23903 30045
rect 23845 30005 23857 30039
rect 23891 30005 23903 30039
rect 24670 30036 24676 30048
rect 24631 30008 24676 30036
rect 23845 29999 23903 30005
rect 24670 29996 24676 30008
rect 24728 30036 24734 30048
rect 27062 30036 27068 30048
rect 24728 30008 27068 30036
rect 24728 29996 24734 30008
rect 27062 29996 27068 30008
rect 27120 29996 27126 30048
rect 27249 30039 27307 30045
rect 27249 30005 27261 30039
rect 27295 30036 27307 30039
rect 27338 30036 27344 30048
rect 27295 30008 27344 30036
rect 27295 30005 27307 30008
rect 27249 29999 27307 30005
rect 27338 29996 27344 30008
rect 27396 29996 27402 30048
rect 27801 30039 27859 30045
rect 27801 30005 27813 30039
rect 27847 30036 27859 30039
rect 28074 30036 28080 30048
rect 27847 30008 28080 30036
rect 27847 30005 27859 30008
rect 27801 29999 27859 30005
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 28626 30036 28632 30048
rect 28587 30008 28632 30036
rect 28626 29996 28632 30008
rect 28684 29996 28690 30048
rect 28736 30036 28764 30076
rect 29273 30073 29285 30107
rect 29319 30104 29331 30107
rect 29822 30104 29828 30116
rect 29319 30076 29828 30104
rect 29319 30073 29331 30076
rect 29273 30067 29331 30073
rect 29822 30064 29828 30076
rect 29880 30064 29886 30116
rect 29454 30036 29460 30048
rect 28736 30008 29460 30036
rect 29454 29996 29460 30008
rect 29512 29996 29518 30048
rect 29917 30039 29975 30045
rect 29917 30005 29929 30039
rect 29963 30036 29975 30039
rect 30374 30036 30380 30048
rect 29963 30008 30380 30036
rect 29963 30005 29975 30008
rect 29917 29999 29975 30005
rect 30374 29996 30380 30008
rect 30432 29996 30438 30048
rect 30558 30036 30564 30048
rect 30519 30008 30564 30036
rect 30558 29996 30564 30008
rect 30616 29996 30622 30048
rect 31202 30036 31208 30048
rect 31163 30008 31208 30036
rect 31202 29996 31208 30008
rect 31260 29996 31266 30048
rect 1104 29946 31832 29968
rect 1104 29894 4791 29946
rect 4843 29894 4855 29946
rect 4907 29894 4919 29946
rect 4971 29894 4983 29946
rect 5035 29894 5047 29946
rect 5099 29894 12473 29946
rect 12525 29894 12537 29946
rect 12589 29894 12601 29946
rect 12653 29894 12665 29946
rect 12717 29894 12729 29946
rect 12781 29894 20155 29946
rect 20207 29894 20219 29946
rect 20271 29894 20283 29946
rect 20335 29894 20347 29946
rect 20399 29894 20411 29946
rect 20463 29894 27837 29946
rect 27889 29894 27901 29946
rect 27953 29894 27965 29946
rect 28017 29894 28029 29946
rect 28081 29894 28093 29946
rect 28145 29894 31832 29946
rect 1104 29872 31832 29894
rect 8573 29835 8631 29841
rect 8573 29801 8585 29835
rect 8619 29832 8631 29835
rect 11238 29832 11244 29844
rect 8619 29804 11244 29832
rect 8619 29801 8631 29804
rect 8573 29795 8631 29801
rect 11238 29792 11244 29804
rect 11296 29792 11302 29844
rect 13173 29835 13231 29841
rect 13173 29801 13185 29835
rect 13219 29832 13231 29835
rect 13354 29832 13360 29844
rect 13219 29804 13360 29832
rect 13219 29801 13231 29804
rect 13173 29795 13231 29801
rect 13354 29792 13360 29804
rect 13412 29792 13418 29844
rect 14366 29792 14372 29844
rect 14424 29832 14430 29844
rect 14829 29835 14887 29841
rect 14829 29832 14841 29835
rect 14424 29804 14841 29832
rect 14424 29792 14430 29804
rect 14829 29801 14841 29804
rect 14875 29832 14887 29835
rect 16850 29832 16856 29844
rect 14875 29804 16856 29832
rect 14875 29801 14887 29804
rect 14829 29795 14887 29801
rect 16850 29792 16856 29804
rect 16908 29792 16914 29844
rect 16942 29792 16948 29844
rect 17000 29832 17006 29844
rect 17770 29832 17776 29844
rect 17000 29804 17776 29832
rect 17000 29792 17006 29804
rect 17770 29792 17776 29804
rect 17828 29792 17834 29844
rect 18141 29835 18199 29841
rect 18141 29801 18153 29835
rect 18187 29832 18199 29835
rect 18230 29832 18236 29844
rect 18187 29804 18236 29832
rect 18187 29801 18199 29804
rect 18141 29795 18199 29801
rect 18230 29792 18236 29804
rect 18288 29832 18294 29844
rect 19426 29832 19432 29844
rect 18288 29804 19432 29832
rect 18288 29792 18294 29804
rect 19426 29792 19432 29804
rect 19484 29792 19490 29844
rect 19978 29792 19984 29844
rect 20036 29832 20042 29844
rect 20165 29835 20223 29841
rect 20165 29832 20177 29835
rect 20036 29804 20177 29832
rect 20036 29792 20042 29804
rect 20165 29801 20177 29804
rect 20211 29801 20223 29835
rect 20165 29795 20223 29801
rect 20346 29792 20352 29844
rect 20404 29832 20410 29844
rect 20714 29832 20720 29844
rect 20404 29804 20720 29832
rect 20404 29792 20410 29804
rect 20714 29792 20720 29804
rect 20772 29792 20778 29844
rect 20901 29835 20959 29841
rect 20901 29801 20913 29835
rect 20947 29832 20959 29835
rect 21358 29832 21364 29844
rect 20947 29804 21364 29832
rect 20947 29801 20959 29804
rect 20901 29795 20959 29801
rect 21358 29792 21364 29804
rect 21416 29792 21422 29844
rect 22094 29792 22100 29844
rect 22152 29832 22158 29844
rect 23661 29835 23719 29841
rect 23661 29832 23673 29835
rect 22152 29804 23673 29832
rect 22152 29792 22158 29804
rect 23661 29801 23673 29804
rect 23707 29832 23719 29835
rect 24118 29832 24124 29844
rect 23707 29804 24124 29832
rect 23707 29801 23719 29804
rect 23661 29795 23719 29801
rect 24118 29792 24124 29804
rect 24176 29792 24182 29844
rect 24210 29792 24216 29844
rect 24268 29832 24274 29844
rect 24854 29832 24860 29844
rect 24268 29804 24860 29832
rect 24268 29792 24274 29804
rect 24854 29792 24860 29804
rect 24912 29792 24918 29844
rect 25222 29792 25228 29844
rect 25280 29832 25286 29844
rect 25685 29835 25743 29841
rect 25685 29832 25697 29835
rect 25280 29804 25697 29832
rect 25280 29792 25286 29804
rect 25685 29801 25697 29804
rect 25731 29801 25743 29835
rect 25866 29832 25872 29844
rect 25827 29804 25872 29832
rect 25685 29795 25743 29801
rect 25866 29792 25872 29804
rect 25924 29832 25930 29844
rect 26142 29832 26148 29844
rect 25924 29804 26148 29832
rect 25924 29792 25930 29804
rect 26142 29792 26148 29804
rect 26200 29792 26206 29844
rect 26326 29792 26332 29844
rect 26384 29792 26390 29844
rect 26602 29832 26608 29844
rect 26563 29804 26608 29832
rect 26602 29792 26608 29804
rect 26660 29792 26666 29844
rect 26970 29792 26976 29844
rect 27028 29832 27034 29844
rect 29178 29832 29184 29844
rect 27028 29804 29184 29832
rect 27028 29792 27034 29804
rect 29178 29792 29184 29804
rect 29236 29792 29242 29844
rect 9861 29767 9919 29773
rect 9861 29733 9873 29767
rect 9907 29764 9919 29767
rect 9950 29764 9956 29776
rect 9907 29736 9956 29764
rect 9907 29733 9919 29736
rect 9861 29727 9919 29733
rect 9950 29724 9956 29736
rect 10008 29724 10014 29776
rect 10502 29724 10508 29776
rect 10560 29764 10566 29776
rect 14182 29764 14188 29776
rect 10560 29736 14188 29764
rect 10560 29724 10566 29736
rect 14182 29724 14188 29736
rect 14240 29724 14246 29776
rect 16206 29764 16212 29776
rect 14292 29736 16212 29764
rect 10965 29699 11023 29705
rect 10965 29665 10977 29699
rect 11011 29696 11023 29699
rect 11146 29696 11152 29708
rect 11011 29668 11152 29696
rect 11011 29665 11023 29668
rect 10965 29659 11023 29665
rect 9398 29588 9404 29640
rect 9456 29628 9462 29640
rect 10321 29631 10379 29637
rect 10321 29628 10333 29631
rect 9456 29600 10333 29628
rect 9456 29588 9462 29600
rect 10321 29597 10333 29600
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 9582 29520 9588 29572
rect 9640 29560 9646 29572
rect 10980 29560 11008 29659
rect 11146 29656 11152 29668
rect 11204 29656 11210 29708
rect 11238 29656 11244 29708
rect 11296 29696 11302 29708
rect 13078 29696 13084 29708
rect 11296 29668 13084 29696
rect 11296 29656 11302 29668
rect 13078 29656 13084 29668
rect 13136 29696 13142 29708
rect 14292 29696 14320 29736
rect 16206 29724 16212 29736
rect 16264 29764 16270 29776
rect 18693 29767 18751 29773
rect 18693 29764 18705 29767
rect 16264 29736 18705 29764
rect 16264 29724 16270 29736
rect 18693 29733 18705 29736
rect 18739 29764 18751 29767
rect 18782 29764 18788 29776
rect 18739 29736 18788 29764
rect 18739 29733 18751 29736
rect 18693 29727 18751 29733
rect 18782 29724 18788 29736
rect 18840 29724 18846 29776
rect 20254 29724 20260 29776
rect 20312 29764 20318 29776
rect 20312 29736 20760 29764
rect 20312 29724 20318 29736
rect 13136 29668 14320 29696
rect 13136 29656 13142 29668
rect 14642 29656 14648 29708
rect 14700 29696 14706 29708
rect 15933 29699 15991 29705
rect 15933 29696 15945 29699
rect 14700 29668 15945 29696
rect 14700 29656 14706 29668
rect 15933 29665 15945 29668
rect 15979 29696 15991 29699
rect 19242 29696 19248 29708
rect 15979 29668 19248 29696
rect 15979 29665 15991 29668
rect 15933 29659 15991 29665
rect 19242 29656 19248 29668
rect 19300 29696 19306 29708
rect 19610 29696 19616 29708
rect 19300 29668 19616 29696
rect 19300 29656 19306 29668
rect 19610 29656 19616 29668
rect 19668 29656 19674 29708
rect 19886 29656 19892 29708
rect 19944 29696 19950 29708
rect 20622 29696 20628 29708
rect 19944 29668 20628 29696
rect 19944 29656 19950 29668
rect 20622 29656 20628 29668
rect 20680 29656 20686 29708
rect 20732 29696 20760 29736
rect 21174 29724 21180 29776
rect 21232 29764 21238 29776
rect 21232 29736 21864 29764
rect 21232 29724 21238 29736
rect 20732 29668 21036 29696
rect 17126 29588 17132 29640
rect 17184 29628 17190 29640
rect 19518 29628 19524 29640
rect 17184 29600 19524 29628
rect 17184 29588 17190 29600
rect 19518 29588 19524 29600
rect 19576 29628 19582 29640
rect 19978 29628 19984 29640
rect 19576 29600 19984 29628
rect 19576 29588 19582 29600
rect 19978 29588 19984 29600
rect 20036 29628 20042 29640
rect 20714 29628 20720 29640
rect 20036 29600 20720 29628
rect 20036 29588 20042 29600
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 21008 29638 21036 29668
rect 21266 29656 21272 29708
rect 21324 29696 21330 29708
rect 21836 29696 21864 29736
rect 21910 29724 21916 29776
rect 21968 29764 21974 29776
rect 22189 29767 22247 29773
rect 22189 29764 22201 29767
rect 21968 29736 22201 29764
rect 21968 29724 21974 29736
rect 22189 29733 22201 29736
rect 22235 29733 22247 29767
rect 22189 29727 22247 29733
rect 22830 29724 22836 29776
rect 22888 29764 22894 29776
rect 23201 29767 23259 29773
rect 23201 29764 23213 29767
rect 22888 29736 23213 29764
rect 22888 29724 22894 29736
rect 23201 29733 23213 29736
rect 23247 29764 23259 29767
rect 23934 29764 23940 29776
rect 23247 29736 23940 29764
rect 23247 29733 23259 29736
rect 23201 29727 23259 29733
rect 23934 29724 23940 29736
rect 23992 29724 23998 29776
rect 24029 29767 24087 29773
rect 24029 29733 24041 29767
rect 24075 29764 24087 29767
rect 26050 29764 26056 29776
rect 24075 29736 26056 29764
rect 24075 29733 24087 29736
rect 24029 29727 24087 29733
rect 26050 29724 26056 29736
rect 26108 29724 26114 29776
rect 26344 29764 26372 29792
rect 28077 29767 28135 29773
rect 28077 29764 28089 29767
rect 26344 29736 28089 29764
rect 28077 29733 28089 29736
rect 28123 29733 28135 29767
rect 28077 29727 28135 29733
rect 28350 29724 28356 29776
rect 28408 29764 28414 29776
rect 30098 29764 30104 29776
rect 28408 29736 30104 29764
rect 28408 29724 28414 29736
rect 30098 29724 30104 29736
rect 30156 29724 30162 29776
rect 21324 29668 21680 29696
rect 21836 29668 22232 29696
rect 21324 29656 21330 29668
rect 21174 29638 21180 29640
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29597 20867 29631
rect 21008 29610 21180 29638
rect 20809 29591 20867 29597
rect 9640 29532 11008 29560
rect 11517 29563 11575 29569
rect 9640 29520 9646 29532
rect 11517 29529 11529 29563
rect 11563 29560 11575 29563
rect 12342 29560 12348 29572
rect 11563 29532 12348 29560
rect 11563 29529 11575 29532
rect 11517 29523 11575 29529
rect 12342 29520 12348 29532
rect 12400 29560 12406 29572
rect 12621 29563 12679 29569
rect 12621 29560 12633 29563
rect 12400 29532 12633 29560
rect 12400 29520 12406 29532
rect 12621 29529 12633 29532
rect 12667 29560 12679 29563
rect 14826 29560 14832 29572
rect 12667 29532 14832 29560
rect 12667 29529 12679 29532
rect 12621 29523 12679 29529
rect 14826 29520 14832 29532
rect 14884 29520 14890 29572
rect 17034 29560 17040 29572
rect 15166 29532 17040 29560
rect 7834 29452 7840 29504
rect 7892 29492 7898 29504
rect 9217 29495 9275 29501
rect 9217 29492 9229 29495
rect 7892 29464 9229 29492
rect 7892 29452 7898 29464
rect 9217 29461 9229 29464
rect 9263 29492 9275 29495
rect 10502 29492 10508 29504
rect 9263 29464 10508 29492
rect 9263 29461 9275 29464
rect 9217 29455 9275 29461
rect 10502 29452 10508 29464
rect 10560 29452 10566 29504
rect 12066 29492 12072 29504
rect 12027 29464 12072 29492
rect 12066 29452 12072 29464
rect 12124 29452 12130 29504
rect 13725 29495 13783 29501
rect 13725 29461 13737 29495
rect 13771 29492 13783 29495
rect 14182 29492 14188 29504
rect 13771 29464 14188 29492
rect 13771 29461 13783 29464
rect 13725 29455 13783 29461
rect 14182 29452 14188 29464
rect 14240 29452 14246 29504
rect 15010 29452 15016 29504
rect 15068 29492 15074 29504
rect 15166 29492 15194 29532
rect 17034 29520 17040 29532
rect 17092 29520 17098 29572
rect 17678 29520 17684 29572
rect 17736 29560 17742 29572
rect 17736 29532 18457 29560
rect 17736 29520 17742 29532
rect 15068 29464 15194 29492
rect 15381 29495 15439 29501
rect 15068 29452 15074 29464
rect 15381 29461 15393 29495
rect 15427 29492 15439 29495
rect 16022 29492 16028 29504
rect 15427 29464 16028 29492
rect 15427 29461 15439 29464
rect 15381 29455 15439 29461
rect 16022 29452 16028 29464
rect 16080 29452 16086 29504
rect 16485 29495 16543 29501
rect 16485 29461 16497 29495
rect 16531 29492 16543 29495
rect 16850 29492 16856 29504
rect 16531 29464 16856 29492
rect 16531 29461 16543 29464
rect 16485 29455 16543 29461
rect 16850 29452 16856 29464
rect 16908 29452 16914 29504
rect 16945 29495 17003 29501
rect 16945 29461 16957 29495
rect 16991 29492 17003 29495
rect 17218 29492 17224 29504
rect 16991 29464 17224 29492
rect 16991 29461 17003 29464
rect 16945 29455 17003 29461
rect 17218 29452 17224 29464
rect 17276 29452 17282 29504
rect 17586 29492 17592 29504
rect 17499 29464 17592 29492
rect 17586 29452 17592 29464
rect 17644 29492 17650 29504
rect 18322 29492 18328 29504
rect 17644 29464 18328 29492
rect 17644 29452 17650 29464
rect 18322 29452 18328 29464
rect 18380 29452 18386 29504
rect 18429 29492 18457 29532
rect 19058 29520 19064 29572
rect 19116 29560 19122 29572
rect 19429 29563 19487 29569
rect 19429 29560 19441 29563
rect 19116 29532 19441 29560
rect 19116 29520 19122 29532
rect 19429 29529 19441 29532
rect 19475 29529 19487 29563
rect 19429 29523 19487 29529
rect 20162 29520 20168 29572
rect 20220 29560 20226 29572
rect 20346 29560 20352 29572
rect 20220 29532 20352 29560
rect 20220 29520 20226 29532
rect 20346 29520 20352 29532
rect 20404 29520 20410 29572
rect 20438 29520 20444 29572
rect 20496 29560 20502 29572
rect 20824 29560 20852 29591
rect 21174 29588 21180 29610
rect 21232 29588 21238 29640
rect 21450 29628 21456 29640
rect 21411 29600 21456 29628
rect 21450 29588 21456 29600
rect 21508 29588 21514 29640
rect 21652 29637 21680 29668
rect 21637 29631 21695 29637
rect 21637 29597 21649 29631
rect 21683 29628 21695 29631
rect 21910 29628 21916 29640
rect 21683 29600 21916 29628
rect 21683 29597 21695 29600
rect 21637 29591 21695 29597
rect 21910 29588 21916 29600
rect 21968 29628 21974 29640
rect 22097 29631 22155 29637
rect 22097 29628 22109 29631
rect 21968 29600 22109 29628
rect 21968 29588 21974 29600
rect 22097 29597 22109 29600
rect 22143 29597 22155 29631
rect 22204 29628 22232 29668
rect 22278 29656 22284 29708
rect 22336 29696 22342 29708
rect 23566 29696 23572 29708
rect 22336 29668 23060 29696
rect 22336 29656 22342 29668
rect 22373 29631 22431 29637
rect 22373 29628 22385 29631
rect 22204 29600 22385 29628
rect 22097 29591 22155 29597
rect 22373 29597 22385 29600
rect 22419 29628 22431 29631
rect 22554 29628 22560 29640
rect 22419 29600 22560 29628
rect 22419 29597 22431 29600
rect 22373 29591 22431 29597
rect 22554 29588 22560 29600
rect 22612 29588 22618 29640
rect 23032 29637 23060 29668
rect 23308 29668 23572 29696
rect 23308 29640 23336 29668
rect 23566 29656 23572 29668
rect 23624 29656 23630 29708
rect 23750 29656 23756 29708
rect 23808 29696 23814 29708
rect 24949 29699 25007 29705
rect 24949 29696 24961 29699
rect 23808 29668 24961 29696
rect 23808 29656 23814 29668
rect 24949 29665 24961 29668
rect 24995 29665 25007 29699
rect 24949 29659 25007 29665
rect 25133 29699 25191 29705
rect 25133 29665 25145 29699
rect 25179 29696 25191 29699
rect 26326 29696 26332 29708
rect 25179 29668 26332 29696
rect 25179 29665 25191 29668
rect 25133 29659 25191 29665
rect 26326 29656 26332 29668
rect 26384 29656 26390 29708
rect 27341 29699 27399 29705
rect 27341 29665 27353 29699
rect 27387 29696 27399 29699
rect 27430 29696 27436 29708
rect 27387 29668 27436 29696
rect 27387 29665 27399 29668
rect 27341 29659 27399 29665
rect 27430 29656 27436 29668
rect 27488 29656 27494 29708
rect 27522 29656 27528 29708
rect 27580 29696 27586 29708
rect 27706 29696 27712 29708
rect 27580 29668 27712 29696
rect 27580 29656 27586 29668
rect 27706 29656 27712 29668
rect 27764 29656 27770 29708
rect 28185 29668 28396 29696
rect 22925 29631 22983 29637
rect 22925 29597 22937 29631
rect 22971 29597 22983 29631
rect 22925 29591 22983 29597
rect 23017 29631 23075 29637
rect 23017 29597 23029 29631
rect 23063 29628 23075 29631
rect 23290 29628 23296 29640
rect 23063 29600 23296 29628
rect 23063 29597 23075 29600
rect 23017 29591 23075 29597
rect 20990 29560 20996 29572
rect 20496 29532 20996 29560
rect 20496 29520 20502 29532
rect 20990 29520 20996 29532
rect 21048 29520 21054 29572
rect 21468 29560 21496 29588
rect 22186 29560 22192 29572
rect 21468 29532 22192 29560
rect 22186 29520 22192 29532
rect 22244 29520 22250 29572
rect 22281 29563 22339 29569
rect 22281 29529 22293 29563
rect 22327 29560 22339 29563
rect 22940 29560 22968 29591
rect 23290 29588 23296 29600
rect 23348 29588 23354 29640
rect 23658 29628 23664 29640
rect 23619 29600 23664 29628
rect 23658 29588 23664 29600
rect 23716 29588 23722 29640
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29628 23903 29631
rect 24670 29628 24676 29640
rect 23891 29600 24676 29628
rect 23891 29597 23903 29600
rect 23845 29591 23903 29597
rect 24670 29588 24676 29600
rect 24728 29588 24734 29640
rect 24854 29628 24860 29640
rect 24815 29600 24860 29628
rect 24854 29588 24860 29600
rect 24912 29588 24918 29640
rect 25225 29631 25283 29637
rect 25225 29597 25237 29631
rect 25271 29628 25283 29631
rect 25590 29628 25596 29640
rect 25271 29600 25596 29628
rect 25271 29597 25283 29600
rect 25225 29591 25283 29597
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 26510 29628 26516 29640
rect 25700 29600 26372 29628
rect 26471 29600 26516 29628
rect 22327 29532 22876 29560
rect 22940 29532 23060 29560
rect 22327 29529 22339 29532
rect 22281 29523 22339 29529
rect 22848 29504 22876 29532
rect 21453 29495 21511 29501
rect 21453 29492 21465 29495
rect 18429 29464 21465 29492
rect 21453 29461 21465 29464
rect 21499 29461 21511 29495
rect 21453 29455 21511 29461
rect 22830 29452 22836 29504
rect 22888 29452 22894 29504
rect 23032 29492 23060 29532
rect 23566 29520 23572 29572
rect 23624 29560 23630 29572
rect 25700 29560 25728 29600
rect 26053 29563 26111 29569
rect 23624 29532 25728 29560
rect 25792 29532 26004 29560
rect 23624 29520 23630 29532
rect 24210 29492 24216 29504
rect 23032 29464 24216 29492
rect 24210 29452 24216 29464
rect 24268 29452 24274 29504
rect 24857 29495 24915 29501
rect 24857 29461 24869 29495
rect 24903 29492 24915 29495
rect 25792 29492 25820 29532
rect 25866 29501 25872 29504
rect 24903 29464 25820 29492
rect 25853 29495 25872 29501
rect 24903 29461 24915 29464
rect 24857 29455 24915 29461
rect 25853 29461 25865 29495
rect 25853 29455 25872 29461
rect 25866 29452 25872 29455
rect 25924 29452 25930 29504
rect 25976 29492 26004 29532
rect 26053 29529 26065 29563
rect 26099 29560 26111 29563
rect 26234 29560 26240 29572
rect 26099 29532 26240 29560
rect 26099 29529 26111 29532
rect 26053 29523 26111 29529
rect 26234 29520 26240 29532
rect 26292 29520 26298 29572
rect 26344 29560 26372 29600
rect 26510 29588 26516 29600
rect 26568 29588 26574 29640
rect 26605 29631 26663 29637
rect 26605 29597 26617 29631
rect 26651 29628 26663 29631
rect 27890 29628 27896 29640
rect 26651 29600 27896 29628
rect 26651 29597 26663 29600
rect 26605 29591 26663 29597
rect 26620 29560 26648 29591
rect 27890 29588 27896 29600
rect 27948 29588 27954 29640
rect 28074 29628 28080 29640
rect 28035 29600 28080 29628
rect 28074 29588 28080 29600
rect 28132 29588 28138 29640
rect 27525 29563 27583 29569
rect 26344 29532 26648 29560
rect 26804 29532 27475 29560
rect 26804 29492 26832 29532
rect 25976 29464 26832 29492
rect 26881 29495 26939 29501
rect 26881 29461 26893 29495
rect 26927 29492 26939 29495
rect 27338 29492 27344 29504
rect 26927 29464 27344 29492
rect 26927 29461 26939 29464
rect 26881 29455 26939 29461
rect 27338 29452 27344 29464
rect 27396 29452 27402 29504
rect 27447 29492 27475 29532
rect 27525 29529 27537 29563
rect 27571 29560 27583 29563
rect 28185 29560 28213 29668
rect 28261 29631 28319 29637
rect 28261 29597 28273 29631
rect 28307 29597 28319 29631
rect 28368 29628 28396 29668
rect 28626 29656 28632 29708
rect 28684 29696 28690 29708
rect 28684 29668 30420 29696
rect 28684 29656 28690 29668
rect 28810 29628 28816 29640
rect 28368 29600 28672 29628
rect 28771 29600 28816 29628
rect 28261 29591 28319 29597
rect 27571 29532 28213 29560
rect 28276 29560 28304 29591
rect 28644 29572 28672 29600
rect 28810 29588 28816 29600
rect 28868 29588 28874 29640
rect 28905 29631 28963 29637
rect 28905 29597 28917 29631
rect 28951 29628 28963 29631
rect 28994 29628 29000 29640
rect 28951 29600 29000 29628
rect 28951 29597 28963 29600
rect 28905 29591 28963 29597
rect 28350 29560 28356 29572
rect 28276 29532 28356 29560
rect 27571 29529 27583 29532
rect 27525 29523 27583 29529
rect 28350 29520 28356 29532
rect 28408 29520 28414 29572
rect 28626 29520 28632 29572
rect 28684 29520 28690 29572
rect 28920 29560 28948 29591
rect 28994 29588 29000 29600
rect 29052 29588 29058 29640
rect 29914 29628 29920 29640
rect 29875 29600 29920 29628
rect 29914 29588 29920 29600
rect 29972 29588 29978 29640
rect 30392 29637 30420 29668
rect 30377 29631 30435 29637
rect 30377 29597 30389 29631
rect 30423 29597 30435 29631
rect 30377 29591 30435 29597
rect 31110 29588 31116 29640
rect 31168 29628 31174 29640
rect 31297 29631 31355 29637
rect 31297 29628 31309 29631
rect 31168 29600 31309 29628
rect 31168 29588 31174 29600
rect 31297 29597 31309 29600
rect 31343 29597 31355 29631
rect 31297 29591 31355 29597
rect 28920 29532 31340 29560
rect 31312 29504 31340 29532
rect 28994 29492 29000 29504
rect 27447 29464 29000 29492
rect 28994 29452 29000 29464
rect 29052 29452 29058 29504
rect 30561 29495 30619 29501
rect 30561 29461 30573 29495
rect 30607 29492 30619 29495
rect 31018 29492 31024 29504
rect 30607 29464 31024 29492
rect 30607 29461 30619 29464
rect 30561 29455 30619 29461
rect 31018 29452 31024 29464
rect 31076 29452 31082 29504
rect 31294 29452 31300 29504
rect 31352 29452 31358 29504
rect 1104 29402 31992 29424
rect 1104 29350 8632 29402
rect 8684 29350 8696 29402
rect 8748 29350 8760 29402
rect 8812 29350 8824 29402
rect 8876 29350 8888 29402
rect 8940 29350 16314 29402
rect 16366 29350 16378 29402
rect 16430 29350 16442 29402
rect 16494 29350 16506 29402
rect 16558 29350 16570 29402
rect 16622 29350 23996 29402
rect 24048 29350 24060 29402
rect 24112 29350 24124 29402
rect 24176 29350 24188 29402
rect 24240 29350 24252 29402
rect 24304 29350 31678 29402
rect 31730 29350 31742 29402
rect 31794 29350 31806 29402
rect 31858 29350 31870 29402
rect 31922 29350 31934 29402
rect 31986 29350 31992 29402
rect 1104 29328 31992 29350
rect 8389 29291 8447 29297
rect 8389 29257 8401 29291
rect 8435 29288 8447 29291
rect 10410 29288 10416 29300
rect 8435 29260 10416 29288
rect 8435 29257 8447 29260
rect 8389 29251 8447 29257
rect 10410 29248 10416 29260
rect 10468 29248 10474 29300
rect 12250 29288 12256 29300
rect 11992 29260 12256 29288
rect 7837 29223 7895 29229
rect 7837 29189 7849 29223
rect 7883 29220 7895 29223
rect 9030 29220 9036 29232
rect 7883 29192 9036 29220
rect 7883 29189 7895 29192
rect 7837 29183 7895 29189
rect 9030 29180 9036 29192
rect 9088 29180 9094 29232
rect 9493 29223 9551 29229
rect 9493 29189 9505 29223
rect 9539 29220 9551 29223
rect 11992 29220 12020 29260
rect 12250 29248 12256 29260
rect 12308 29248 12314 29300
rect 12437 29291 12495 29297
rect 12437 29257 12449 29291
rect 12483 29288 12495 29291
rect 12802 29288 12808 29300
rect 12483 29260 12808 29288
rect 12483 29257 12495 29260
rect 12437 29251 12495 29257
rect 12802 29248 12808 29260
rect 12860 29288 12866 29300
rect 13630 29288 13636 29300
rect 12860 29260 13636 29288
rect 12860 29248 12866 29260
rect 13630 29248 13636 29260
rect 13688 29248 13694 29300
rect 15197 29291 15255 29297
rect 15197 29257 15209 29291
rect 15243 29288 15255 29291
rect 15470 29288 15476 29300
rect 15243 29260 15476 29288
rect 15243 29257 15255 29260
rect 15197 29251 15255 29257
rect 9539 29192 12020 29220
rect 9539 29189 9551 29192
rect 9493 29183 9551 29189
rect 12066 29180 12072 29232
rect 12124 29220 12130 29232
rect 13722 29220 13728 29232
rect 12124 29192 13728 29220
rect 12124 29180 12130 29192
rect 11146 29112 11152 29164
rect 11204 29152 11210 29164
rect 11793 29155 11851 29161
rect 11793 29152 11805 29155
rect 11204 29124 11805 29152
rect 11204 29112 11210 29124
rect 11793 29121 11805 29124
rect 11839 29152 11851 29155
rect 11882 29152 11888 29164
rect 11839 29124 11888 29152
rect 11839 29121 11851 29124
rect 11793 29115 11851 29121
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 8941 29087 8999 29093
rect 8941 29053 8953 29087
rect 8987 29084 8999 29087
rect 10505 29087 10563 29093
rect 10505 29084 10517 29087
rect 8987 29056 10517 29084
rect 8987 29053 8999 29056
rect 8941 29047 8999 29053
rect 10505 29053 10517 29056
rect 10551 29084 10563 29087
rect 12176 29084 12204 29192
rect 13722 29180 13728 29192
rect 13780 29220 13786 29232
rect 15212 29220 15240 29251
rect 15470 29248 15476 29260
rect 15528 29248 15534 29300
rect 16022 29248 16028 29300
rect 16080 29288 16086 29300
rect 16945 29291 17003 29297
rect 16945 29288 16957 29291
rect 16080 29260 16957 29288
rect 16080 29248 16086 29260
rect 16945 29257 16957 29260
rect 16991 29288 17003 29291
rect 17402 29288 17408 29300
rect 16991 29260 17408 29288
rect 16991 29257 17003 29260
rect 16945 29251 17003 29257
rect 17402 29248 17408 29260
rect 17460 29288 17466 29300
rect 18690 29288 18696 29300
rect 17460 29260 18696 29288
rect 17460 29248 17466 29260
rect 18690 29248 18696 29260
rect 18748 29288 18754 29300
rect 20438 29288 20444 29300
rect 18748 29260 20444 29288
rect 18748 29248 18754 29260
rect 20438 29248 20444 29260
rect 20496 29248 20502 29300
rect 20622 29288 20628 29300
rect 20583 29260 20628 29288
rect 20622 29248 20628 29260
rect 20680 29248 20686 29300
rect 22278 29288 22284 29300
rect 20916 29260 22284 29288
rect 13780 29192 15240 29220
rect 13780 29180 13786 29192
rect 15562 29180 15568 29232
rect 15620 29220 15626 29232
rect 17497 29223 17555 29229
rect 17497 29220 17509 29223
rect 15620 29192 17509 29220
rect 15620 29180 15626 29192
rect 17497 29189 17509 29192
rect 17543 29220 17555 29223
rect 20916 29220 20944 29260
rect 22278 29248 22284 29260
rect 22336 29248 22342 29300
rect 22370 29248 22376 29300
rect 22428 29288 22434 29300
rect 22428 29260 22508 29288
rect 22428 29248 22434 29260
rect 17543 29192 20944 29220
rect 17543 29189 17555 29192
rect 17497 29183 17555 29189
rect 21450 29186 21456 29232
rect 21376 29180 21456 29186
rect 21508 29180 21514 29232
rect 22480 29229 22508 29260
rect 22554 29248 22560 29300
rect 22612 29288 22618 29300
rect 25409 29291 25467 29297
rect 22612 29260 25360 29288
rect 22612 29248 22618 29260
rect 22465 29223 22523 29229
rect 22465 29189 22477 29223
rect 22511 29189 22523 29223
rect 23569 29223 23627 29229
rect 23569 29220 23581 29223
rect 22465 29183 22523 29189
rect 22572 29192 23581 29220
rect 21376 29171 21494 29180
rect 21361 29165 21494 29171
rect 15838 29112 15844 29164
rect 15896 29152 15902 29164
rect 17770 29152 17776 29164
rect 15896 29124 17776 29152
rect 15896 29112 15902 29124
rect 17770 29112 17776 29124
rect 17828 29112 17834 29164
rect 18046 29152 18052 29164
rect 18007 29124 18052 29152
rect 18046 29112 18052 29124
rect 18104 29112 18110 29164
rect 18230 29112 18236 29164
rect 18288 29152 18294 29164
rect 19061 29155 19119 29161
rect 19061 29152 19073 29155
rect 18288 29124 19073 29152
rect 18288 29112 18294 29124
rect 19061 29121 19073 29124
rect 19107 29152 19119 29155
rect 19242 29152 19248 29164
rect 19107 29124 19248 29152
rect 19107 29121 19119 29124
rect 19061 29115 19119 29121
rect 19242 29112 19248 29124
rect 19300 29112 19306 29164
rect 19886 29152 19892 29164
rect 19847 29124 19892 29152
rect 19886 29112 19892 29124
rect 19944 29112 19950 29164
rect 19981 29155 20039 29161
rect 19981 29121 19993 29155
rect 20027 29121 20039 29155
rect 19981 29115 20039 29121
rect 10551 29056 12204 29084
rect 10551 29053 10563 29056
rect 10505 29047 10563 29053
rect 14366 29044 14372 29096
rect 14424 29084 14430 29096
rect 14645 29087 14703 29093
rect 14645 29084 14657 29087
rect 14424 29056 14657 29084
rect 14424 29044 14430 29056
rect 14645 29053 14657 29056
rect 14691 29084 14703 29087
rect 16758 29084 16764 29096
rect 14691 29056 16764 29084
rect 14691 29053 14703 29056
rect 14645 29047 14703 29053
rect 16758 29044 16764 29056
rect 16816 29044 16822 29096
rect 17034 29044 17040 29096
rect 17092 29084 17098 29096
rect 19996 29084 20024 29115
rect 20070 29112 20076 29164
rect 20128 29152 20134 29164
rect 20128 29124 20173 29152
rect 20128 29112 20134 29124
rect 20438 29112 20444 29164
rect 20496 29152 20502 29164
rect 20533 29155 20591 29161
rect 20533 29152 20545 29155
rect 20496 29124 20545 29152
rect 20496 29112 20502 29124
rect 20533 29121 20545 29124
rect 20579 29121 20591 29155
rect 20533 29115 20591 29121
rect 20714 29112 20720 29164
rect 20772 29152 20778 29164
rect 21177 29158 21235 29161
rect 20916 29155 21235 29158
rect 20916 29152 21189 29155
rect 20772 29130 21189 29152
rect 20772 29124 20944 29130
rect 20772 29112 20778 29124
rect 21177 29121 21189 29130
rect 21223 29121 21235 29155
rect 21361 29131 21373 29165
rect 21407 29158 21494 29165
rect 21407 29131 21419 29158
rect 21361 29125 21419 29131
rect 22112 29150 22324 29156
rect 22572 29150 22600 29192
rect 23569 29189 23581 29192
rect 23615 29189 23627 29223
rect 24397 29223 24455 29229
rect 24397 29220 24409 29223
rect 23569 29183 23627 29189
rect 24136 29192 24409 29220
rect 22112 29128 22600 29150
rect 21177 29115 21235 29121
rect 21269 29087 21327 29093
rect 21269 29084 21281 29087
rect 17092 29056 20024 29084
rect 20364 29056 21281 29084
rect 17092 29044 17098 29056
rect 9950 29016 9956 29028
rect 9911 28988 9956 29016
rect 9950 28976 9956 28988
rect 10008 28976 10014 29028
rect 11149 29019 11207 29025
rect 11149 28985 11161 29019
rect 11195 29016 11207 29019
rect 11330 29016 11336 29028
rect 11195 28988 11336 29016
rect 11195 28985 11207 28988
rect 11149 28979 11207 28985
rect 11330 28976 11336 28988
rect 11388 28976 11394 29028
rect 12989 29019 13047 29025
rect 12989 28985 13001 29019
rect 13035 29016 13047 29019
rect 14734 29016 14740 29028
rect 13035 28988 14740 29016
rect 13035 28985 13047 28988
rect 12989 28979 13047 28985
rect 14734 28976 14740 28988
rect 14792 28976 14798 29028
rect 15562 28976 15568 29028
rect 15620 29016 15626 29028
rect 16206 29016 16212 29028
rect 15620 28988 15884 29016
rect 16167 28988 16212 29016
rect 15620 28976 15626 28988
rect 13541 28951 13599 28957
rect 13541 28917 13553 28951
rect 13587 28948 13599 28951
rect 13630 28948 13636 28960
rect 13587 28920 13636 28948
rect 13587 28917 13599 28920
rect 13541 28911 13599 28917
rect 13630 28908 13636 28920
rect 13688 28908 13694 28960
rect 14093 28951 14151 28957
rect 14093 28917 14105 28951
rect 14139 28948 14151 28951
rect 14182 28948 14188 28960
rect 14139 28920 14188 28948
rect 14139 28917 14151 28920
rect 14093 28911 14151 28917
rect 14182 28908 14188 28920
rect 14240 28908 14246 28960
rect 15746 28948 15752 28960
rect 15707 28920 15752 28948
rect 15746 28908 15752 28920
rect 15804 28908 15810 28960
rect 15856 28948 15884 28988
rect 16206 28976 16212 28988
rect 16264 28976 16270 29028
rect 17218 28976 17224 29028
rect 17276 29016 17282 29028
rect 18509 29019 18567 29025
rect 18509 29016 18521 29019
rect 17276 28988 18521 29016
rect 17276 28976 17282 28988
rect 18509 28985 18521 28988
rect 18555 28985 18567 29019
rect 18509 28979 18567 28985
rect 18782 28976 18788 29028
rect 18840 29016 18846 29028
rect 20254 29016 20260 29028
rect 18840 28988 20260 29016
rect 18840 28976 18846 28988
rect 20254 28976 20260 28988
rect 20312 28976 20318 29028
rect 20364 28948 20392 29056
rect 21269 29053 21281 29056
rect 21315 29053 21327 29087
rect 22112 29084 22140 29128
rect 22296 29122 22600 29128
rect 22649 29155 22707 29161
rect 22649 29121 22661 29155
rect 22695 29152 22707 29155
rect 22738 29152 22744 29164
rect 22695 29124 22744 29152
rect 22695 29121 22707 29124
rect 22649 29115 22707 29121
rect 22664 29084 22692 29115
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 23290 29112 23296 29164
rect 23348 29152 23354 29164
rect 23348 29124 23393 29152
rect 23348 29112 23354 29124
rect 23658 29112 23664 29164
rect 23716 29152 23722 29164
rect 24026 29152 24032 29164
rect 23716 29124 23761 29152
rect 23828 29124 24032 29152
rect 23716 29112 23722 29124
rect 23477 29087 23535 29093
rect 21269 29047 21327 29053
rect 21578 29056 22140 29084
rect 22296 29056 22692 29084
rect 22848 29056 23440 29084
rect 21082 28976 21088 29028
rect 21140 29016 21146 29028
rect 21140 28988 21312 29016
rect 21140 28976 21146 28988
rect 15856 28920 20392 28948
rect 21284 28948 21312 28988
rect 21578 28948 21606 29056
rect 22296 29028 22324 29056
rect 22186 28976 22192 29028
rect 22244 28976 22250 29028
rect 22278 28976 22284 29028
rect 22336 28976 22342 29028
rect 22848 29025 22876 29056
rect 22833 29019 22891 29025
rect 22833 28985 22845 29019
rect 22879 28985 22891 29019
rect 23290 29016 23296 29028
rect 23251 28988 23296 29016
rect 22833 28979 22891 28985
rect 23290 28976 23296 28988
rect 23348 28976 23354 29028
rect 23412 29016 23440 29056
rect 23477 29053 23489 29087
rect 23523 29084 23535 29087
rect 23828 29084 23856 29124
rect 24026 29112 24032 29124
rect 24084 29112 24090 29164
rect 24136 29084 24164 29192
rect 24397 29189 24409 29192
rect 24443 29189 24455 29223
rect 24397 29183 24455 29189
rect 24688 29164 24716 29260
rect 25222 29220 25228 29232
rect 24872 29192 25228 29220
rect 24302 29112 24308 29164
rect 24360 29152 24366 29164
rect 24581 29155 24639 29161
rect 24581 29152 24593 29155
rect 24360 29124 24593 29152
rect 24360 29112 24366 29124
rect 24581 29121 24593 29124
rect 24627 29121 24639 29155
rect 24581 29115 24639 29121
rect 24670 29112 24676 29164
rect 24728 29152 24734 29164
rect 24872 29161 24900 29192
rect 25222 29180 25228 29192
rect 25280 29180 25286 29232
rect 25332 29220 25360 29260
rect 25409 29257 25421 29291
rect 25455 29288 25467 29291
rect 26326 29288 26332 29300
rect 25455 29260 26332 29288
rect 25455 29257 25467 29260
rect 25409 29251 25467 29257
rect 26326 29248 26332 29260
rect 26384 29248 26390 29300
rect 26605 29291 26663 29297
rect 26605 29257 26617 29291
rect 26651 29288 26663 29291
rect 27982 29288 27988 29300
rect 26651 29260 27988 29288
rect 26651 29257 26663 29260
rect 26605 29251 26663 29257
rect 27982 29248 27988 29260
rect 28040 29248 28046 29300
rect 28258 29248 28264 29300
rect 28316 29248 28322 29300
rect 28442 29248 28448 29300
rect 28500 29248 28506 29300
rect 28626 29248 28632 29300
rect 28684 29288 28690 29300
rect 28905 29291 28963 29297
rect 28905 29288 28917 29291
rect 28684 29260 28917 29288
rect 28684 29248 28690 29260
rect 28905 29257 28917 29260
rect 28951 29288 28963 29291
rect 30190 29288 30196 29300
rect 28951 29260 29500 29288
rect 30151 29260 30196 29288
rect 28951 29257 28963 29260
rect 28905 29251 28963 29257
rect 25593 29223 25651 29229
rect 25593 29220 25605 29223
rect 25332 29192 25605 29220
rect 25593 29189 25605 29192
rect 25639 29189 25651 29223
rect 25593 29183 25651 29189
rect 25866 29180 25872 29232
rect 25924 29220 25930 29232
rect 25924 29192 27292 29220
rect 25924 29180 25930 29192
rect 24857 29155 24915 29161
rect 24728 29124 24821 29152
rect 24728 29112 24734 29124
rect 24857 29121 24869 29155
rect 24903 29121 24915 29155
rect 24857 29115 24915 29121
rect 24946 29112 24952 29164
rect 25004 29152 25010 29164
rect 25004 29124 25049 29152
rect 25004 29112 25010 29124
rect 25130 29112 25136 29164
rect 25188 29152 25194 29164
rect 25188 29124 25652 29152
rect 25188 29112 25194 29124
rect 24394 29084 24400 29096
rect 23523 29056 23856 29084
rect 23952 29056 24164 29084
rect 24228 29056 24400 29084
rect 23523 29053 23535 29056
rect 23477 29047 23535 29053
rect 23566 29016 23572 29028
rect 23412 28988 23572 29016
rect 23566 28976 23572 28988
rect 23624 28976 23630 29028
rect 23658 28976 23664 29028
rect 23716 29016 23722 29028
rect 23952 29016 23980 29056
rect 23716 28988 23980 29016
rect 23716 28976 23722 28988
rect 24026 28976 24032 29028
rect 24084 29016 24090 29028
rect 24228 29016 24256 29056
rect 24394 29044 24400 29056
rect 24452 29084 24458 29096
rect 25222 29084 25228 29096
rect 24452 29056 25228 29084
rect 24452 29044 24458 29056
rect 25222 29044 25228 29056
rect 25280 29044 25286 29096
rect 25624 29084 25652 29124
rect 25682 29112 25688 29164
rect 25740 29152 25746 29164
rect 26421 29155 26479 29161
rect 26421 29152 26433 29155
rect 25740 29124 26433 29152
rect 25740 29112 25746 29124
rect 26421 29121 26433 29124
rect 26467 29121 26479 29155
rect 26421 29115 26479 29121
rect 26510 29112 26516 29164
rect 26568 29152 26574 29164
rect 26605 29155 26663 29161
rect 26605 29152 26617 29155
rect 26568 29124 26617 29152
rect 26568 29112 26574 29124
rect 26605 29121 26617 29124
rect 26651 29121 26663 29155
rect 26970 29152 26976 29164
rect 26605 29115 26663 29121
rect 26712 29124 26976 29152
rect 25961 29087 26019 29093
rect 25961 29084 25973 29087
rect 25624 29056 25973 29084
rect 25961 29053 25973 29056
rect 26007 29053 26019 29087
rect 25961 29047 26019 29053
rect 26326 29044 26332 29096
rect 26384 29084 26390 29096
rect 26712 29084 26740 29124
rect 26970 29112 26976 29124
rect 27028 29152 27034 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 27028 29124 27169 29152
rect 27028 29112 27034 29124
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 27264 29152 27292 29192
rect 27522 29180 27528 29232
rect 27580 29220 27586 29232
rect 28077 29223 28135 29229
rect 28077 29220 28089 29223
rect 27580 29192 28089 29220
rect 27580 29180 27586 29192
rect 28077 29189 28089 29192
rect 28123 29189 28135 29223
rect 28077 29183 28135 29189
rect 28276 29161 28304 29248
rect 28460 29164 28488 29248
rect 29472 29220 29500 29260
rect 30190 29248 30196 29260
rect 30248 29248 30254 29300
rect 32398 29220 32404 29232
rect 28644 29192 29408 29220
rect 29472 29192 32404 29220
rect 27985 29155 28043 29161
rect 27264 29124 27844 29152
rect 27157 29115 27215 29121
rect 26384 29056 26740 29084
rect 26384 29044 26390 29056
rect 26786 29044 26792 29096
rect 26844 29084 26850 29096
rect 27249 29087 27307 29093
rect 27249 29084 27261 29087
rect 26844 29056 27261 29084
rect 26844 29044 26850 29056
rect 27249 29053 27261 29056
rect 27295 29053 27307 29087
rect 27614 29084 27620 29096
rect 27249 29047 27307 29053
rect 27356 29056 27620 29084
rect 24084 28988 24256 29016
rect 24084 28976 24090 28988
rect 24302 28976 24308 29028
rect 24360 29016 24366 29028
rect 26142 29016 26148 29028
rect 24360 28988 26148 29016
rect 24360 28976 24366 28988
rect 26142 28976 26148 28988
rect 26200 28976 26206 29028
rect 26418 28976 26424 29028
rect 26476 29016 26482 29028
rect 26694 29016 26700 29028
rect 26476 28988 26700 29016
rect 26476 28976 26482 28988
rect 26694 28976 26700 28988
rect 26752 28976 26758 29028
rect 27062 28976 27068 29028
rect 27120 29016 27126 29028
rect 27356 29016 27384 29056
rect 27614 29044 27620 29056
rect 27672 29044 27678 29096
rect 27706 29044 27712 29096
rect 27764 29044 27770 29096
rect 27120 28988 27384 29016
rect 27120 28976 27126 28988
rect 27430 28976 27436 29028
rect 27488 29016 27494 29028
rect 27525 29019 27583 29025
rect 27525 29016 27537 29019
rect 27488 28988 27537 29016
rect 27488 28976 27494 28988
rect 27525 28985 27537 28988
rect 27571 28985 27583 29019
rect 27525 28979 27583 28985
rect 21284 28920 21606 28948
rect 22204 28948 22232 28976
rect 24394 28948 24400 28960
rect 22204 28920 24400 28948
rect 24394 28908 24400 28920
rect 24452 28908 24458 28960
rect 25314 28908 25320 28960
rect 25372 28948 25378 28960
rect 25593 28951 25651 28957
rect 25593 28948 25605 28951
rect 25372 28920 25605 28948
rect 25372 28908 25378 28920
rect 25593 28917 25605 28920
rect 25639 28917 25651 28951
rect 25593 28911 25651 28917
rect 26510 28908 26516 28960
rect 26568 28948 26574 28960
rect 26786 28948 26792 28960
rect 26568 28920 26792 28948
rect 26568 28908 26574 28920
rect 26786 28908 26792 28920
rect 26844 28908 26850 28960
rect 26970 28908 26976 28960
rect 27028 28948 27034 28960
rect 27246 28948 27252 28960
rect 27028 28920 27252 28948
rect 27028 28908 27034 28920
rect 27246 28908 27252 28920
rect 27304 28908 27310 28960
rect 27341 28951 27399 28957
rect 27341 28917 27353 28951
rect 27387 28948 27399 28951
rect 27614 28948 27620 28960
rect 27387 28920 27620 28948
rect 27387 28917 27399 28920
rect 27341 28911 27399 28917
rect 27614 28908 27620 28920
rect 27672 28948 27678 28960
rect 27724 28948 27752 29044
rect 27816 29016 27844 29124
rect 27985 29121 27997 29155
rect 28031 29121 28043 29155
rect 27985 29115 28043 29121
rect 28261 29155 28319 29161
rect 28261 29121 28273 29155
rect 28307 29121 28319 29155
rect 28261 29115 28319 29121
rect 28000 29016 28028 29115
rect 28350 29112 28356 29164
rect 28408 29112 28414 29164
rect 28442 29112 28448 29164
rect 28500 29112 28506 29164
rect 27816 28988 28028 29016
rect 28261 29019 28319 29025
rect 28261 28985 28273 29019
rect 28307 29016 28319 29019
rect 28368 29016 28396 29112
rect 28644 29096 28672 29192
rect 29380 29161 29408 29192
rect 32398 29180 32404 29192
rect 32456 29180 32462 29232
rect 28721 29155 28779 29161
rect 28721 29121 28733 29155
rect 28767 29121 28779 29155
rect 28721 29115 28779 29121
rect 28905 29155 28963 29161
rect 28905 29121 28917 29155
rect 28951 29152 28963 29155
rect 29365 29155 29423 29161
rect 28951 29124 29040 29152
rect 28951 29121 28963 29124
rect 28905 29115 28963 29121
rect 28626 29044 28632 29096
rect 28684 29044 28690 29096
rect 28736 29084 28764 29115
rect 29012 29084 29040 29124
rect 29365 29121 29377 29155
rect 29411 29121 29423 29155
rect 29365 29115 29423 29121
rect 29454 29112 29460 29164
rect 29512 29152 29518 29164
rect 29549 29155 29607 29161
rect 29549 29152 29561 29155
rect 29512 29124 29561 29152
rect 29512 29112 29518 29124
rect 29549 29121 29561 29124
rect 29595 29152 29607 29155
rect 29822 29152 29828 29164
rect 29595 29124 29828 29152
rect 29595 29121 29607 29124
rect 29549 29115 29607 29121
rect 29822 29112 29828 29124
rect 29880 29112 29886 29164
rect 30006 29152 30012 29164
rect 29967 29124 30012 29152
rect 30006 29112 30012 29124
rect 30064 29112 30070 29164
rect 30374 29112 30380 29164
rect 30432 29152 30438 29164
rect 31021 29155 31079 29161
rect 31021 29152 31033 29155
rect 30432 29124 31033 29152
rect 30432 29112 30438 29124
rect 31021 29121 31033 29124
rect 31067 29121 31079 29155
rect 31021 29115 31079 29121
rect 32858 29084 32864 29096
rect 28736 29056 28948 29084
rect 29012 29056 32864 29084
rect 28920 29028 28948 29056
rect 29380 29028 29408 29056
rect 32858 29044 32864 29056
rect 32916 29044 32922 29096
rect 28307 28988 28396 29016
rect 28307 28985 28319 28988
rect 28261 28979 28319 28985
rect 28902 28976 28908 29028
rect 28960 28976 28966 29028
rect 29362 28976 29368 29028
rect 29420 28976 29426 29028
rect 29457 29019 29515 29025
rect 29457 28985 29469 29019
rect 29503 29016 29515 29019
rect 29730 29016 29736 29028
rect 29503 28988 29736 29016
rect 29503 28985 29515 28988
rect 29457 28979 29515 28985
rect 29730 28976 29736 28988
rect 29788 28976 29794 29028
rect 31202 29016 31208 29028
rect 31163 28988 31208 29016
rect 31202 28976 31208 28988
rect 31260 28976 31266 29028
rect 28810 28948 28816 28960
rect 27672 28920 28816 28948
rect 27672 28908 27678 28920
rect 28810 28908 28816 28920
rect 28868 28908 28874 28960
rect 29178 28908 29184 28960
rect 29236 28948 29242 28960
rect 30190 28948 30196 28960
rect 29236 28920 30196 28948
rect 29236 28908 29242 28920
rect 30190 28908 30196 28920
rect 30248 28908 30254 28960
rect 1104 28858 31832 28880
rect 1104 28806 4791 28858
rect 4843 28806 4855 28858
rect 4907 28806 4919 28858
rect 4971 28806 4983 28858
rect 5035 28806 5047 28858
rect 5099 28806 12473 28858
rect 12525 28806 12537 28858
rect 12589 28806 12601 28858
rect 12653 28806 12665 28858
rect 12717 28806 12729 28858
rect 12781 28806 20155 28858
rect 20207 28806 20219 28858
rect 20271 28806 20283 28858
rect 20335 28806 20347 28858
rect 20399 28806 20411 28858
rect 20463 28806 27837 28858
rect 27889 28806 27901 28858
rect 27953 28806 27965 28858
rect 28017 28806 28029 28858
rect 28081 28806 28093 28858
rect 28145 28806 31832 28858
rect 1104 28784 31832 28806
rect 9858 28744 9864 28756
rect 9819 28716 9864 28744
rect 9858 28704 9864 28716
rect 9916 28704 9922 28756
rect 11790 28704 11796 28756
rect 11848 28744 11854 28756
rect 11977 28747 12035 28753
rect 11977 28744 11989 28747
rect 11848 28716 11989 28744
rect 11848 28704 11854 28716
rect 11977 28713 11989 28716
rect 12023 28713 12035 28747
rect 11977 28707 12035 28713
rect 12066 28704 12072 28756
rect 12124 28744 12130 28756
rect 12529 28747 12587 28753
rect 12529 28744 12541 28747
rect 12124 28716 12541 28744
rect 12124 28704 12130 28716
rect 12529 28713 12541 28716
rect 12575 28713 12587 28747
rect 12529 28707 12587 28713
rect 13725 28747 13783 28753
rect 13725 28713 13737 28747
rect 13771 28744 13783 28747
rect 13814 28744 13820 28756
rect 13771 28716 13820 28744
rect 13771 28713 13783 28716
rect 13725 28707 13783 28713
rect 6362 28636 6368 28688
rect 6420 28676 6426 28688
rect 11808 28676 11836 28704
rect 6420 28648 11836 28676
rect 6420 28636 6426 28648
rect 12434 28636 12440 28688
rect 12492 28676 12498 28688
rect 13740 28676 13768 28707
rect 13814 28704 13820 28716
rect 13872 28704 13878 28756
rect 15841 28747 15899 28753
rect 15841 28713 15853 28747
rect 15887 28744 15899 28747
rect 16022 28744 16028 28756
rect 15887 28716 16028 28744
rect 15887 28713 15899 28716
rect 15841 28707 15899 28713
rect 16022 28704 16028 28716
rect 16080 28704 16086 28756
rect 17126 28744 17132 28756
rect 17087 28716 17132 28744
rect 17126 28704 17132 28716
rect 17184 28704 17190 28756
rect 17402 28704 17408 28756
rect 17460 28744 17466 28756
rect 18046 28744 18052 28756
rect 17460 28716 18052 28744
rect 17460 28704 17466 28716
rect 18046 28704 18052 28716
rect 18104 28704 18110 28756
rect 18506 28704 18512 28756
rect 18564 28744 18570 28756
rect 20254 28744 20260 28756
rect 18564 28716 20260 28744
rect 18564 28704 18570 28716
rect 20254 28704 20260 28716
rect 20312 28704 20318 28756
rect 20349 28747 20407 28753
rect 20349 28713 20361 28747
rect 20395 28744 20407 28747
rect 20530 28744 20536 28756
rect 20395 28716 20536 28744
rect 20395 28713 20407 28716
rect 20349 28707 20407 28713
rect 20530 28704 20536 28716
rect 20588 28704 20594 28756
rect 21542 28704 21548 28756
rect 21600 28744 21606 28756
rect 22002 28744 22008 28756
rect 21600 28716 22008 28744
rect 21600 28704 21606 28716
rect 22002 28704 22008 28716
rect 22060 28704 22066 28756
rect 22833 28747 22891 28753
rect 22582 28716 22706 28744
rect 17586 28676 17592 28688
rect 12492 28648 13768 28676
rect 17547 28648 17592 28676
rect 12492 28636 12498 28648
rect 17586 28636 17592 28648
rect 17644 28636 17650 28688
rect 17770 28636 17776 28688
rect 17828 28676 17834 28688
rect 21269 28679 21327 28685
rect 21269 28676 21281 28679
rect 17828 28648 21281 28676
rect 17828 28636 17834 28648
rect 21269 28645 21281 28648
rect 21315 28645 21327 28679
rect 21269 28639 21327 28645
rect 21818 28636 21824 28688
rect 21876 28676 21882 28688
rect 22582 28676 22610 28716
rect 21876 28648 22610 28676
rect 22678 28676 22706 28716
rect 22833 28713 22845 28747
rect 22879 28744 22891 28747
rect 23106 28744 23112 28756
rect 22879 28716 23112 28744
rect 22879 28713 22891 28716
rect 22833 28707 22891 28713
rect 23106 28704 23112 28716
rect 23164 28704 23170 28756
rect 23198 28704 23204 28756
rect 23256 28744 23262 28756
rect 23382 28744 23388 28756
rect 23256 28716 23388 28744
rect 23256 28704 23262 28716
rect 23382 28704 23388 28716
rect 23440 28704 23446 28756
rect 23474 28704 23480 28756
rect 23532 28744 23538 28756
rect 23532 28716 23704 28744
rect 23532 28704 23538 28716
rect 22922 28676 22928 28688
rect 22678 28648 22928 28676
rect 21876 28636 21882 28648
rect 22922 28636 22928 28648
rect 22980 28676 22986 28688
rect 23566 28676 23572 28688
rect 22980 28648 23572 28676
rect 22980 28636 22986 28648
rect 23566 28636 23572 28648
rect 23624 28636 23630 28688
rect 7469 28611 7527 28617
rect 7469 28577 7481 28611
rect 7515 28608 7527 28611
rect 10873 28611 10931 28617
rect 10873 28608 10885 28611
rect 7515 28580 10885 28608
rect 7515 28577 7527 28580
rect 7469 28571 7527 28577
rect 10873 28577 10885 28580
rect 10919 28608 10931 28611
rect 19702 28608 19708 28620
rect 10919 28580 19708 28608
rect 10919 28577 10931 28580
rect 10873 28571 10931 28577
rect 19702 28568 19708 28580
rect 19760 28568 19766 28620
rect 20438 28608 20444 28620
rect 19812 28580 20444 28608
rect 1578 28540 1584 28552
rect 1539 28512 1584 28540
rect 1578 28500 1584 28512
rect 1636 28500 1642 28552
rect 8021 28543 8079 28549
rect 8021 28509 8033 28543
rect 8067 28540 8079 28543
rect 9030 28540 9036 28552
rect 8067 28512 9036 28540
rect 8067 28509 8079 28512
rect 8021 28503 8079 28509
rect 9030 28500 9036 28512
rect 9088 28500 9094 28552
rect 11054 28540 11060 28552
rect 9232 28512 11060 28540
rect 4154 28364 4160 28416
rect 4212 28404 4218 28416
rect 8481 28407 8539 28413
rect 8481 28404 8493 28407
rect 4212 28376 8493 28404
rect 4212 28364 4218 28376
rect 8481 28373 8493 28376
rect 8527 28404 8539 28407
rect 9232 28404 9260 28512
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 13170 28540 13176 28552
rect 13083 28512 13176 28540
rect 13170 28500 13176 28512
rect 13228 28540 13234 28552
rect 13228 28512 17954 28540
rect 13228 28500 13234 28512
rect 14182 28432 14188 28484
rect 14240 28472 14246 28484
rect 14737 28475 14795 28481
rect 14737 28472 14749 28475
rect 14240 28444 14749 28472
rect 14240 28432 14246 28444
rect 14737 28441 14749 28444
rect 14783 28472 14795 28475
rect 15746 28472 15752 28484
rect 14783 28444 15752 28472
rect 14783 28441 14795 28444
rect 14737 28435 14795 28441
rect 15746 28432 15752 28444
rect 15804 28432 15810 28484
rect 16850 28472 16856 28484
rect 15856 28444 16856 28472
rect 8527 28376 9260 28404
rect 9309 28407 9367 28413
rect 8527 28373 8539 28376
rect 8481 28367 8539 28373
rect 9309 28373 9321 28407
rect 9355 28404 9367 28407
rect 9398 28404 9404 28416
rect 9355 28376 9404 28404
rect 9355 28373 9367 28376
rect 9309 28367 9367 28373
rect 9398 28364 9404 28376
rect 9456 28364 9462 28416
rect 10410 28404 10416 28416
rect 10323 28376 10416 28404
rect 10410 28364 10416 28376
rect 10468 28404 10474 28416
rect 10870 28404 10876 28416
rect 10468 28376 10876 28404
rect 10468 28364 10474 28376
rect 10870 28364 10876 28376
rect 10928 28364 10934 28416
rect 11514 28404 11520 28416
rect 11475 28376 11520 28404
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 15194 28404 15200 28416
rect 15155 28376 15200 28404
rect 15194 28364 15200 28376
rect 15252 28364 15258 28416
rect 15286 28364 15292 28416
rect 15344 28404 15350 28416
rect 15856 28404 15884 28444
rect 16850 28432 16856 28444
rect 16908 28432 16914 28484
rect 17926 28472 17954 28512
rect 18230 28500 18236 28552
rect 18288 28540 18294 28552
rect 18690 28540 18696 28552
rect 18288 28512 18696 28540
rect 18288 28500 18294 28512
rect 18690 28500 18696 28512
rect 18748 28500 18754 28552
rect 19812 28540 19840 28580
rect 20438 28568 20444 28580
rect 20496 28568 20502 28620
rect 20714 28608 20720 28620
rect 20548 28580 20720 28608
rect 18797 28512 19840 28540
rect 19889 28543 19947 28549
rect 18797 28472 18825 28512
rect 19889 28509 19901 28543
rect 19935 28509 19947 28543
rect 19889 28503 19947 28509
rect 17926 28444 18825 28472
rect 19334 28432 19340 28484
rect 19392 28472 19398 28484
rect 19904 28472 19932 28503
rect 19978 28500 19984 28552
rect 20036 28540 20042 28552
rect 20548 28549 20576 28580
rect 20714 28568 20720 28580
rect 20772 28568 20778 28620
rect 20806 28568 20812 28620
rect 20864 28608 20870 28620
rect 21085 28611 21143 28617
rect 21085 28608 21097 28611
rect 20864 28580 21097 28608
rect 20864 28568 20870 28580
rect 21085 28577 21097 28580
rect 21131 28577 21143 28611
rect 23676 28608 23704 28716
rect 23750 28704 23756 28756
rect 23808 28744 23814 28756
rect 25590 28744 25596 28756
rect 23808 28716 25596 28744
rect 23808 28704 23814 28716
rect 25590 28704 25596 28716
rect 25648 28704 25654 28756
rect 25774 28744 25780 28756
rect 25735 28716 25780 28744
rect 25774 28704 25780 28716
rect 25832 28704 25838 28756
rect 25866 28704 25872 28756
rect 25924 28704 25930 28756
rect 26510 28704 26516 28756
rect 26568 28744 26574 28756
rect 26878 28744 26884 28756
rect 26568 28716 26884 28744
rect 26568 28704 26574 28716
rect 26878 28704 26884 28716
rect 26936 28704 26942 28756
rect 26970 28704 26976 28756
rect 27028 28744 27034 28756
rect 28353 28747 28411 28753
rect 28353 28744 28365 28747
rect 27028 28716 27073 28744
rect 27159 28716 28365 28744
rect 27028 28704 27034 28716
rect 23937 28679 23995 28685
rect 23937 28645 23949 28679
rect 23983 28676 23995 28679
rect 24578 28676 24584 28688
rect 23983 28648 24584 28676
rect 23983 28645 23995 28648
rect 23937 28639 23995 28645
rect 24578 28636 24584 28648
rect 24636 28676 24642 28688
rect 24946 28676 24952 28688
rect 24636 28648 24952 28676
rect 24636 28636 24642 28648
rect 24946 28636 24952 28648
rect 25004 28636 25010 28688
rect 25038 28636 25044 28688
rect 25096 28676 25102 28688
rect 25133 28679 25191 28685
rect 25133 28676 25145 28679
rect 25096 28648 25145 28676
rect 25096 28636 25102 28648
rect 25133 28645 25145 28648
rect 25179 28645 25191 28679
rect 25884 28676 25912 28704
rect 25133 28639 25191 28645
rect 25332 28648 25912 28676
rect 26605 28679 26663 28685
rect 25332 28620 25360 28648
rect 26605 28645 26617 28679
rect 26651 28645 26663 28679
rect 26605 28639 26663 28645
rect 23753 28611 23811 28617
rect 23753 28608 23765 28611
rect 21085 28571 21143 28577
rect 21284 28580 23440 28608
rect 23676 28580 23765 28608
rect 20533 28543 20591 28549
rect 20533 28540 20545 28543
rect 20036 28512 20545 28540
rect 20036 28500 20042 28512
rect 20533 28509 20545 28512
rect 20579 28509 20591 28543
rect 20533 28503 20591 28509
rect 20625 28543 20683 28549
rect 20625 28509 20637 28543
rect 20671 28540 20683 28543
rect 21284 28540 21312 28580
rect 23412 28574 23440 28580
rect 23753 28577 23765 28580
rect 23799 28577 23811 28611
rect 24118 28608 24124 28620
rect 20671 28512 21312 28540
rect 21361 28543 21419 28549
rect 20671 28509 20683 28512
rect 20625 28503 20683 28509
rect 21361 28509 21373 28543
rect 21407 28540 21419 28543
rect 21910 28540 21916 28552
rect 21407 28512 21916 28540
rect 21407 28509 21419 28512
rect 21361 28503 21419 28509
rect 21910 28500 21916 28512
rect 21968 28500 21974 28552
rect 22186 28540 22192 28552
rect 22099 28512 22192 28540
rect 22186 28500 22192 28512
rect 22244 28542 22250 28552
rect 22244 28540 22265 28542
rect 22244 28512 22508 28540
rect 22244 28500 22250 28512
rect 20346 28472 20352 28484
rect 19392 28444 19932 28472
rect 20307 28444 20352 28472
rect 19392 28432 19398 28444
rect 20346 28432 20352 28444
rect 20404 28432 20410 28484
rect 20438 28432 20444 28484
rect 20496 28472 20502 28484
rect 21085 28475 21143 28481
rect 21085 28472 21097 28475
rect 20496 28444 21097 28472
rect 20496 28432 20502 28444
rect 21085 28441 21097 28444
rect 21131 28441 21143 28475
rect 21085 28435 21143 28441
rect 21174 28432 21180 28484
rect 21232 28472 21238 28484
rect 21450 28472 21456 28484
rect 21232 28444 21456 28472
rect 21232 28432 21238 28444
rect 21450 28432 21456 28444
rect 21508 28432 21514 28484
rect 22005 28475 22063 28481
rect 22005 28441 22017 28475
rect 22051 28472 22063 28475
rect 22480 28472 22508 28512
rect 22554 28500 22560 28552
rect 22612 28540 22618 28552
rect 23412 28546 23474 28574
rect 23753 28571 23811 28577
rect 23952 28580 24124 28608
rect 22756 28540 22892 28542
rect 22612 28514 22892 28540
rect 23032 28540 23152 28542
rect 23446 28540 23474 28546
rect 23952 28540 23980 28580
rect 24118 28568 24124 28580
rect 24176 28568 24182 28620
rect 24210 28568 24216 28620
rect 24268 28608 24274 28620
rect 24673 28611 24731 28617
rect 24673 28608 24685 28611
rect 24268 28580 24685 28608
rect 24268 28568 24274 28580
rect 24673 28577 24685 28580
rect 24719 28577 24731 28611
rect 24673 28571 24731 28577
rect 24857 28611 24915 28617
rect 24857 28577 24869 28611
rect 24903 28608 24915 28611
rect 25314 28608 25320 28620
rect 24903 28580 25320 28608
rect 24903 28577 24915 28580
rect 24857 28571 24915 28577
rect 25314 28568 25320 28580
rect 25372 28568 25378 28620
rect 25590 28568 25596 28620
rect 25648 28568 25654 28620
rect 25774 28568 25780 28620
rect 25832 28608 25838 28620
rect 25869 28611 25927 28617
rect 25869 28608 25881 28611
rect 25832 28580 25881 28608
rect 25832 28568 25838 28580
rect 25869 28577 25881 28580
rect 25915 28577 25927 28611
rect 26620 28608 26648 28639
rect 26786 28636 26792 28688
rect 26844 28676 26850 28688
rect 27159 28676 27187 28716
rect 28353 28713 28365 28716
rect 28399 28713 28411 28747
rect 28721 28747 28779 28753
rect 28353 28707 28411 28713
rect 28460 28716 28672 28744
rect 28460 28676 28488 28716
rect 26844 28648 27187 28676
rect 27392 28648 28488 28676
rect 28644 28676 28672 28716
rect 28721 28713 28733 28747
rect 28767 28744 28779 28747
rect 31386 28744 31392 28756
rect 28767 28716 31392 28744
rect 28767 28713 28779 28716
rect 28721 28707 28779 28713
rect 31386 28704 31392 28716
rect 31444 28704 31450 28756
rect 30006 28676 30012 28688
rect 28644 28648 30012 28676
rect 26844 28636 26850 28648
rect 27392 28608 27420 28648
rect 30006 28636 30012 28648
rect 30064 28636 30070 28688
rect 29086 28608 29092 28620
rect 26620 28580 27420 28608
rect 27451 28580 28212 28608
rect 25869 28571 25927 28577
rect 23032 28518 23244 28540
rect 22612 28512 22784 28514
rect 22612 28500 22618 28512
rect 22649 28475 22707 28481
rect 22051 28444 22140 28472
rect 22480 28444 22607 28472
rect 22051 28441 22063 28444
rect 22005 28435 22063 28441
rect 22112 28416 22140 28444
rect 15344 28376 15884 28404
rect 16577 28407 16635 28413
rect 15344 28364 15350 28376
rect 16577 28373 16589 28407
rect 16623 28404 16635 28407
rect 16666 28404 16672 28416
rect 16623 28376 16672 28404
rect 16623 28373 16635 28376
rect 16577 28367 16635 28373
rect 16666 28364 16672 28376
rect 16724 28364 16730 28416
rect 17954 28364 17960 28416
rect 18012 28404 18018 28416
rect 18141 28407 18199 28413
rect 18141 28404 18153 28407
rect 18012 28376 18153 28404
rect 18012 28364 18018 28376
rect 18141 28373 18153 28376
rect 18187 28373 18199 28407
rect 18141 28367 18199 28373
rect 18785 28407 18843 28413
rect 18785 28373 18797 28407
rect 18831 28404 18843 28407
rect 19610 28404 19616 28416
rect 18831 28376 19616 28404
rect 18831 28373 18843 28376
rect 18785 28367 18843 28373
rect 19610 28364 19616 28376
rect 19668 28364 19674 28416
rect 19797 28407 19855 28413
rect 19797 28373 19809 28407
rect 19843 28404 19855 28407
rect 20714 28404 20720 28416
rect 19843 28376 20720 28404
rect 19843 28373 19855 28376
rect 19797 28367 19855 28373
rect 20714 28364 20720 28376
rect 20772 28364 20778 28416
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 21358 28404 21364 28416
rect 20864 28376 21364 28404
rect 20864 28364 20870 28376
rect 21358 28364 21364 28376
rect 21416 28364 21422 28416
rect 21542 28364 21548 28416
rect 21600 28404 21606 28416
rect 21821 28407 21879 28413
rect 21821 28404 21833 28407
rect 21600 28376 21833 28404
rect 21600 28364 21606 28376
rect 21821 28373 21833 28376
rect 21867 28373 21879 28407
rect 21821 28367 21879 28373
rect 22094 28364 22100 28416
rect 22152 28404 22158 28416
rect 22278 28404 22284 28416
rect 22152 28376 22284 28404
rect 22152 28364 22158 28376
rect 22278 28364 22284 28376
rect 22336 28364 22342 28416
rect 22579 28404 22607 28444
rect 22649 28441 22661 28475
rect 22695 28472 22707 28475
rect 22738 28472 22744 28484
rect 22695 28444 22744 28472
rect 22695 28441 22707 28444
rect 22649 28435 22707 28441
rect 22738 28432 22744 28444
rect 22796 28432 22802 28484
rect 22864 28481 22892 28514
rect 22940 28514 23244 28518
rect 22940 28490 23060 28514
rect 23124 28512 23244 28514
rect 23446 28512 23980 28540
rect 24029 28543 24087 28549
rect 23216 28506 23244 28512
rect 24029 28509 24041 28543
rect 24075 28540 24087 28543
rect 24578 28540 24584 28552
rect 24075 28512 24584 28540
rect 24075 28509 24087 28512
rect 22849 28475 22907 28481
rect 22849 28441 22861 28475
rect 22895 28441 22907 28475
rect 22849 28435 22907 28441
rect 22940 28404 22968 28490
rect 23216 28478 23416 28506
rect 24029 28503 24087 28509
rect 24578 28500 24584 28512
rect 24636 28500 24642 28552
rect 24762 28540 24768 28552
rect 24723 28512 24768 28540
rect 24762 28500 24768 28512
rect 24820 28500 24826 28552
rect 24949 28543 25007 28549
rect 24949 28509 24961 28543
rect 24995 28540 25007 28543
rect 25406 28540 25412 28552
rect 24995 28512 25412 28540
rect 24995 28509 25007 28512
rect 24949 28503 25007 28509
rect 25406 28500 25412 28512
rect 25464 28500 25470 28552
rect 25608 28540 25636 28568
rect 26145 28543 26203 28549
rect 25608 28512 26004 28540
rect 23388 28472 23416 28478
rect 23934 28472 23940 28484
rect 23388 28444 23940 28472
rect 23934 28432 23940 28444
rect 23992 28432 23998 28484
rect 24118 28432 24124 28484
rect 24176 28472 24182 28484
rect 25774 28472 25780 28484
rect 24176 28444 25780 28472
rect 24176 28432 24182 28444
rect 25774 28432 25780 28444
rect 25832 28432 25838 28484
rect 23033 28413 23039 28416
rect 22579 28376 22968 28404
rect 23017 28407 23039 28413
rect 23017 28373 23029 28407
rect 23017 28367 23039 28373
rect 23033 28364 23039 28367
rect 23091 28364 23097 28416
rect 23566 28404 23572 28416
rect 23527 28376 23572 28404
rect 23566 28364 23572 28376
rect 23624 28364 23630 28416
rect 23750 28364 23756 28416
rect 23808 28404 23814 28416
rect 25593 28407 25651 28413
rect 25593 28404 25605 28407
rect 23808 28376 25605 28404
rect 23808 28364 23814 28376
rect 25593 28373 25605 28376
rect 25639 28373 25651 28407
rect 25593 28367 25651 28373
rect 25682 28364 25688 28416
rect 25740 28404 25746 28416
rect 25866 28404 25872 28416
rect 25740 28376 25872 28404
rect 25740 28364 25746 28376
rect 25866 28364 25872 28376
rect 25924 28364 25930 28416
rect 25976 28404 26004 28512
rect 26145 28509 26157 28543
rect 26191 28540 26203 28543
rect 26234 28540 26240 28552
rect 26191 28512 26240 28540
rect 26191 28509 26203 28512
rect 26145 28503 26203 28509
rect 26234 28500 26240 28512
rect 26292 28500 26298 28552
rect 26786 28540 26792 28552
rect 26747 28512 26792 28540
rect 26786 28500 26792 28512
rect 26844 28500 26850 28552
rect 26881 28543 26939 28549
rect 26881 28509 26893 28543
rect 26927 28509 26939 28543
rect 26881 28503 26939 28509
rect 27065 28543 27123 28549
rect 27065 28509 27077 28543
rect 27111 28540 27123 28543
rect 27451 28540 27479 28580
rect 27111 28512 27479 28540
rect 27525 28543 27583 28549
rect 27111 28509 27123 28512
rect 27065 28503 27123 28509
rect 27525 28509 27537 28543
rect 27571 28540 27583 28543
rect 27798 28540 27804 28552
rect 27571 28512 27804 28540
rect 27571 28509 27583 28512
rect 27525 28503 27583 28509
rect 26896 28472 26924 28503
rect 27540 28472 27568 28503
rect 27798 28500 27804 28512
rect 27856 28500 27862 28552
rect 28184 28542 28212 28580
rect 28376 28580 29092 28608
rect 28258 28542 28264 28552
rect 28184 28514 28264 28542
rect 28258 28500 28264 28514
rect 28316 28500 28322 28552
rect 28376 28549 28404 28580
rect 29086 28568 29092 28580
rect 29144 28568 29150 28620
rect 28358 28543 28416 28549
rect 28358 28509 28370 28543
rect 28404 28509 28416 28543
rect 28358 28503 28416 28509
rect 28537 28543 28595 28549
rect 28537 28509 28549 28543
rect 28583 28540 28595 28543
rect 29454 28540 29460 28552
rect 28583 28512 29460 28540
rect 28583 28509 28595 28512
rect 28537 28503 28595 28509
rect 29454 28500 29460 28512
rect 29512 28500 29518 28552
rect 29917 28543 29975 28549
rect 29917 28509 29929 28543
rect 29963 28540 29975 28543
rect 30006 28540 30012 28552
rect 29963 28512 30012 28540
rect 29963 28509 29975 28512
rect 29917 28503 29975 28509
rect 30006 28500 30012 28512
rect 30064 28500 30070 28552
rect 30377 28543 30435 28549
rect 30377 28509 30389 28543
rect 30423 28509 30435 28543
rect 30377 28503 30435 28509
rect 27706 28472 27712 28484
rect 26896 28444 27568 28472
rect 27667 28444 27712 28472
rect 27706 28432 27712 28444
rect 27764 28432 27770 28484
rect 27890 28472 27896 28484
rect 27851 28444 27896 28472
rect 27890 28432 27896 28444
rect 27948 28432 27954 28484
rect 29178 28472 29184 28484
rect 28460 28444 29184 28472
rect 26878 28404 26884 28416
rect 25976 28376 26884 28404
rect 26878 28364 26884 28376
rect 26936 28364 26942 28416
rect 27062 28364 27068 28416
rect 27120 28404 27126 28416
rect 27614 28404 27620 28416
rect 27120 28376 27620 28404
rect 27120 28364 27126 28376
rect 27614 28364 27620 28376
rect 27672 28364 27678 28416
rect 28258 28364 28264 28416
rect 28316 28404 28322 28416
rect 28460 28404 28488 28444
rect 29178 28432 29184 28444
rect 29236 28432 29242 28484
rect 30392 28472 30420 28503
rect 30558 28500 30564 28552
rect 30616 28540 30622 28552
rect 31021 28543 31079 28549
rect 31021 28540 31033 28543
rect 30616 28512 31033 28540
rect 30616 28500 30622 28512
rect 31021 28509 31033 28512
rect 31067 28509 31079 28543
rect 31021 28503 31079 28509
rect 31294 28500 31300 28552
rect 31352 28500 31358 28552
rect 31312 28472 31340 28500
rect 32398 28472 32404 28484
rect 30392 28444 32404 28472
rect 32398 28432 32404 28444
rect 32456 28432 32462 28484
rect 28316 28376 28488 28404
rect 28316 28364 28322 28376
rect 28534 28364 28540 28416
rect 28592 28404 28598 28416
rect 28994 28404 29000 28416
rect 28592 28376 29000 28404
rect 28592 28364 28598 28376
rect 28994 28364 29000 28376
rect 29052 28364 29058 28416
rect 29086 28364 29092 28416
rect 29144 28404 29150 28416
rect 29454 28404 29460 28416
rect 29144 28376 29460 28404
rect 29144 28364 29150 28376
rect 29454 28364 29460 28376
rect 29512 28364 29518 28416
rect 29822 28404 29828 28416
rect 29783 28376 29828 28404
rect 29822 28364 29828 28376
rect 29880 28364 29886 28416
rect 30374 28364 30380 28416
rect 30432 28404 30438 28416
rect 30469 28407 30527 28413
rect 30469 28404 30481 28407
rect 30432 28376 30481 28404
rect 30432 28364 30438 28376
rect 30469 28373 30481 28376
rect 30515 28373 30527 28407
rect 30469 28367 30527 28373
rect 31205 28407 31263 28413
rect 31205 28373 31217 28407
rect 31251 28404 31263 28407
rect 31294 28404 31300 28416
rect 31251 28376 31300 28404
rect 31251 28373 31263 28376
rect 31205 28367 31263 28373
rect 31294 28364 31300 28376
rect 31352 28364 31358 28416
rect 1104 28314 31992 28336
rect 1104 28262 8632 28314
rect 8684 28262 8696 28314
rect 8748 28262 8760 28314
rect 8812 28262 8824 28314
rect 8876 28262 8888 28314
rect 8940 28262 16314 28314
rect 16366 28262 16378 28314
rect 16430 28262 16442 28314
rect 16494 28262 16506 28314
rect 16558 28262 16570 28314
rect 16622 28262 23996 28314
rect 24048 28262 24060 28314
rect 24112 28262 24124 28314
rect 24176 28262 24188 28314
rect 24240 28262 24252 28314
rect 24304 28262 31678 28314
rect 31730 28262 31742 28314
rect 31794 28262 31806 28314
rect 31858 28262 31870 28314
rect 31922 28262 31934 28314
rect 31986 28262 31992 28314
rect 1104 28240 31992 28262
rect 7285 28203 7343 28209
rect 7285 28169 7297 28203
rect 7331 28200 7343 28203
rect 9582 28200 9588 28212
rect 7331 28172 9588 28200
rect 7331 28169 7343 28172
rect 7285 28163 7343 28169
rect 9582 28160 9588 28172
rect 9640 28160 9646 28212
rect 13909 28203 13967 28209
rect 13909 28169 13921 28203
rect 13955 28200 13967 28203
rect 14550 28200 14556 28212
rect 13955 28172 14556 28200
rect 13955 28169 13967 28172
rect 13909 28163 13967 28169
rect 14550 28160 14556 28172
rect 14608 28160 14614 28212
rect 14734 28200 14740 28212
rect 14695 28172 14740 28200
rect 14734 28160 14740 28172
rect 14792 28160 14798 28212
rect 15289 28203 15347 28209
rect 15289 28169 15301 28203
rect 15335 28200 15347 28203
rect 15378 28200 15384 28212
rect 15335 28172 15384 28200
rect 15335 28169 15347 28172
rect 15289 28163 15347 28169
rect 15378 28160 15384 28172
rect 15436 28160 15442 28212
rect 15930 28160 15936 28212
rect 15988 28200 15994 28212
rect 16209 28203 16267 28209
rect 16209 28200 16221 28203
rect 15988 28172 16221 28200
rect 15988 28160 15994 28172
rect 16209 28169 16221 28172
rect 16255 28169 16267 28203
rect 16209 28163 16267 28169
rect 18417 28203 18475 28209
rect 18417 28169 18429 28203
rect 18463 28200 18475 28203
rect 18598 28200 18604 28212
rect 18463 28172 18604 28200
rect 18463 28169 18475 28172
rect 18417 28163 18475 28169
rect 18598 28160 18604 28172
rect 18656 28160 18662 28212
rect 18690 28160 18696 28212
rect 18748 28200 18754 28212
rect 19061 28203 19119 28209
rect 19061 28200 19073 28203
rect 18748 28172 19073 28200
rect 18748 28160 18754 28172
rect 19061 28169 19073 28172
rect 19107 28169 19119 28203
rect 19061 28163 19119 28169
rect 19150 28160 19156 28212
rect 19208 28200 19214 28212
rect 19334 28200 19340 28212
rect 19208 28172 19340 28200
rect 19208 28160 19214 28172
rect 19334 28160 19340 28172
rect 19392 28160 19398 28212
rect 19610 28160 19616 28212
rect 19668 28200 19674 28212
rect 21174 28200 21180 28212
rect 19668 28172 21180 28200
rect 19668 28160 19674 28172
rect 21174 28160 21180 28172
rect 21232 28160 21238 28212
rect 21361 28203 21419 28209
rect 21361 28169 21373 28203
rect 21407 28200 21419 28203
rect 21818 28200 21824 28212
rect 21407 28172 21824 28200
rect 21407 28169 21419 28172
rect 21361 28163 21419 28169
rect 21818 28160 21824 28172
rect 21876 28160 21882 28212
rect 23474 28200 23480 28212
rect 22848 28172 23480 28200
rect 9493 28135 9551 28141
rect 9493 28101 9505 28135
rect 9539 28132 9551 28135
rect 11422 28132 11428 28144
rect 9539 28104 11428 28132
rect 9539 28101 9551 28104
rect 9493 28095 9551 28101
rect 11422 28092 11428 28104
rect 11480 28132 11486 28144
rect 11974 28132 11980 28144
rect 11480 28104 11980 28132
rect 11480 28092 11486 28104
rect 11974 28092 11980 28104
rect 12032 28092 12038 28144
rect 12802 28132 12808 28144
rect 12763 28104 12808 28132
rect 12802 28092 12808 28104
rect 12860 28092 12866 28144
rect 13262 28132 13268 28144
rect 13175 28104 13268 28132
rect 13262 28092 13268 28104
rect 13320 28132 13326 28144
rect 14918 28132 14924 28144
rect 13320 28104 14924 28132
rect 13320 28092 13326 28104
rect 14918 28092 14924 28104
rect 14976 28092 14982 28144
rect 16574 28092 16580 28144
rect 16632 28132 16638 28144
rect 17218 28132 17224 28144
rect 16632 28104 17224 28132
rect 16632 28092 16638 28104
rect 17218 28092 17224 28104
rect 17276 28092 17282 28144
rect 20441 28135 20499 28141
rect 20441 28132 20453 28135
rect 18429 28104 20453 28132
rect 13354 28024 13360 28076
rect 13412 28064 13418 28076
rect 18313 28067 18371 28073
rect 18313 28064 18325 28067
rect 13412 28036 18325 28064
rect 13412 28024 13418 28036
rect 18313 28033 18325 28036
rect 18359 28033 18371 28067
rect 18313 28027 18371 28033
rect 10502 27956 10508 28008
rect 10560 27996 10566 28008
rect 12161 27999 12219 28005
rect 12161 27996 12173 27999
rect 10560 27968 12173 27996
rect 10560 27956 10566 27968
rect 12161 27965 12173 27968
rect 12207 27996 12219 27999
rect 13906 27996 13912 28008
rect 12207 27968 13912 27996
rect 12207 27965 12219 27968
rect 12161 27959 12219 27965
rect 13906 27956 13912 27968
rect 13964 27996 13970 28008
rect 14366 27996 14372 28008
rect 13964 27968 14372 27996
rect 13964 27956 13970 27968
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 18429 27996 18457 28104
rect 20441 28101 20453 28104
rect 20487 28101 20499 28135
rect 22005 28135 22063 28141
rect 22005 28132 22017 28135
rect 20441 28095 20499 28101
rect 20732 28104 22017 28132
rect 18509 28067 18567 28073
rect 18509 28033 18521 28067
rect 18555 28064 18567 28067
rect 18782 28064 18788 28076
rect 18555 28036 18788 28064
rect 18555 28033 18567 28036
rect 18509 28027 18567 28033
rect 18782 28024 18788 28036
rect 18840 28024 18846 28076
rect 18972 28073 18978 28076
rect 18969 28027 18978 28073
rect 19030 28064 19036 28076
rect 19030 28036 19069 28064
rect 18972 28024 18978 28027
rect 19030 28024 19036 28036
rect 19150 28024 19156 28076
rect 19208 28064 19214 28076
rect 19208 28036 19253 28064
rect 19208 28024 19214 28036
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 19705 28067 19763 28073
rect 19705 28064 19717 28067
rect 19392 28036 19717 28064
rect 19392 28024 19398 28036
rect 19705 28033 19717 28036
rect 19751 28064 19763 28067
rect 20254 28064 20260 28076
rect 19751 28036 20260 28064
rect 19751 28033 19763 28036
rect 19705 28027 19763 28033
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20349 28067 20407 28073
rect 20349 28033 20361 28067
rect 20395 28064 20407 28067
rect 20530 28064 20536 28076
rect 20395 28036 20536 28064
rect 20395 28033 20407 28036
rect 20349 28027 20407 28033
rect 20530 28024 20536 28036
rect 20588 28024 20594 28076
rect 20625 28067 20683 28073
rect 20625 28033 20637 28067
rect 20671 28033 20683 28067
rect 20625 28027 20683 28033
rect 19168 27996 19196 28024
rect 14608 27968 18457 27996
rect 18511 27968 19196 27996
rect 14608 27956 14614 27968
rect 8294 27888 8300 27940
rect 8352 27928 8358 27940
rect 8849 27931 8907 27937
rect 8849 27928 8861 27931
rect 8352 27900 8861 27928
rect 8352 27888 8358 27900
rect 8849 27897 8861 27900
rect 8895 27897 8907 27931
rect 8849 27891 8907 27897
rect 10597 27931 10655 27937
rect 10597 27897 10609 27931
rect 10643 27928 10655 27931
rect 11330 27928 11336 27940
rect 10643 27900 11336 27928
rect 10643 27897 10655 27900
rect 10597 27891 10655 27897
rect 11330 27888 11336 27900
rect 11388 27888 11394 27940
rect 11790 27888 11796 27940
rect 11848 27928 11854 27940
rect 11974 27928 11980 27940
rect 11848 27900 11980 27928
rect 11848 27888 11854 27900
rect 11974 27888 11980 27900
rect 12032 27928 12038 27940
rect 15286 27928 15292 27940
rect 12032 27900 15292 27928
rect 12032 27888 12038 27900
rect 15286 27888 15292 27900
rect 15344 27888 15350 27940
rect 15746 27888 15752 27940
rect 15804 27928 15810 27940
rect 18511 27928 18539 27968
rect 19610 27956 19616 28008
rect 19668 27996 19674 28008
rect 19668 27968 20024 27996
rect 19668 27956 19674 27968
rect 19794 27928 19800 27940
rect 15804 27900 18539 27928
rect 18616 27900 19800 27928
rect 15804 27888 15810 27900
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 7837 27863 7895 27869
rect 7837 27829 7849 27863
rect 7883 27860 7895 27863
rect 8110 27860 8116 27872
rect 7883 27832 8116 27860
rect 7883 27829 7895 27832
rect 7837 27823 7895 27829
rect 8110 27820 8116 27832
rect 8168 27820 8174 27872
rect 8386 27860 8392 27872
rect 8347 27832 8392 27860
rect 8386 27820 8392 27832
rect 8444 27820 8450 27872
rect 9674 27820 9680 27872
rect 9732 27860 9738 27872
rect 9953 27863 10011 27869
rect 9953 27860 9965 27863
rect 9732 27832 9965 27860
rect 9732 27820 9738 27832
rect 9953 27829 9965 27832
rect 9999 27829 10011 27863
rect 9953 27823 10011 27829
rect 11149 27863 11207 27869
rect 11149 27829 11161 27863
rect 11195 27860 11207 27863
rect 11238 27860 11244 27872
rect 11195 27832 11244 27860
rect 11195 27829 11207 27832
rect 11149 27823 11207 27829
rect 11238 27820 11244 27832
rect 11296 27820 11302 27872
rect 12066 27820 12072 27872
rect 12124 27860 12130 27872
rect 12802 27860 12808 27872
rect 12124 27832 12808 27860
rect 12124 27820 12130 27832
rect 12802 27820 12808 27832
rect 12860 27820 12866 27872
rect 15102 27820 15108 27872
rect 15160 27860 15166 27872
rect 15654 27860 15660 27872
rect 15160 27832 15660 27860
rect 15160 27820 15166 27832
rect 15654 27820 15660 27832
rect 15712 27860 15718 27872
rect 17773 27863 17831 27869
rect 17773 27860 17785 27863
rect 15712 27832 17785 27860
rect 15712 27820 15718 27832
rect 17773 27829 17785 27832
rect 17819 27860 17831 27863
rect 18616 27860 18644 27900
rect 19794 27888 19800 27900
rect 19852 27928 19858 27940
rect 19889 27931 19947 27937
rect 19889 27928 19901 27931
rect 19852 27900 19901 27928
rect 19852 27888 19858 27900
rect 19889 27897 19901 27900
rect 19935 27897 19947 27931
rect 19996 27928 20024 27968
rect 20070 27956 20076 28008
rect 20128 27996 20134 28008
rect 20640 27996 20668 28027
rect 20128 27968 20668 27996
rect 20128 27956 20134 27968
rect 20625 27931 20683 27937
rect 20625 27928 20637 27931
rect 19996 27900 20637 27928
rect 19889 27891 19947 27897
rect 20625 27897 20637 27900
rect 20671 27928 20683 27931
rect 20732 27928 20760 28104
rect 22005 28101 22017 28104
rect 22051 28101 22063 28135
rect 22186 28132 22192 28144
rect 22147 28104 22192 28132
rect 22005 28095 22063 28101
rect 22186 28092 22192 28104
rect 22244 28092 22250 28144
rect 22278 28092 22284 28144
rect 22336 28132 22342 28144
rect 22848 28132 22876 28172
rect 23474 28160 23480 28172
rect 23532 28160 23538 28212
rect 23658 28160 23664 28212
rect 23716 28200 23722 28212
rect 24029 28203 24087 28209
rect 24029 28200 24041 28203
rect 23716 28172 24041 28200
rect 23716 28160 23722 28172
rect 24029 28169 24041 28172
rect 24075 28169 24087 28203
rect 24029 28163 24087 28169
rect 24121 28203 24179 28209
rect 24121 28169 24133 28203
rect 24167 28200 24179 28203
rect 24210 28200 24216 28212
rect 24167 28172 24216 28200
rect 24167 28169 24179 28172
rect 24121 28163 24179 28169
rect 24210 28160 24216 28172
rect 24268 28160 24274 28212
rect 27982 28200 27988 28212
rect 24320 28172 27988 28200
rect 22336 28104 22876 28132
rect 22336 28092 22342 28104
rect 20806 28024 20812 28076
rect 20864 28064 20870 28076
rect 21085 28067 21143 28073
rect 21085 28064 21097 28067
rect 20864 28036 21097 28064
rect 20864 28024 20870 28036
rect 21085 28033 21097 28036
rect 21131 28033 21143 28067
rect 21085 28027 21143 28033
rect 21269 28067 21327 28073
rect 21269 28033 21281 28067
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 20898 27956 20904 28008
rect 20956 27996 20962 28008
rect 21284 27996 21312 28027
rect 21634 28024 21640 28076
rect 21692 28064 21698 28076
rect 22738 28064 22744 28076
rect 21692 28036 22744 28064
rect 21692 28024 21698 28036
rect 22738 28024 22744 28036
rect 22796 28024 22802 28076
rect 22848 28073 22876 28104
rect 23566 28092 23572 28144
rect 23624 28132 23630 28144
rect 23934 28132 23940 28144
rect 23624 28104 23940 28132
rect 23624 28092 23630 28104
rect 23934 28092 23940 28104
rect 23992 28092 23998 28144
rect 24320 28132 24348 28172
rect 27982 28160 27988 28172
rect 28040 28160 28046 28212
rect 28166 28200 28172 28212
rect 28127 28172 28172 28200
rect 28166 28160 28172 28172
rect 28224 28160 28230 28212
rect 30193 28203 30251 28209
rect 28376 28172 30144 28200
rect 24044 28104 24348 28132
rect 22833 28067 22891 28073
rect 22833 28033 22845 28067
rect 22879 28033 22891 28067
rect 22833 28027 22891 28033
rect 22925 28067 22983 28073
rect 22925 28033 22937 28067
rect 22971 28033 22983 28067
rect 22925 28027 22983 28033
rect 20956 27968 21312 27996
rect 20956 27956 20962 27968
rect 21818 27956 21824 28008
rect 21876 27996 21882 28008
rect 22940 27996 22968 28027
rect 23014 28024 23020 28076
rect 23072 28073 23078 28076
rect 23072 28067 23094 28073
rect 23082 28033 23094 28067
rect 23198 28064 23204 28076
rect 23159 28036 23204 28064
rect 23072 28027 23094 28033
rect 23072 28024 23078 28027
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 23385 28067 23443 28073
rect 23385 28033 23397 28067
rect 23431 28064 23443 28067
rect 24044 28064 24072 28104
rect 24394 28092 24400 28144
rect 24452 28132 24458 28144
rect 25406 28132 25412 28144
rect 24452 28104 25412 28132
rect 24452 28092 24458 28104
rect 25406 28092 25412 28104
rect 25464 28092 25470 28144
rect 26602 28132 26608 28144
rect 25516 28104 26608 28132
rect 23431 28036 24072 28064
rect 23431 28033 23443 28036
rect 23385 28027 23443 28033
rect 24118 28024 24124 28076
rect 24176 28064 24182 28076
rect 24213 28067 24271 28073
rect 24213 28064 24225 28067
rect 24176 28036 24225 28064
rect 24176 28024 24182 28036
rect 24213 28033 24225 28036
rect 24259 28033 24271 28067
rect 24213 28027 24271 28033
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28064 24915 28067
rect 24946 28064 24952 28076
rect 24903 28036 24952 28064
rect 24903 28033 24915 28036
rect 24857 28027 24915 28033
rect 24946 28024 24952 28036
rect 25004 28024 25010 28076
rect 25222 28064 25228 28076
rect 25183 28036 25228 28064
rect 25222 28024 25228 28036
rect 25280 28024 25286 28076
rect 25516 28064 25544 28104
rect 26602 28092 26608 28104
rect 26660 28092 26666 28144
rect 26694 28092 26700 28144
rect 26752 28132 26758 28144
rect 28376 28132 28404 28172
rect 28810 28132 28816 28144
rect 26752 28104 27384 28132
rect 26752 28092 26758 28104
rect 26046 28064 26052 28076
rect 25332 28036 25544 28064
rect 26007 28036 26052 28064
rect 24394 27996 24400 28008
rect 21876 27968 22892 27996
rect 22940 27968 24400 27996
rect 21876 27956 21882 27968
rect 20671 27900 20760 27928
rect 20671 27897 20683 27900
rect 20625 27891 20683 27897
rect 21266 27888 21272 27940
rect 21324 27928 21330 27940
rect 22373 27931 22431 27937
rect 22373 27928 22385 27931
rect 21324 27900 22385 27928
rect 21324 27888 21330 27900
rect 22373 27897 22385 27900
rect 22419 27897 22431 27931
rect 22373 27891 22431 27897
rect 22554 27888 22560 27940
rect 22612 27888 22618 27940
rect 22864 27928 22892 27968
rect 24394 27956 24400 27968
rect 24452 27956 24458 28008
rect 24578 27956 24584 28008
rect 24636 27996 24642 28008
rect 25332 27996 25360 28036
rect 26046 28024 26052 28036
rect 26104 28024 26110 28076
rect 26142 28024 26148 28076
rect 26200 28064 26206 28076
rect 26330 28067 26388 28073
rect 26200 28036 26245 28064
rect 26200 28024 26206 28036
rect 26330 28033 26342 28067
rect 26376 28064 26388 28067
rect 26786 28064 26792 28076
rect 26376 28036 26792 28064
rect 26376 28033 26388 28036
rect 26330 28027 26388 28033
rect 26786 28024 26792 28036
rect 26844 28024 26850 28076
rect 26970 28024 26976 28076
rect 27028 28064 27034 28076
rect 27356 28073 27384 28104
rect 27448 28104 28404 28132
rect 28460 28104 28816 28132
rect 27448 28073 27476 28104
rect 27249 28067 27307 28073
rect 27249 28064 27261 28067
rect 27028 28036 27261 28064
rect 27028 28024 27034 28036
rect 27249 28033 27261 28036
rect 27295 28033 27307 28067
rect 27249 28027 27307 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28033 27399 28067
rect 27341 28027 27399 28033
rect 27433 28067 27491 28073
rect 27433 28033 27445 28067
rect 27479 28033 27491 28067
rect 27433 28027 27491 28033
rect 27614 28024 27620 28076
rect 27672 28064 27678 28076
rect 28074 28064 28080 28076
rect 27672 28036 28080 28064
rect 27672 28024 27678 28036
rect 28074 28024 28080 28036
rect 28132 28024 28138 28076
rect 28350 28064 28356 28076
rect 28311 28036 28356 28064
rect 28350 28024 28356 28036
rect 28408 28024 28414 28076
rect 28460 28073 28488 28104
rect 28810 28092 28816 28104
rect 28868 28092 28874 28144
rect 29270 28132 29276 28144
rect 29231 28104 29276 28132
rect 29270 28092 29276 28104
rect 29328 28092 29334 28144
rect 29454 28132 29460 28144
rect 29415 28104 29460 28132
rect 29454 28092 29460 28104
rect 29512 28092 29518 28144
rect 30116 28132 30144 28172
rect 30193 28169 30205 28203
rect 30239 28200 30251 28203
rect 30239 28172 30880 28200
rect 30239 28169 30251 28172
rect 30193 28163 30251 28169
rect 30742 28132 30748 28144
rect 30116 28104 30748 28132
rect 30742 28092 30748 28104
rect 30800 28092 30806 28144
rect 28445 28067 28503 28073
rect 28445 28033 28457 28067
rect 28491 28033 28503 28067
rect 28445 28027 28503 28033
rect 28629 28070 28687 28073
rect 28629 28067 28764 28070
rect 28629 28033 28641 28067
rect 28675 28042 28764 28067
rect 28675 28033 28687 28042
rect 28629 28027 28687 28033
rect 24636 27968 25360 27996
rect 24636 27956 24642 27968
rect 25406 27956 25412 28008
rect 25464 27996 25470 28008
rect 26237 27999 26295 28005
rect 26237 27996 26249 27999
rect 25464 27968 26249 27996
rect 25464 27956 25470 27968
rect 26237 27965 26249 27968
rect 26283 27965 26295 27999
rect 26237 27959 26295 27965
rect 22864 27900 23980 27928
rect 17819 27832 18644 27860
rect 17819 27829 17831 27832
rect 17773 27823 17831 27829
rect 19058 27820 19064 27872
rect 19116 27860 19122 27872
rect 22186 27860 22192 27872
rect 19116 27832 22192 27860
rect 19116 27820 19122 27832
rect 22186 27820 22192 27832
rect 22244 27820 22250 27872
rect 22572 27860 22600 27888
rect 23845 27863 23903 27869
rect 23845 27860 23857 27863
rect 22572 27832 23857 27860
rect 23845 27829 23857 27832
rect 23891 27829 23903 27863
rect 23952 27860 23980 27900
rect 24210 27888 24216 27940
rect 24268 27928 24274 27940
rect 24268 27900 25728 27928
rect 24268 27888 24274 27900
rect 24854 27860 24860 27872
rect 23952 27832 24860 27860
rect 23845 27823 23903 27829
rect 24854 27820 24860 27832
rect 24912 27820 24918 27872
rect 25222 27860 25228 27872
rect 25183 27832 25228 27860
rect 25222 27820 25228 27832
rect 25280 27820 25286 27872
rect 25409 27863 25467 27869
rect 25409 27829 25421 27863
rect 25455 27860 25467 27863
rect 25590 27860 25596 27872
rect 25455 27832 25596 27860
rect 25455 27829 25467 27832
rect 25409 27823 25467 27829
rect 25590 27820 25596 27832
rect 25648 27820 25654 27872
rect 25700 27860 25728 27900
rect 25774 27888 25780 27940
rect 25832 27928 25838 27940
rect 25869 27931 25927 27937
rect 25869 27928 25881 27931
rect 25832 27900 25881 27928
rect 25832 27888 25838 27900
rect 25869 27897 25881 27900
rect 25915 27897 25927 27931
rect 26252 27928 26280 27959
rect 26602 27956 26608 28008
rect 26660 27996 26666 28008
rect 27525 27999 27583 28005
rect 27525 27996 27537 27999
rect 26660 27968 27537 27996
rect 26660 27956 26666 27968
rect 27525 27965 27537 27968
rect 27571 27965 27583 27999
rect 27525 27959 27583 27965
rect 27798 27956 27804 28008
rect 27856 27996 27862 28008
rect 27856 27968 28580 27996
rect 27856 27956 27862 27968
rect 26252 27900 26832 27928
rect 25869 27891 25927 27897
rect 26804 27872 26832 27900
rect 26878 27888 26884 27940
rect 26936 27928 26942 27940
rect 26936 27900 28488 27928
rect 26936 27888 26942 27900
rect 28460 27872 28488 27900
rect 26694 27860 26700 27872
rect 25700 27832 26700 27860
rect 26694 27820 26700 27832
rect 26752 27820 26758 27872
rect 26786 27820 26792 27872
rect 26844 27820 26850 27872
rect 27430 27820 27436 27872
rect 27488 27860 27494 27872
rect 27709 27863 27767 27869
rect 27709 27860 27721 27863
rect 27488 27832 27721 27860
rect 27488 27820 27494 27832
rect 27709 27829 27721 27832
rect 27755 27829 27767 27863
rect 28442 27860 28448 27872
rect 28403 27832 28448 27860
rect 27709 27823 27767 27829
rect 28442 27820 28448 27832
rect 28500 27820 28506 27872
rect 28552 27860 28580 27968
rect 28736 27928 28764 28042
rect 29089 28067 29147 28073
rect 29089 28033 29101 28067
rect 29135 28064 29147 28067
rect 29546 28064 29552 28076
rect 29135 28036 29552 28064
rect 29135 28033 29147 28036
rect 29089 28027 29147 28033
rect 29546 28024 29552 28036
rect 29604 28064 29610 28076
rect 30006 28064 30012 28076
rect 29604 28036 30012 28064
rect 29604 28024 29610 28036
rect 30006 28024 30012 28036
rect 30064 28024 30070 28076
rect 30098 28024 30104 28076
rect 30156 28064 30162 28076
rect 30193 28067 30251 28073
rect 30193 28064 30205 28067
rect 30156 28036 30205 28064
rect 30156 28024 30162 28036
rect 30193 28033 30205 28036
rect 30239 28033 30251 28067
rect 30193 28027 30251 28033
rect 28810 27956 28816 28008
rect 28868 27996 28874 28008
rect 29917 27999 29975 28005
rect 29917 27996 29929 27999
rect 28868 27968 29929 27996
rect 28868 27956 28874 27968
rect 29917 27965 29929 27968
rect 29963 27996 29975 27999
rect 30282 27996 30288 28008
rect 29963 27968 30288 27996
rect 29963 27965 29975 27968
rect 29917 27959 29975 27965
rect 30282 27956 30288 27968
rect 30340 27956 30346 28008
rect 29822 27928 29828 27940
rect 28736 27900 29828 27928
rect 29822 27888 29828 27900
rect 29880 27888 29886 27940
rect 30101 27931 30159 27937
rect 30101 27897 30113 27931
rect 30147 27928 30159 27931
rect 30190 27928 30196 27940
rect 30147 27900 30196 27928
rect 30147 27897 30159 27900
rect 30101 27891 30159 27897
rect 30190 27888 30196 27900
rect 30248 27888 30254 27940
rect 30852 27928 30880 28172
rect 31018 28064 31024 28076
rect 30979 28036 31024 28064
rect 31018 28024 31024 28036
rect 31076 28024 31082 28076
rect 31018 27928 31024 27940
rect 30852 27900 31024 27928
rect 31018 27888 31024 27900
rect 31076 27888 31082 27940
rect 29454 27860 29460 27872
rect 28552 27832 29460 27860
rect 29454 27820 29460 27832
rect 29512 27820 29518 27872
rect 30282 27820 30288 27872
rect 30340 27860 30346 27872
rect 31205 27863 31263 27869
rect 31205 27860 31217 27863
rect 30340 27832 31217 27860
rect 30340 27820 30346 27832
rect 31205 27829 31217 27832
rect 31251 27829 31263 27863
rect 31205 27823 31263 27829
rect 1104 27770 31832 27792
rect 1104 27718 4791 27770
rect 4843 27718 4855 27770
rect 4907 27718 4919 27770
rect 4971 27718 4983 27770
rect 5035 27718 5047 27770
rect 5099 27718 12473 27770
rect 12525 27718 12537 27770
rect 12589 27718 12601 27770
rect 12653 27718 12665 27770
rect 12717 27718 12729 27770
rect 12781 27718 20155 27770
rect 20207 27718 20219 27770
rect 20271 27718 20283 27770
rect 20335 27718 20347 27770
rect 20399 27718 20411 27770
rect 20463 27718 27837 27770
rect 27889 27718 27901 27770
rect 27953 27718 27965 27770
rect 28017 27718 28029 27770
rect 28081 27718 28093 27770
rect 28145 27718 31832 27770
rect 1104 27696 31832 27718
rect 8386 27616 8392 27668
rect 8444 27656 8450 27668
rect 12986 27656 12992 27668
rect 8444 27628 12992 27656
rect 8444 27616 8450 27628
rect 12986 27616 12992 27628
rect 13044 27616 13050 27668
rect 14366 27616 14372 27668
rect 14424 27656 14430 27668
rect 15378 27656 15384 27668
rect 14424 27628 15384 27656
rect 14424 27616 14430 27628
rect 15378 27616 15384 27628
rect 15436 27616 15442 27668
rect 15746 27616 15752 27668
rect 15804 27656 15810 27668
rect 16574 27656 16580 27668
rect 15804 27628 16580 27656
rect 15804 27616 15810 27628
rect 16574 27616 16580 27628
rect 16632 27616 16638 27668
rect 16853 27659 16911 27665
rect 16853 27625 16865 27659
rect 16899 27656 16911 27659
rect 16942 27656 16948 27668
rect 16899 27628 16948 27656
rect 16899 27625 16911 27628
rect 16853 27619 16911 27625
rect 16942 27616 16948 27628
rect 17000 27656 17006 27668
rect 17402 27656 17408 27668
rect 17000 27628 17408 27656
rect 17000 27616 17006 27628
rect 17402 27616 17408 27628
rect 17460 27616 17466 27668
rect 17494 27616 17500 27668
rect 17552 27656 17558 27668
rect 17552 27628 17597 27656
rect 17552 27616 17558 27628
rect 17862 27616 17868 27668
rect 17920 27656 17926 27668
rect 19889 27659 19947 27665
rect 17920 27628 18920 27656
rect 17920 27616 17926 27628
rect 9030 27548 9036 27600
rect 9088 27588 9094 27600
rect 10042 27588 10048 27600
rect 9088 27560 10048 27588
rect 9088 27548 9094 27560
rect 10042 27548 10048 27560
rect 10100 27588 10106 27600
rect 11517 27591 11575 27597
rect 11517 27588 11529 27591
rect 10100 27560 11529 27588
rect 10100 27548 10106 27560
rect 11517 27557 11529 27560
rect 11563 27588 11575 27591
rect 11790 27588 11796 27600
rect 11563 27560 11796 27588
rect 11563 27557 11575 27560
rect 11517 27551 11575 27557
rect 11790 27548 11796 27560
rect 11848 27548 11854 27600
rect 12621 27591 12679 27597
rect 12621 27557 12633 27591
rect 12667 27588 12679 27591
rect 12894 27588 12900 27600
rect 12667 27560 12900 27588
rect 12667 27557 12679 27560
rect 12621 27551 12679 27557
rect 9309 27523 9367 27529
rect 9309 27489 9321 27523
rect 9355 27520 9367 27523
rect 10134 27520 10140 27532
rect 9355 27492 10140 27520
rect 9355 27489 9367 27492
rect 9309 27483 9367 27489
rect 10134 27480 10140 27492
rect 10192 27520 10198 27532
rect 10318 27520 10324 27532
rect 10192 27492 10324 27520
rect 10192 27480 10198 27492
rect 10318 27480 10324 27492
rect 10376 27480 10382 27532
rect 10410 27480 10416 27532
rect 10468 27520 10474 27532
rect 12636 27520 12664 27551
rect 12894 27548 12900 27560
rect 12952 27548 12958 27600
rect 13630 27588 13636 27600
rect 13004 27560 13636 27588
rect 13004 27520 13032 27560
rect 13630 27548 13636 27560
rect 13688 27588 13694 27600
rect 15657 27591 15715 27597
rect 15657 27588 15669 27591
rect 13688 27560 15669 27588
rect 13688 27548 13694 27560
rect 15657 27557 15669 27560
rect 15703 27588 15715 27591
rect 17954 27588 17960 27600
rect 15703 27560 17960 27588
rect 15703 27557 15715 27560
rect 15657 27551 15715 27557
rect 17954 27548 17960 27560
rect 18012 27548 18018 27600
rect 18049 27591 18107 27597
rect 18049 27557 18061 27591
rect 18095 27588 18107 27591
rect 18322 27588 18328 27600
rect 18095 27560 18328 27588
rect 18095 27557 18107 27560
rect 18049 27551 18107 27557
rect 18322 27548 18328 27560
rect 18380 27548 18386 27600
rect 18414 27548 18420 27600
rect 18472 27548 18478 27600
rect 18785 27591 18843 27597
rect 18785 27557 18797 27591
rect 18831 27588 18843 27591
rect 18892 27588 18920 27628
rect 19889 27625 19901 27659
rect 19935 27656 19947 27659
rect 20254 27656 20260 27668
rect 19935 27628 20260 27656
rect 19935 27625 19947 27628
rect 19889 27619 19947 27625
rect 20254 27616 20260 27628
rect 20312 27616 20318 27668
rect 20806 27616 20812 27668
rect 20864 27656 20870 27668
rect 21177 27659 21235 27665
rect 21177 27656 21189 27659
rect 20864 27628 21189 27656
rect 20864 27616 20870 27628
rect 21177 27625 21189 27628
rect 21223 27625 21235 27659
rect 21177 27619 21235 27625
rect 21266 27616 21272 27668
rect 21324 27656 21330 27668
rect 21542 27656 21548 27668
rect 21324 27628 21548 27656
rect 21324 27616 21330 27628
rect 21542 27616 21548 27628
rect 21600 27616 21606 27668
rect 21634 27616 21640 27668
rect 21692 27656 21698 27668
rect 21692 27628 22416 27656
rect 21692 27616 21698 27628
rect 18831 27560 18920 27588
rect 18831 27557 18843 27560
rect 18785 27551 18843 27557
rect 19334 27548 19340 27600
rect 19392 27588 19398 27600
rect 20070 27588 20076 27600
rect 19392 27560 20076 27588
rect 19392 27548 19398 27560
rect 20070 27548 20076 27560
rect 20128 27548 20134 27600
rect 22281 27591 22339 27597
rect 22281 27588 22293 27591
rect 21100 27560 22293 27588
rect 10468 27492 12664 27520
rect 12728 27492 13032 27520
rect 10468 27480 10474 27492
rect 11238 27412 11244 27464
rect 11296 27452 11302 27464
rect 12158 27452 12164 27464
rect 11296 27424 12164 27452
rect 11296 27412 11302 27424
rect 12158 27412 12164 27424
rect 12216 27452 12222 27464
rect 12728 27452 12756 27492
rect 13538 27480 13544 27532
rect 13596 27520 13602 27532
rect 13725 27523 13783 27529
rect 13725 27520 13737 27523
rect 13596 27492 13737 27520
rect 13596 27480 13602 27492
rect 13725 27489 13737 27492
rect 13771 27520 13783 27523
rect 14553 27523 14611 27529
rect 14553 27520 14565 27523
rect 13771 27492 14565 27520
rect 13771 27489 13783 27492
rect 13725 27483 13783 27489
rect 14553 27489 14565 27492
rect 14599 27520 14611 27523
rect 17034 27520 17040 27532
rect 14599 27492 17040 27520
rect 14599 27489 14611 27492
rect 14553 27483 14611 27489
rect 17034 27480 17040 27492
rect 17092 27480 17098 27532
rect 17586 27480 17592 27532
rect 17644 27520 17650 27532
rect 18432 27520 18460 27548
rect 18877 27523 18935 27529
rect 18877 27520 18889 27523
rect 17644 27492 18352 27520
rect 18432 27492 18889 27520
rect 17644 27480 17650 27492
rect 12216 27424 12756 27452
rect 12216 27412 12222 27424
rect 14182 27412 14188 27464
rect 14240 27452 14246 27464
rect 16114 27452 16120 27464
rect 14240 27424 16120 27452
rect 14240 27412 14246 27424
rect 16114 27412 16120 27424
rect 16172 27452 16178 27464
rect 16209 27455 16267 27461
rect 16209 27452 16221 27455
rect 16172 27424 16221 27452
rect 16172 27412 16178 27424
rect 16209 27421 16221 27424
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 17126 27412 17132 27464
rect 17184 27452 17190 27464
rect 17313 27455 17371 27461
rect 17313 27452 17325 27455
rect 17184 27424 17325 27452
rect 17184 27412 17190 27424
rect 17313 27421 17325 27424
rect 17359 27421 17371 27455
rect 17313 27415 17371 27421
rect 17497 27455 17555 27461
rect 17497 27421 17509 27455
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 17957 27455 18015 27461
rect 17957 27421 17969 27455
rect 18003 27452 18015 27455
rect 18230 27452 18236 27464
rect 18003 27424 18236 27452
rect 18003 27421 18015 27424
rect 17957 27415 18015 27421
rect 3878 27344 3884 27396
rect 3936 27384 3942 27396
rect 7374 27384 7380 27396
rect 3936 27356 7380 27384
rect 3936 27344 3942 27356
rect 7374 27344 7380 27356
rect 7432 27344 7438 27396
rect 8018 27384 8024 27396
rect 7979 27356 8024 27384
rect 8018 27344 8024 27356
rect 8076 27344 8082 27396
rect 10318 27344 10324 27396
rect 10376 27384 10382 27396
rect 12066 27384 12072 27396
rect 10376 27356 12072 27384
rect 10376 27344 10382 27356
rect 12066 27344 12072 27356
rect 12124 27344 12130 27396
rect 13998 27344 14004 27396
rect 14056 27384 14062 27396
rect 14826 27384 14832 27396
rect 14056 27356 14832 27384
rect 14056 27344 14062 27356
rect 14826 27344 14832 27356
rect 14884 27384 14890 27396
rect 15013 27387 15071 27393
rect 15013 27384 15025 27387
rect 14884 27356 15025 27384
rect 14884 27344 14890 27356
rect 15013 27353 15025 27356
rect 15059 27353 15071 27387
rect 15013 27347 15071 27353
rect 15654 27344 15660 27396
rect 15712 27384 15718 27396
rect 17512 27384 17540 27415
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 18324 27452 18352 27492
rect 18877 27489 18889 27492
rect 18923 27489 18935 27523
rect 18877 27483 18935 27489
rect 18984 27492 20668 27520
rect 18414 27452 18420 27464
rect 18324 27424 18420 27452
rect 18414 27412 18420 27424
rect 18472 27452 18478 27464
rect 18601 27455 18659 27461
rect 18472 27446 18555 27452
rect 18601 27446 18613 27455
rect 18472 27424 18613 27446
rect 18472 27412 18478 27424
rect 18527 27421 18613 27424
rect 18647 27421 18659 27455
rect 18527 27418 18659 27421
rect 18601 27415 18659 27418
rect 18690 27412 18696 27464
rect 18748 27452 18754 27464
rect 18748 27424 18793 27452
rect 18748 27412 18754 27424
rect 15712 27356 17540 27384
rect 15712 27344 15718 27356
rect 17586 27344 17592 27396
rect 17644 27384 17650 27396
rect 18984 27384 19012 27492
rect 19334 27412 19340 27464
rect 19392 27452 19398 27464
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 19392 27424 19625 27452
rect 19392 27412 19398 27424
rect 19613 27421 19625 27424
rect 19659 27421 19671 27455
rect 19886 27452 19892 27464
rect 19847 27424 19892 27452
rect 19613 27415 19671 27421
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 20254 27452 20260 27464
rect 20088 27424 20260 27452
rect 17644 27356 19012 27384
rect 19705 27387 19763 27393
rect 17644 27344 17650 27356
rect 19705 27353 19717 27387
rect 19751 27384 19763 27387
rect 20088 27384 20116 27424
rect 20254 27412 20260 27424
rect 20312 27412 20318 27464
rect 20533 27455 20591 27461
rect 20533 27421 20545 27455
rect 20579 27421 20591 27455
rect 20640 27452 20668 27492
rect 20714 27480 20720 27532
rect 20772 27520 20778 27532
rect 20772 27492 20817 27520
rect 20772 27480 20778 27492
rect 21100 27464 21128 27560
rect 22281 27557 22293 27560
rect 22327 27557 22339 27591
rect 22281 27551 22339 27557
rect 21266 27520 21272 27532
rect 21227 27492 21272 27520
rect 21266 27480 21272 27492
rect 21324 27480 21330 27532
rect 22388 27520 22416 27628
rect 22204 27492 22416 27520
rect 22678 27628 23416 27656
rect 20640 27424 21036 27452
rect 20533 27415 20591 27421
rect 19751 27356 20116 27384
rect 19751 27353 19763 27356
rect 19705 27347 19763 27353
rect 20162 27344 20168 27396
rect 20220 27384 20226 27396
rect 20349 27387 20407 27393
rect 20349 27384 20361 27387
rect 20220 27356 20361 27384
rect 20220 27344 20226 27356
rect 20349 27353 20361 27356
rect 20395 27353 20407 27387
rect 20349 27347 20407 27353
rect 6362 27316 6368 27328
rect 6323 27288 6368 27316
rect 6362 27276 6368 27288
rect 6420 27276 6426 27328
rect 6917 27319 6975 27325
rect 6917 27285 6929 27319
rect 6963 27316 6975 27319
rect 7282 27316 7288 27328
rect 6963 27288 7288 27316
rect 6963 27285 6975 27288
rect 6917 27279 6975 27285
rect 7282 27276 7288 27288
rect 7340 27276 7346 27328
rect 8573 27319 8631 27325
rect 8573 27285 8585 27319
rect 8619 27316 8631 27319
rect 9030 27316 9036 27328
rect 8619 27288 9036 27316
rect 8619 27285 8631 27288
rect 8573 27279 8631 27285
rect 9030 27276 9036 27288
rect 9088 27276 9094 27328
rect 9398 27276 9404 27328
rect 9456 27316 9462 27328
rect 9861 27319 9919 27325
rect 9861 27316 9873 27319
rect 9456 27288 9873 27316
rect 9456 27276 9462 27288
rect 9861 27285 9873 27288
rect 9907 27316 9919 27319
rect 10873 27319 10931 27325
rect 10873 27316 10885 27319
rect 9907 27288 10885 27316
rect 9907 27285 9919 27288
rect 9861 27279 9919 27285
rect 10873 27285 10885 27288
rect 10919 27285 10931 27319
rect 10873 27279 10931 27285
rect 11606 27276 11612 27328
rect 11664 27316 11670 27328
rect 11882 27316 11888 27328
rect 11664 27288 11888 27316
rect 11664 27276 11670 27288
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 13173 27319 13231 27325
rect 13173 27285 13185 27319
rect 13219 27316 13231 27319
rect 16758 27316 16764 27328
rect 13219 27288 16764 27316
rect 13219 27285 13231 27288
rect 13173 27279 13231 27285
rect 16758 27276 16764 27288
rect 16816 27276 16822 27328
rect 16850 27276 16856 27328
rect 16908 27316 16914 27328
rect 20548 27316 20576 27415
rect 16908 27288 20576 27316
rect 16908 27276 16914 27288
rect 20714 27276 20720 27328
rect 20772 27316 20778 27328
rect 20898 27316 20904 27328
rect 20772 27288 20904 27316
rect 20772 27276 20778 27288
rect 20898 27276 20904 27288
rect 20956 27276 20962 27328
rect 21008 27316 21036 27424
rect 21082 27412 21088 27464
rect 21140 27412 21146 27464
rect 21177 27455 21235 27461
rect 21177 27421 21189 27455
rect 21223 27452 21235 27455
rect 21223 27424 21312 27452
rect 21223 27421 21235 27424
rect 21177 27415 21235 27421
rect 21284 27396 21312 27424
rect 22204 27396 22232 27492
rect 22557 27455 22615 27461
rect 22557 27421 22569 27455
rect 22603 27452 22615 27455
rect 22678 27452 22706 27628
rect 22833 27591 22891 27597
rect 22833 27557 22845 27591
rect 22879 27588 22891 27591
rect 23290 27588 23296 27600
rect 22879 27560 23296 27588
rect 22879 27557 22891 27560
rect 22833 27551 22891 27557
rect 23290 27548 23296 27560
rect 23348 27548 23354 27600
rect 23388 27588 23416 27628
rect 23566 27616 23572 27668
rect 23624 27656 23630 27668
rect 24765 27659 24823 27665
rect 24765 27656 24777 27659
rect 23624 27628 24777 27656
rect 23624 27616 23630 27628
rect 24765 27625 24777 27628
rect 24811 27625 24823 27659
rect 24765 27619 24823 27625
rect 24854 27616 24860 27668
rect 24912 27656 24918 27668
rect 25590 27656 25596 27668
rect 24912 27628 25596 27656
rect 24912 27616 24918 27628
rect 25590 27616 25596 27628
rect 25648 27616 25654 27668
rect 26053 27659 26111 27665
rect 26053 27625 26065 27659
rect 26099 27656 26111 27659
rect 26142 27656 26148 27668
rect 26099 27628 26148 27656
rect 26099 27625 26111 27628
rect 26053 27619 26111 27625
rect 26142 27616 26148 27628
rect 26200 27616 26206 27668
rect 28905 27659 28963 27665
rect 26620 27628 27381 27656
rect 23388 27560 24900 27588
rect 22738 27480 22744 27532
rect 22796 27520 22802 27532
rect 24578 27520 24584 27532
rect 22796 27492 24584 27520
rect 22796 27480 22802 27492
rect 24578 27480 24584 27492
rect 24636 27480 24642 27532
rect 22603 27424 22706 27452
rect 22603 27421 22615 27424
rect 22557 27415 22615 27421
rect 23198 27412 23204 27464
rect 23256 27452 23262 27464
rect 23293 27455 23351 27461
rect 23293 27452 23305 27455
rect 23256 27424 23305 27452
rect 23256 27412 23262 27424
rect 23293 27421 23305 27424
rect 23339 27421 23351 27455
rect 23293 27415 23351 27421
rect 23385 27455 23443 27461
rect 23385 27421 23397 27455
rect 23431 27421 23443 27455
rect 23385 27415 23443 27421
rect 23569 27455 23627 27461
rect 23569 27421 23581 27455
rect 23615 27421 23627 27455
rect 23569 27415 23627 27421
rect 23661 27455 23719 27461
rect 23661 27421 23673 27455
rect 23707 27421 23719 27455
rect 23661 27415 23719 27421
rect 23845 27455 23903 27461
rect 23845 27421 23857 27455
rect 23891 27452 23903 27455
rect 24210 27452 24216 27464
rect 23891 27424 24216 27452
rect 23891 27421 23903 27424
rect 23845 27415 23903 27421
rect 21266 27344 21272 27396
rect 21324 27344 21330 27396
rect 21376 27356 22094 27384
rect 21376 27316 21404 27356
rect 21008 27288 21404 27316
rect 21545 27319 21603 27325
rect 21545 27285 21557 27319
rect 21591 27316 21603 27319
rect 21634 27316 21640 27328
rect 21591 27288 21640 27316
rect 21591 27285 21603 27288
rect 21545 27279 21603 27285
rect 21634 27276 21640 27288
rect 21692 27276 21698 27328
rect 22066 27316 22094 27356
rect 22186 27344 22192 27396
rect 22244 27344 22250 27396
rect 22278 27344 22284 27396
rect 22336 27384 22342 27396
rect 22336 27356 22692 27384
rect 22336 27344 22342 27356
rect 22664 27325 22692 27356
rect 22830 27344 22836 27396
rect 22888 27384 22894 27396
rect 23388 27384 23416 27415
rect 23584 27384 23612 27415
rect 22888 27356 23416 27384
rect 23446 27356 23612 27384
rect 22888 27344 22894 27356
rect 22465 27319 22523 27325
rect 22465 27316 22477 27319
rect 22066 27288 22477 27316
rect 22465 27285 22477 27288
rect 22511 27285 22523 27319
rect 22465 27279 22523 27285
rect 22649 27319 22707 27325
rect 22649 27285 22661 27319
rect 22695 27285 22707 27319
rect 22649 27279 22707 27285
rect 22922 27276 22928 27328
rect 22980 27316 22986 27328
rect 23446 27316 23474 27356
rect 22980 27288 23474 27316
rect 22980 27276 22986 27288
rect 23566 27276 23572 27328
rect 23624 27316 23630 27328
rect 23676 27316 23704 27415
rect 24210 27412 24216 27424
rect 24268 27412 24274 27464
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27421 24823 27455
rect 24872 27452 24900 27560
rect 26234 27548 26240 27600
rect 26292 27588 26298 27600
rect 26292 27560 26337 27588
rect 26292 27548 26298 27560
rect 24949 27523 25007 27529
rect 24949 27489 24961 27523
rect 24995 27520 25007 27523
rect 26620 27520 26648 27628
rect 26697 27591 26755 27597
rect 26697 27557 26709 27591
rect 26743 27588 26755 27591
rect 26878 27588 26884 27600
rect 26743 27560 26884 27588
rect 26743 27557 26755 27560
rect 26697 27551 26755 27557
rect 26878 27548 26884 27560
rect 26936 27548 26942 27600
rect 26970 27548 26976 27600
rect 27028 27588 27034 27600
rect 27249 27591 27307 27597
rect 27249 27588 27261 27591
rect 27028 27560 27261 27588
rect 27028 27548 27034 27560
rect 27249 27557 27261 27560
rect 27295 27557 27307 27591
rect 27353 27588 27381 27628
rect 27882 27628 28300 27656
rect 27882 27588 27910 27628
rect 27353 27560 27910 27588
rect 27985 27591 28043 27597
rect 27249 27551 27307 27557
rect 27985 27557 27997 27591
rect 28031 27588 28043 27591
rect 28272 27588 28300 27628
rect 28905 27625 28917 27659
rect 28951 27656 28963 27659
rect 29086 27656 29092 27668
rect 28951 27628 29092 27656
rect 28951 27625 28963 27628
rect 28905 27619 28963 27625
rect 29086 27616 29092 27628
rect 29144 27616 29150 27668
rect 29638 27616 29644 27668
rect 29696 27656 29702 27668
rect 29733 27659 29791 27665
rect 29733 27656 29745 27659
rect 29696 27628 29745 27656
rect 29696 27616 29702 27628
rect 29733 27625 29745 27628
rect 29779 27625 29791 27659
rect 29733 27619 29791 27625
rect 29917 27659 29975 27665
rect 29917 27625 29929 27659
rect 29963 27656 29975 27659
rect 30558 27656 30564 27668
rect 29963 27628 30564 27656
rect 29963 27625 29975 27628
rect 29917 27619 29975 27625
rect 30558 27616 30564 27628
rect 30616 27616 30622 27668
rect 30653 27591 30711 27597
rect 30653 27588 30665 27591
rect 28031 27560 28212 27588
rect 28272 27560 30665 27588
rect 28031 27557 28043 27560
rect 27985 27551 28043 27557
rect 27614 27520 27620 27532
rect 24995 27492 26648 27520
rect 26804 27492 27620 27520
rect 24995 27489 25007 27492
rect 24949 27483 25007 27489
rect 25222 27452 25228 27464
rect 24872 27424 25228 27452
rect 23934 27344 23940 27396
rect 23992 27384 23998 27396
rect 24320 27390 24624 27418
rect 24765 27415 24823 27421
rect 24320 27384 24348 27390
rect 23992 27356 24348 27384
rect 24596 27384 24624 27390
rect 24780 27384 24808 27415
rect 25222 27412 25228 27424
rect 25280 27412 25286 27464
rect 25498 27412 25504 27464
rect 25556 27452 25562 27464
rect 25685 27455 25743 27461
rect 25685 27452 25697 27455
rect 25556 27424 25697 27452
rect 25556 27412 25562 27424
rect 25685 27421 25697 27424
rect 25731 27452 25743 27455
rect 25958 27452 25964 27464
rect 25731 27424 25964 27452
rect 25731 27421 25743 27424
rect 25685 27415 25743 27421
rect 25958 27412 25964 27424
rect 26016 27412 26022 27464
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27452 26111 27455
rect 26142 27452 26148 27464
rect 26099 27424 26148 27452
rect 26099 27421 26111 27424
rect 26053 27415 26111 27421
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 26804 27452 26832 27492
rect 27614 27480 27620 27492
rect 27672 27480 27678 27532
rect 28077 27523 28135 27529
rect 26528 27424 26832 27452
rect 26973 27455 27031 27461
rect 26326 27384 26332 27396
rect 24596 27356 26332 27384
rect 23992 27344 23998 27356
rect 26326 27344 26332 27356
rect 26384 27344 26390 27396
rect 23624 27288 23704 27316
rect 23624 27276 23630 27288
rect 24026 27276 24032 27328
rect 24084 27316 24090 27328
rect 24581 27319 24639 27325
rect 24581 27316 24593 27319
rect 24084 27288 24593 27316
rect 24084 27276 24090 27288
rect 24581 27285 24593 27288
rect 24627 27285 24639 27319
rect 24581 27279 24639 27285
rect 24854 27276 24860 27328
rect 24912 27316 24918 27328
rect 25314 27316 25320 27328
rect 24912 27288 25320 27316
rect 24912 27276 24918 27288
rect 25314 27276 25320 27288
rect 25372 27276 25378 27328
rect 25682 27276 25688 27328
rect 25740 27316 25746 27328
rect 26528 27316 26556 27424
rect 26973 27421 26985 27455
rect 27019 27421 27031 27455
rect 26973 27415 27031 27421
rect 26602 27344 26608 27396
rect 26660 27384 26666 27396
rect 26988 27384 27016 27415
rect 27522 27412 27528 27464
rect 27580 27452 27586 27464
rect 27724 27462 27910 27490
rect 28077 27489 28089 27523
rect 28123 27489 28135 27523
rect 28184 27528 28212 27560
rect 30653 27557 30665 27560
rect 30699 27557 30711 27591
rect 30653 27551 30711 27557
rect 28184 27520 28213 27528
rect 28718 27520 28724 27532
rect 28184 27500 28724 27520
rect 28185 27492 28724 27500
rect 28077 27483 28135 27489
rect 27724 27452 27752 27462
rect 27580 27424 27752 27452
rect 27882 27461 27910 27462
rect 27882 27455 27963 27461
rect 27882 27426 27917 27455
rect 27580 27412 27586 27424
rect 27905 27421 27917 27426
rect 27951 27421 27963 27455
rect 27905 27415 27963 27421
rect 27991 27452 28028 27454
rect 28092 27452 28120 27483
rect 28718 27480 28724 27492
rect 28776 27480 28782 27532
rect 28810 27480 28816 27532
rect 28868 27480 28874 27532
rect 28994 27480 29000 27532
rect 29052 27520 29058 27532
rect 29052 27492 29500 27520
rect 29052 27480 29058 27492
rect 27991 27424 28120 27452
rect 26660 27356 27016 27384
rect 26660 27344 26666 27356
rect 27614 27344 27620 27396
rect 27672 27384 27678 27396
rect 27709 27387 27767 27393
rect 27709 27384 27721 27387
rect 27672 27356 27721 27384
rect 27672 27344 27678 27356
rect 27709 27353 27721 27356
rect 27755 27353 27767 27387
rect 27709 27347 27767 27353
rect 27798 27344 27804 27396
rect 27856 27384 27862 27396
rect 27991 27384 28019 27424
rect 28166 27412 28172 27464
rect 28224 27461 28230 27464
rect 28224 27455 28239 27461
rect 28227 27421 28239 27455
rect 28224 27415 28239 27421
rect 28224 27412 28230 27415
rect 28828 27384 28856 27480
rect 29086 27384 29092 27396
rect 27856 27356 28019 27384
rect 28346 27356 28856 27384
rect 29047 27356 29092 27384
rect 27856 27344 27862 27356
rect 25740 27288 26556 27316
rect 26881 27319 26939 27325
rect 25740 27276 25746 27288
rect 26881 27285 26893 27319
rect 26927 27316 26939 27319
rect 26970 27316 26976 27328
rect 26927 27288 26976 27316
rect 26927 27285 26939 27288
rect 26881 27279 26939 27285
rect 26970 27276 26976 27288
rect 27028 27276 27034 27328
rect 27062 27276 27068 27328
rect 27120 27316 27126 27328
rect 28346 27316 28374 27356
rect 29086 27344 29092 27356
rect 29144 27344 29150 27396
rect 28718 27316 28724 27328
rect 27120 27288 28374 27316
rect 28679 27288 28724 27316
rect 27120 27276 27126 27288
rect 28718 27276 28724 27288
rect 28776 27276 28782 27328
rect 28902 27325 28908 27328
rect 28889 27319 28908 27325
rect 28889 27285 28901 27319
rect 28889 27279 28908 27285
rect 28902 27276 28908 27279
rect 28960 27276 28966 27328
rect 29472 27316 29500 27492
rect 29546 27480 29552 27532
rect 29604 27520 29610 27532
rect 30558 27520 30564 27532
rect 29604 27492 30144 27520
rect 30519 27492 30564 27520
rect 29604 27480 29610 27492
rect 29871 27421 29929 27427
rect 29871 27396 29883 27421
rect 29822 27344 29828 27396
rect 29880 27387 29883 27396
rect 29917 27387 29929 27421
rect 30116 27393 30144 27492
rect 30558 27480 30564 27492
rect 30616 27480 30622 27532
rect 30190 27412 30196 27464
rect 30248 27452 30254 27464
rect 30745 27455 30803 27461
rect 30745 27452 30757 27455
rect 30248 27424 30757 27452
rect 30248 27412 30254 27424
rect 30745 27421 30757 27424
rect 30791 27421 30803 27455
rect 30745 27415 30803 27421
rect 30837 27455 30895 27461
rect 30837 27421 30849 27455
rect 30883 27421 30895 27455
rect 30837 27415 30895 27421
rect 29880 27381 29929 27387
rect 30101 27387 30159 27393
rect 29880 27356 29914 27381
rect 29880 27344 29886 27356
rect 30101 27353 30113 27387
rect 30147 27353 30159 27387
rect 30101 27347 30159 27353
rect 30852 27316 30880 27415
rect 29472 27288 30880 27316
rect 1104 27226 31992 27248
rect 1104 27174 8632 27226
rect 8684 27174 8696 27226
rect 8748 27174 8760 27226
rect 8812 27174 8824 27226
rect 8876 27174 8888 27226
rect 8940 27174 16314 27226
rect 16366 27174 16378 27226
rect 16430 27174 16442 27226
rect 16494 27174 16506 27226
rect 16558 27174 16570 27226
rect 16622 27174 23996 27226
rect 24048 27174 24060 27226
rect 24112 27174 24124 27226
rect 24176 27174 24188 27226
rect 24240 27174 24252 27226
rect 24304 27174 31678 27226
rect 31730 27174 31742 27226
rect 31794 27174 31806 27226
rect 31858 27174 31870 27226
rect 31922 27174 31934 27226
rect 31986 27174 31992 27226
rect 1104 27152 31992 27174
rect 8389 27115 8447 27121
rect 8389 27081 8401 27115
rect 8435 27112 8447 27115
rect 8478 27112 8484 27124
rect 8435 27084 8484 27112
rect 8435 27081 8447 27084
rect 8389 27075 8447 27081
rect 8478 27072 8484 27084
rect 8536 27112 8542 27124
rect 9582 27112 9588 27124
rect 8536 27084 9588 27112
rect 8536 27072 8542 27084
rect 9582 27072 9588 27084
rect 9640 27072 9646 27124
rect 10042 27112 10048 27124
rect 10003 27084 10048 27112
rect 10042 27072 10048 27084
rect 10100 27072 10106 27124
rect 11054 27072 11060 27124
rect 11112 27112 11118 27124
rect 11149 27115 11207 27121
rect 11149 27112 11161 27115
rect 11112 27084 11161 27112
rect 11112 27072 11118 27084
rect 11149 27081 11161 27084
rect 11195 27112 11207 27115
rect 13262 27112 13268 27124
rect 11195 27084 13268 27112
rect 11195 27081 11207 27084
rect 11149 27075 11207 27081
rect 13262 27072 13268 27084
rect 13320 27072 13326 27124
rect 15197 27115 15255 27121
rect 15197 27081 15209 27115
rect 15243 27112 15255 27115
rect 15286 27112 15292 27124
rect 15243 27084 15292 27112
rect 15243 27081 15255 27084
rect 15197 27075 15255 27081
rect 15286 27072 15292 27084
rect 15344 27072 15350 27124
rect 15654 27112 15660 27124
rect 15615 27084 15660 27112
rect 15654 27072 15660 27084
rect 15712 27072 15718 27124
rect 17420 27084 19833 27112
rect 6270 27004 6276 27056
rect 6328 27044 6334 27056
rect 6733 27047 6791 27053
rect 6733 27044 6745 27047
rect 6328 27016 6745 27044
rect 6328 27004 6334 27016
rect 6733 27013 6745 27016
rect 6779 27044 6791 27047
rect 10318 27044 10324 27056
rect 6779 27016 10324 27044
rect 6779 27013 6791 27016
rect 6733 27007 6791 27013
rect 10318 27004 10324 27016
rect 10376 27004 10382 27056
rect 11790 27004 11796 27056
rect 11848 27044 11854 27056
rect 12437 27047 12495 27053
rect 12437 27044 12449 27047
rect 11848 27016 12449 27044
rect 11848 27004 11854 27016
rect 12437 27013 12449 27016
rect 12483 27044 12495 27047
rect 16022 27044 16028 27056
rect 12483 27016 16028 27044
rect 12483 27013 12495 27016
rect 12437 27007 12495 27013
rect 16022 27004 16028 27016
rect 16080 27044 16086 27056
rect 16482 27044 16488 27056
rect 16080 27016 16488 27044
rect 16080 27004 16086 27016
rect 16482 27004 16488 27016
rect 16540 27004 16546 27056
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 17126 27044 17132 27056
rect 16816 27016 17132 27044
rect 16816 27004 16822 27016
rect 17126 27004 17132 27016
rect 17184 27004 17190 27056
rect 9122 26936 9128 26988
rect 9180 26976 9186 26988
rect 16209 26979 16267 26985
rect 16209 26976 16221 26979
rect 9180 26948 16221 26976
rect 9180 26936 9186 26948
rect 16209 26945 16221 26948
rect 16255 26945 16267 26979
rect 16209 26939 16267 26945
rect 17034 26936 17040 26988
rect 17092 26976 17098 26988
rect 17221 26979 17279 26985
rect 17221 26976 17233 26979
rect 17092 26948 17233 26976
rect 17092 26936 17098 26948
rect 17221 26945 17233 26948
rect 17267 26945 17279 26979
rect 17221 26939 17279 26945
rect 17310 26936 17316 26988
rect 17368 26936 17374 26988
rect 17420 26985 17448 27084
rect 17957 27047 18015 27053
rect 17957 27013 17969 27047
rect 18003 27044 18015 27047
rect 18230 27044 18236 27056
rect 18003 27016 18236 27044
rect 18003 27013 18015 27016
rect 17957 27007 18015 27013
rect 18230 27004 18236 27016
rect 18288 27044 18294 27056
rect 19805 27044 19833 27084
rect 19886 27072 19892 27124
rect 19944 27112 19950 27124
rect 21085 27115 21143 27121
rect 19944 27084 20668 27112
rect 19944 27072 19950 27084
rect 20162 27044 20168 27056
rect 18288 27016 19773 27044
rect 19805 27016 20168 27044
rect 18288 27004 18294 27016
rect 17405 26979 17463 26985
rect 17405 26945 17417 26979
rect 17451 26945 17463 26979
rect 17405 26939 17463 26945
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 18141 26979 18199 26985
rect 18141 26976 18153 26979
rect 18104 26948 18153 26976
rect 18104 26936 18110 26948
rect 18141 26945 18153 26948
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 18877 26979 18935 26985
rect 18877 26945 18889 26979
rect 18923 26976 18935 26979
rect 19058 26976 19064 26988
rect 18923 26948 19064 26976
rect 18923 26945 18935 26948
rect 18877 26939 18935 26945
rect 19058 26936 19064 26948
rect 19116 26936 19122 26988
rect 19150 26936 19156 26988
rect 19208 26976 19214 26988
rect 19337 26979 19395 26985
rect 19337 26976 19349 26979
rect 19208 26948 19349 26976
rect 19208 26936 19214 26948
rect 19337 26945 19349 26948
rect 19383 26945 19395 26979
rect 19337 26939 19395 26945
rect 19521 26979 19579 26985
rect 19521 26945 19533 26979
rect 19567 26976 19579 26979
rect 19610 26976 19616 26988
rect 19567 26948 19616 26976
rect 19567 26945 19579 26948
rect 19521 26939 19579 26945
rect 19610 26936 19616 26948
rect 19668 26936 19674 26988
rect 19745 26976 19773 27016
rect 20162 27004 20168 27016
rect 20220 27004 20226 27056
rect 20533 27047 20591 27053
rect 20303 27013 20361 27019
rect 20303 26979 20315 27013
rect 20349 26979 20361 27013
rect 20533 27013 20545 27047
rect 20579 27013 20591 27047
rect 20640 27044 20668 27084
rect 21085 27081 21097 27115
rect 21131 27112 21143 27115
rect 21358 27112 21364 27124
rect 21131 27084 21364 27112
rect 21131 27081 21143 27084
rect 21085 27075 21143 27081
rect 21358 27072 21364 27084
rect 21416 27072 21422 27124
rect 21453 27115 21511 27121
rect 21453 27081 21465 27115
rect 21499 27112 21511 27115
rect 22922 27112 22928 27124
rect 21499 27084 22928 27112
rect 21499 27081 21511 27084
rect 21453 27075 21511 27081
rect 22922 27072 22928 27084
rect 22980 27072 22986 27124
rect 23370 27112 23376 27124
rect 23032 27084 23376 27112
rect 23032 27044 23060 27084
rect 23370 27072 23376 27084
rect 23428 27072 23434 27124
rect 23474 27072 23480 27124
rect 23532 27112 23538 27124
rect 24026 27112 24032 27124
rect 23532 27084 24032 27112
rect 23532 27072 23538 27084
rect 24026 27072 24032 27084
rect 24084 27072 24090 27124
rect 24397 27115 24455 27121
rect 24397 27081 24409 27115
rect 24443 27081 24455 27115
rect 24397 27075 24455 27081
rect 20640 27016 22692 27044
rect 20533 27007 20591 27013
rect 20303 26976 20361 26979
rect 19745 26973 20361 26976
rect 19745 26948 20346 26973
rect 7837 26911 7895 26917
rect 7837 26877 7849 26911
rect 7883 26908 7895 26911
rect 9490 26908 9496 26920
rect 7883 26880 9496 26908
rect 7883 26877 7895 26880
rect 7837 26871 7895 26877
rect 9490 26868 9496 26880
rect 9548 26908 9554 26920
rect 14093 26911 14151 26917
rect 14093 26908 14105 26911
rect 9548 26880 14105 26908
rect 9548 26868 9554 26880
rect 14093 26877 14105 26880
rect 14139 26908 14151 26911
rect 14182 26908 14188 26920
rect 14139 26880 14188 26908
rect 14139 26877 14151 26880
rect 14093 26871 14151 26877
rect 14182 26868 14188 26880
rect 14240 26868 14246 26920
rect 17328 26908 17356 26936
rect 17052 26880 17356 26908
rect 17052 26852 17080 26880
rect 17494 26868 17500 26920
rect 17552 26908 17558 26920
rect 18230 26908 18236 26920
rect 17552 26880 18236 26908
rect 17552 26868 17558 26880
rect 18230 26868 18236 26880
rect 18288 26868 18294 26920
rect 18598 26908 18604 26920
rect 18559 26880 18604 26908
rect 18598 26868 18604 26880
rect 18656 26868 18662 26920
rect 18966 26868 18972 26920
rect 19024 26908 19030 26920
rect 20548 26908 20576 27007
rect 20993 26979 21051 26985
rect 20993 26945 21005 26979
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26976 21327 26979
rect 21358 26976 21364 26988
rect 21315 26948 21364 26976
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 19024 26880 20576 26908
rect 19024 26868 19030 26880
rect 8941 26843 8999 26849
rect 8941 26809 8953 26843
rect 8987 26840 8999 26843
rect 11606 26840 11612 26852
rect 8987 26812 11612 26840
rect 8987 26809 8999 26812
rect 8941 26803 8999 26809
rect 11606 26800 11612 26812
rect 11664 26800 11670 26852
rect 11974 26800 11980 26852
rect 12032 26840 12038 26852
rect 15378 26840 15384 26852
rect 12032 26812 15384 26840
rect 12032 26800 12038 26812
rect 15378 26800 15384 26812
rect 15436 26800 15442 26852
rect 16206 26840 16212 26852
rect 15488 26812 16212 26840
rect 7282 26772 7288 26784
rect 7243 26744 7288 26772
rect 7282 26732 7288 26744
rect 7340 26732 7346 26784
rect 9493 26775 9551 26781
rect 9493 26741 9505 26775
rect 9539 26772 9551 26775
rect 9582 26772 9588 26784
rect 9539 26744 9588 26772
rect 9539 26741 9551 26744
rect 9493 26735 9551 26741
rect 9582 26732 9588 26744
rect 9640 26732 9646 26784
rect 10502 26772 10508 26784
rect 10463 26744 10508 26772
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 10870 26732 10876 26784
rect 10928 26772 10934 26784
rect 11793 26775 11851 26781
rect 11793 26772 11805 26775
rect 10928 26744 11805 26772
rect 10928 26732 10934 26744
rect 11793 26741 11805 26744
rect 11839 26741 11851 26775
rect 12986 26772 12992 26784
rect 12947 26744 12992 26772
rect 11793 26735 11851 26741
rect 12986 26732 12992 26744
rect 13044 26732 13050 26784
rect 13446 26772 13452 26784
rect 13407 26744 13452 26772
rect 13446 26732 13452 26744
rect 13504 26732 13510 26784
rect 13630 26732 13636 26784
rect 13688 26772 13694 26784
rect 14553 26775 14611 26781
rect 14553 26772 14565 26775
rect 13688 26744 14565 26772
rect 13688 26732 13694 26744
rect 14553 26741 14565 26744
rect 14599 26772 14611 26775
rect 15102 26772 15108 26784
rect 14599 26744 15108 26772
rect 14599 26741 14611 26744
rect 14553 26735 14611 26741
rect 15102 26732 15108 26744
rect 15160 26732 15166 26784
rect 15286 26732 15292 26784
rect 15344 26772 15350 26784
rect 15488 26772 15516 26812
rect 16206 26800 16212 26812
rect 16264 26800 16270 26852
rect 17034 26800 17040 26852
rect 17092 26800 17098 26852
rect 17310 26800 17316 26852
rect 17368 26840 17374 26852
rect 17368 26812 18078 26840
rect 17368 26800 17374 26812
rect 15344 26744 15516 26772
rect 15344 26732 15350 26744
rect 16574 26732 16580 26784
rect 16632 26772 16638 26784
rect 17126 26772 17132 26784
rect 16632 26744 17132 26772
rect 16632 26732 16638 26744
rect 17126 26732 17132 26744
rect 17184 26732 17190 26784
rect 17405 26775 17463 26781
rect 17405 26741 17417 26775
rect 17451 26772 17463 26775
rect 17954 26772 17960 26784
rect 17451 26744 17960 26772
rect 17451 26741 17463 26744
rect 17405 26735 17463 26741
rect 17954 26732 17960 26744
rect 18012 26732 18018 26784
rect 18050 26772 18078 26812
rect 18322 26800 18328 26852
rect 18380 26840 18386 26852
rect 19705 26843 19763 26849
rect 19705 26840 19717 26843
rect 18380 26812 19717 26840
rect 18380 26800 18386 26812
rect 19705 26809 19717 26812
rect 19751 26809 19763 26843
rect 20165 26843 20223 26849
rect 20165 26840 20177 26843
rect 19705 26803 19763 26809
rect 19805 26812 20177 26840
rect 18693 26775 18751 26781
rect 18693 26772 18705 26775
rect 18050 26744 18705 26772
rect 18693 26741 18705 26744
rect 18739 26741 18751 26775
rect 18693 26735 18751 26741
rect 18779 26732 18785 26784
rect 18837 26772 18843 26784
rect 19426 26772 19432 26784
rect 18837 26744 18882 26772
rect 19387 26744 19432 26772
rect 18837 26732 18843 26744
rect 19426 26732 19432 26744
rect 19484 26732 19490 26784
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 19805 26772 19833 26812
rect 20165 26809 20177 26812
rect 20211 26809 20223 26843
rect 20530 26840 20536 26852
rect 20165 26803 20223 26809
rect 20364 26812 20536 26840
rect 19668 26744 19833 26772
rect 19668 26732 19674 26744
rect 19886 26732 19892 26784
rect 19944 26772 19950 26784
rect 20070 26772 20076 26784
rect 19944 26744 20076 26772
rect 19944 26732 19950 26744
rect 20070 26732 20076 26744
rect 20128 26732 20134 26784
rect 20364 26781 20392 26812
rect 20530 26800 20536 26812
rect 20588 26800 20594 26852
rect 21008 26840 21036 26939
rect 21358 26936 21364 26948
rect 21416 26936 21422 26988
rect 21450 26936 21456 26988
rect 21508 26976 21514 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21508 26948 22017 26976
rect 21508 26936 21514 26948
rect 22005 26945 22017 26948
rect 22051 26976 22063 26979
rect 22186 26976 22192 26988
rect 22051 26948 22192 26976
rect 22051 26945 22063 26948
rect 22005 26939 22063 26945
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 22554 26976 22560 26988
rect 22515 26948 22560 26976
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 22664 26985 22692 27016
rect 22750 27016 23060 27044
rect 22649 26979 22707 26985
rect 22649 26945 22661 26979
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 21542 26868 21548 26920
rect 21600 26908 21606 26920
rect 21600 26880 22232 26908
rect 21600 26868 21606 26880
rect 22094 26840 22100 26852
rect 21008 26812 22100 26840
rect 22094 26800 22100 26812
rect 22152 26800 22158 26852
rect 22204 26840 22232 26880
rect 22278 26868 22284 26920
rect 22336 26908 22342 26920
rect 22750 26908 22778 27016
rect 23658 27004 23664 27056
rect 23716 27044 23722 27056
rect 23934 27044 23940 27056
rect 23716 27016 23940 27044
rect 23716 27004 23722 27016
rect 23934 27004 23940 27016
rect 23992 27004 23998 27056
rect 24412 27044 24440 27075
rect 26142 27072 26148 27124
rect 26200 27112 26206 27124
rect 27341 27115 27399 27121
rect 26200 27084 27200 27112
rect 26200 27072 26206 27084
rect 27172 27053 27200 27084
rect 27341 27081 27353 27115
rect 27387 27112 27399 27115
rect 27890 27112 27896 27124
rect 27387 27084 27896 27112
rect 27387 27081 27399 27084
rect 27341 27075 27399 27081
rect 27890 27072 27896 27084
rect 27948 27072 27954 27124
rect 27982 27072 27988 27124
rect 28040 27112 28046 27124
rect 28169 27115 28227 27121
rect 28169 27112 28181 27115
rect 28040 27084 28181 27112
rect 28040 27072 28046 27084
rect 28169 27081 28181 27084
rect 28215 27081 28227 27115
rect 28350 27112 28356 27124
rect 28311 27084 28356 27112
rect 28169 27075 28227 27081
rect 28350 27072 28356 27084
rect 28408 27072 28414 27124
rect 28460 27084 29776 27112
rect 27157 27047 27215 27053
rect 24412 27016 26004 27044
rect 22833 26979 22891 26985
rect 22833 26945 22845 26979
rect 22879 26945 22891 26979
rect 22833 26939 22891 26945
rect 22336 26880 22778 26908
rect 22848 26908 22876 26939
rect 22922 26936 22928 26988
rect 22980 26976 22986 26988
rect 22980 26948 23025 26976
rect 22980 26936 22986 26948
rect 23198 26936 23204 26988
rect 23256 26976 23262 26988
rect 23474 26976 23480 26988
rect 23256 26948 23480 26976
rect 23256 26936 23262 26948
rect 23474 26936 23480 26948
rect 23532 26936 23538 26988
rect 24210 26976 24216 26988
rect 24171 26948 24216 26976
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 24394 26936 24400 26988
rect 24452 26976 24458 26988
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 24452 26948 25053 26976
rect 24452 26936 24458 26948
rect 25041 26945 25053 26948
rect 25087 26976 25099 26979
rect 25087 26948 25268 26976
rect 25087 26945 25099 26948
rect 25041 26939 25099 26945
rect 23290 26908 23296 26920
rect 22848 26880 23296 26908
rect 22336 26868 22342 26880
rect 23290 26868 23296 26880
rect 23348 26868 23354 26920
rect 23382 26868 23388 26920
rect 23440 26908 23446 26920
rect 23753 26911 23811 26917
rect 23753 26908 23765 26911
rect 23440 26880 23765 26908
rect 23440 26868 23446 26880
rect 23753 26877 23765 26880
rect 23799 26877 23811 26911
rect 23753 26871 23811 26877
rect 23842 26868 23848 26920
rect 23900 26908 23906 26920
rect 24118 26908 24124 26920
rect 23900 26880 23945 26908
rect 24079 26880 24124 26908
rect 23900 26868 23906 26880
rect 24118 26868 24124 26880
rect 24176 26868 24182 26920
rect 24302 26868 24308 26920
rect 24360 26908 24366 26920
rect 25240 26908 25268 26948
rect 25314 26936 25320 26988
rect 25372 26985 25378 26988
rect 25372 26979 25408 26985
rect 25396 26945 25408 26979
rect 25372 26939 25408 26945
rect 25372 26936 25378 26939
rect 25498 26936 25504 26988
rect 25556 26976 25562 26988
rect 25976 26976 26004 27016
rect 26064 27016 27005 27044
rect 26064 26976 26092 27016
rect 25556 26948 25601 26976
rect 25976 26948 26092 26976
rect 26191 26979 26249 26985
rect 25556 26936 25562 26948
rect 26191 26945 26203 26979
rect 26237 26945 26249 26979
rect 26326 26976 26332 26988
rect 26287 26948 26332 26976
rect 26191 26939 26249 26945
rect 26206 26908 26234 26939
rect 26326 26936 26332 26948
rect 26384 26936 26390 26988
rect 26418 26936 26424 26988
rect 26476 26976 26482 26988
rect 26605 26979 26663 26985
rect 26476 26948 26521 26976
rect 26476 26936 26482 26948
rect 26605 26945 26617 26979
rect 26651 26976 26663 26979
rect 26878 26976 26884 26988
rect 26651 26948 26884 26976
rect 26651 26945 26663 26948
rect 26605 26939 26663 26945
rect 26878 26936 26884 26948
rect 26936 26936 26942 26988
rect 26786 26908 26792 26920
rect 24360 26880 25176 26908
rect 25240 26880 26096 26908
rect 26206 26880 26792 26908
rect 24360 26868 24366 26880
rect 23014 26840 23020 26852
rect 22204 26812 23020 26840
rect 23014 26800 23020 26812
rect 23072 26800 23078 26852
rect 23198 26800 23204 26852
rect 23256 26840 23262 26852
rect 23256 26812 23520 26840
rect 23256 26800 23262 26812
rect 20349 26775 20407 26781
rect 20349 26741 20361 26775
rect 20395 26741 20407 26775
rect 20349 26735 20407 26741
rect 20438 26732 20444 26784
rect 20496 26772 20502 26784
rect 22554 26772 22560 26784
rect 20496 26744 22560 26772
rect 20496 26732 20502 26744
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 23109 26775 23167 26781
rect 23109 26741 23121 26775
rect 23155 26772 23167 26775
rect 23382 26772 23388 26784
rect 23155 26744 23388 26772
rect 23155 26741 23167 26744
rect 23109 26735 23167 26741
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 23492 26772 23520 26812
rect 23566 26800 23572 26852
rect 23624 26840 23630 26852
rect 24394 26840 24400 26852
rect 23624 26812 24400 26840
rect 23624 26800 23630 26812
rect 24394 26800 24400 26812
rect 24452 26800 24458 26852
rect 25148 26840 25176 26880
rect 25866 26840 25872 26852
rect 25148 26812 25268 26840
rect 24857 26775 24915 26781
rect 24857 26772 24869 26775
rect 23492 26744 24869 26772
rect 24857 26741 24869 26744
rect 24903 26741 24915 26775
rect 25240 26772 25268 26812
rect 25424 26812 25872 26840
rect 25424 26772 25452 26812
rect 25866 26800 25872 26812
rect 25924 26800 25930 26852
rect 26068 26840 26096 26880
rect 26786 26868 26792 26880
rect 26844 26868 26850 26920
rect 26977 26908 27005 27016
rect 27157 27013 27169 27047
rect 27203 27044 27215 27047
rect 28460 27044 28488 27084
rect 27203 27016 28488 27044
rect 27203 27013 27215 27016
rect 27157 27007 27215 27013
rect 28810 27004 28816 27056
rect 28868 27044 28874 27056
rect 29181 27047 29239 27053
rect 29181 27044 29193 27047
rect 28868 27016 29193 27044
rect 28868 27004 28874 27016
rect 29181 27013 29193 27016
rect 29227 27013 29239 27047
rect 29181 27007 29239 27013
rect 29270 27004 29276 27056
rect 29328 27044 29334 27056
rect 29641 27047 29699 27053
rect 29641 27044 29653 27047
rect 29328 27016 29653 27044
rect 29328 27004 29334 27016
rect 29641 27013 29653 27016
rect 29687 27013 29699 27047
rect 29641 27007 29699 27013
rect 27246 26936 27252 26988
rect 27304 26976 27310 26988
rect 27433 26979 27491 26985
rect 27433 26976 27445 26979
rect 27304 26948 27445 26976
rect 27304 26936 27310 26948
rect 27433 26945 27445 26948
rect 27479 26945 27491 26979
rect 27433 26939 27491 26945
rect 27522 26936 27528 26988
rect 27580 26976 27586 26988
rect 27580 26948 27625 26976
rect 27580 26936 27586 26948
rect 27706 26936 27712 26988
rect 27764 26976 27770 26988
rect 27764 26948 27809 26976
rect 27764 26936 27770 26948
rect 27890 26936 27896 26988
rect 27948 26976 27954 26988
rect 28534 26976 28540 26988
rect 27948 26948 28540 26976
rect 27948 26936 27954 26948
rect 28534 26936 28540 26948
rect 28592 26936 28598 26988
rect 28902 26936 28908 26988
rect 28960 26976 28966 26988
rect 29362 26976 29368 26988
rect 28960 26948 29368 26976
rect 28960 26936 28966 26948
rect 29362 26936 29368 26948
rect 29420 26936 29426 26988
rect 29546 26976 29552 26988
rect 29507 26948 29552 26976
rect 29546 26936 29552 26948
rect 29604 26936 29610 26988
rect 28721 26911 28779 26917
rect 28721 26908 28733 26911
rect 26977 26880 28733 26908
rect 28721 26877 28733 26880
rect 28767 26877 28779 26911
rect 28721 26871 28779 26877
rect 29273 26911 29331 26917
rect 29273 26877 29285 26911
rect 29319 26908 29331 26911
rect 29748 26908 29776 27084
rect 29822 27072 29828 27124
rect 29880 27112 29886 27124
rect 30190 27112 30196 27124
rect 29880 27084 30196 27112
rect 29880 27072 29886 27084
rect 30190 27072 30196 27084
rect 30248 27072 30254 27124
rect 30466 27112 30472 27124
rect 30427 27084 30472 27112
rect 30466 27072 30472 27084
rect 30524 27072 30530 27124
rect 31297 27115 31355 27121
rect 31297 27081 31309 27115
rect 31343 27112 31355 27115
rect 31478 27112 31484 27124
rect 31343 27084 31484 27112
rect 31343 27081 31355 27084
rect 31297 27075 31355 27081
rect 31478 27072 31484 27084
rect 31536 27072 31542 27124
rect 30098 27044 30104 27056
rect 30059 27016 30104 27044
rect 30098 27004 30104 27016
rect 30156 27004 30162 27056
rect 30929 27047 30987 27053
rect 30929 27013 30941 27047
rect 30975 27044 30987 27047
rect 31018 27044 31024 27056
rect 30975 27016 31024 27044
rect 30975 27013 30987 27016
rect 30929 27007 30987 27013
rect 31018 27004 31024 27016
rect 31076 27044 31082 27056
rect 31662 27044 31668 27056
rect 31076 27016 31668 27044
rect 31076 27004 31082 27016
rect 31662 27004 31668 27016
rect 31720 27004 31726 27056
rect 30190 26936 30196 26988
rect 30248 26976 30254 26988
rect 30285 26979 30343 26985
rect 30285 26976 30297 26979
rect 30248 26948 30297 26976
rect 30248 26936 30254 26948
rect 30285 26945 30297 26948
rect 30331 26945 30343 26979
rect 30285 26939 30343 26945
rect 31113 26979 31171 26985
rect 31113 26945 31125 26979
rect 31159 26976 31171 26979
rect 31202 26976 31208 26988
rect 31159 26948 31208 26976
rect 31159 26945 31171 26948
rect 31113 26939 31171 26945
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 31754 26908 31760 26920
rect 29319 26880 29500 26908
rect 29748 26880 31760 26908
rect 29319 26877 29331 26880
rect 29273 26871 29331 26877
rect 29362 26840 29368 26852
rect 26068 26812 29368 26840
rect 29362 26800 29368 26812
rect 29420 26800 29426 26852
rect 29472 26840 29500 26880
rect 31754 26868 31760 26880
rect 31812 26868 31818 26920
rect 30926 26840 30932 26852
rect 29472 26812 30932 26840
rect 30926 26800 30932 26812
rect 30984 26800 30990 26852
rect 25240 26744 25452 26772
rect 24857 26735 24915 26741
rect 25590 26732 25596 26784
rect 25648 26772 25654 26784
rect 25961 26775 26019 26781
rect 25961 26772 25973 26775
rect 25648 26744 25973 26772
rect 25648 26732 25654 26744
rect 25961 26741 25973 26744
rect 26007 26741 26019 26775
rect 25961 26735 26019 26741
rect 26234 26732 26240 26784
rect 26292 26772 26298 26784
rect 26786 26772 26792 26784
rect 26292 26744 26792 26772
rect 26292 26732 26298 26744
rect 26786 26732 26792 26744
rect 26844 26732 26850 26784
rect 26878 26732 26884 26784
rect 26936 26772 26942 26784
rect 27062 26772 27068 26784
rect 26936 26744 27068 26772
rect 26936 26732 26942 26744
rect 27062 26732 27068 26744
rect 27120 26732 27126 26784
rect 27522 26732 27528 26784
rect 27580 26772 27586 26784
rect 27890 26772 27896 26784
rect 27580 26744 27896 26772
rect 27580 26732 27586 26744
rect 27890 26732 27896 26744
rect 27948 26732 27954 26784
rect 28074 26732 28080 26784
rect 28132 26772 28138 26784
rect 28167 26772 28173 26784
rect 28132 26744 28173 26772
rect 28132 26732 28138 26744
rect 28167 26732 28173 26744
rect 28225 26732 28231 26784
rect 28331 26775 28389 26781
rect 28331 26741 28343 26775
rect 28377 26772 28389 26775
rect 28718 26772 28724 26784
rect 28377 26744 28724 26772
rect 28377 26741 28389 26744
rect 28331 26735 28389 26741
rect 28718 26732 28724 26744
rect 28776 26732 28782 26784
rect 29270 26732 29276 26784
rect 29328 26772 29334 26784
rect 29822 26772 29828 26784
rect 29328 26744 29828 26772
rect 29328 26732 29334 26744
rect 29822 26732 29828 26744
rect 29880 26732 29886 26784
rect 1104 26682 31832 26704
rect 1104 26630 4791 26682
rect 4843 26630 4855 26682
rect 4907 26630 4919 26682
rect 4971 26630 4983 26682
rect 5035 26630 5047 26682
rect 5099 26630 12473 26682
rect 12525 26630 12537 26682
rect 12589 26630 12601 26682
rect 12653 26630 12665 26682
rect 12717 26630 12729 26682
rect 12781 26630 20155 26682
rect 20207 26630 20219 26682
rect 20271 26630 20283 26682
rect 20335 26630 20347 26682
rect 20399 26630 20411 26682
rect 20463 26630 27837 26682
rect 27889 26630 27901 26682
rect 27953 26630 27965 26682
rect 28017 26630 28029 26682
rect 28081 26630 28093 26682
rect 28145 26630 31832 26682
rect 1104 26608 31832 26630
rect 8573 26571 8631 26577
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 10962 26568 10968 26580
rect 8619 26540 10968 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 10962 26528 10968 26540
rect 11020 26528 11026 26580
rect 11517 26571 11575 26577
rect 11517 26537 11529 26571
rect 11563 26568 11575 26571
rect 12250 26568 12256 26580
rect 11563 26540 12256 26568
rect 11563 26537 11575 26540
rect 11517 26531 11575 26537
rect 12250 26528 12256 26540
rect 12308 26528 12314 26580
rect 12342 26528 12348 26580
rect 12400 26568 12406 26580
rect 12529 26571 12587 26577
rect 12529 26568 12541 26571
rect 12400 26540 12541 26568
rect 12400 26528 12406 26540
rect 12529 26537 12541 26540
rect 12575 26537 12587 26571
rect 13078 26568 13084 26580
rect 12529 26531 12587 26537
rect 12636 26540 13084 26568
rect 10594 26460 10600 26512
rect 10652 26500 10658 26512
rect 10873 26503 10931 26509
rect 10873 26500 10885 26503
rect 10652 26472 10885 26500
rect 10652 26460 10658 26472
rect 10873 26469 10885 26472
rect 10919 26469 10931 26503
rect 10873 26463 10931 26469
rect 11606 26460 11612 26512
rect 11664 26500 11670 26512
rect 12636 26500 12664 26540
rect 13078 26528 13084 26540
rect 13136 26528 13142 26580
rect 13262 26528 13268 26580
rect 13320 26568 13326 26580
rect 13630 26568 13636 26580
rect 13320 26540 13636 26568
rect 13320 26528 13326 26540
rect 13630 26528 13636 26540
rect 13688 26528 13694 26580
rect 14642 26568 14648 26580
rect 14603 26540 14648 26568
rect 14642 26528 14648 26540
rect 14700 26528 14706 26580
rect 16206 26568 16212 26580
rect 15228 26540 16212 26568
rect 11664 26472 12664 26500
rect 11664 26460 11670 26472
rect 5166 26392 5172 26444
rect 5224 26432 5230 26444
rect 5813 26435 5871 26441
rect 5813 26432 5825 26435
rect 5224 26404 5825 26432
rect 5224 26392 5230 26404
rect 5813 26401 5825 26404
rect 5859 26432 5871 26435
rect 10413 26435 10471 26441
rect 10413 26432 10425 26435
rect 5859 26404 10425 26432
rect 5859 26401 5871 26404
rect 5813 26395 5871 26401
rect 10413 26401 10425 26404
rect 10459 26432 10471 26435
rect 11790 26432 11796 26444
rect 10459 26404 11796 26432
rect 10459 26401 10471 26404
rect 10413 26395 10471 26401
rect 11790 26392 11796 26404
rect 11848 26392 11854 26444
rect 12250 26392 12256 26444
rect 12308 26432 12314 26444
rect 15228 26432 15256 26540
rect 16206 26528 16212 26540
rect 16264 26568 16270 26580
rect 16850 26568 16856 26580
rect 16264 26540 16856 26568
rect 16264 26528 16270 26540
rect 16850 26528 16856 26540
rect 16908 26528 16914 26580
rect 17034 26528 17040 26580
rect 17092 26568 17098 26580
rect 17129 26571 17187 26577
rect 17129 26568 17141 26571
rect 17092 26540 17141 26568
rect 17092 26528 17098 26540
rect 17129 26537 17141 26540
rect 17175 26537 17187 26571
rect 17129 26531 17187 26537
rect 17221 26571 17279 26577
rect 17221 26537 17233 26571
rect 17267 26568 17279 26571
rect 17586 26568 17592 26580
rect 17267 26540 17592 26568
rect 17267 26537 17279 26540
rect 17221 26531 17279 26537
rect 17586 26528 17592 26540
rect 17644 26528 17650 26580
rect 17862 26528 17868 26580
rect 17920 26568 17926 26580
rect 18877 26571 18935 26577
rect 18877 26568 18889 26571
rect 17920 26540 18889 26568
rect 17920 26528 17926 26540
rect 18877 26537 18889 26540
rect 18923 26537 18935 26571
rect 18877 26531 18935 26537
rect 19981 26571 20039 26577
rect 19981 26537 19993 26571
rect 20027 26568 20039 26571
rect 20530 26568 20536 26580
rect 20027 26540 20536 26568
rect 20027 26537 20039 26540
rect 19981 26531 20039 26537
rect 20530 26528 20536 26540
rect 20588 26528 20594 26580
rect 20901 26571 20959 26577
rect 20901 26537 20913 26571
rect 20947 26537 20959 26571
rect 22002 26568 22008 26580
rect 20901 26531 20959 26537
rect 21008 26540 22008 26568
rect 15286 26460 15292 26512
rect 15344 26500 15350 26512
rect 16574 26500 16580 26512
rect 15344 26472 16580 26500
rect 15344 26460 15350 26472
rect 16574 26460 16580 26472
rect 16632 26460 16638 26512
rect 16960 26472 18078 26500
rect 12308 26404 15256 26432
rect 15841 26435 15899 26441
rect 12308 26392 12314 26404
rect 15841 26401 15853 26435
rect 15887 26432 15899 26435
rect 15887 26404 16804 26432
rect 15887 26401 15899 26404
rect 15841 26395 15899 26401
rect 1578 26364 1584 26376
rect 1539 26336 1584 26364
rect 1578 26324 1584 26336
rect 1636 26324 1642 26376
rect 9306 26364 9312 26376
rect 9267 26336 9312 26364
rect 9306 26324 9312 26336
rect 9364 26324 9370 26376
rect 9398 26324 9404 26376
rect 9456 26364 9462 26376
rect 12894 26364 12900 26376
rect 9456 26336 12900 26364
rect 9456 26324 9462 26336
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26333 15807 26367
rect 15930 26364 15936 26376
rect 15891 26336 15936 26364
rect 15749 26327 15807 26333
rect 6365 26299 6423 26305
rect 6365 26265 6377 26299
rect 6411 26296 6423 26299
rect 6822 26296 6828 26308
rect 6411 26268 6828 26296
rect 6411 26265 6423 26268
rect 6365 26259 6423 26265
rect 6822 26256 6828 26268
rect 6880 26256 6886 26308
rect 6917 26299 6975 26305
rect 6917 26265 6929 26299
rect 6963 26296 6975 26299
rect 7926 26296 7932 26308
rect 6963 26268 7788 26296
rect 7887 26268 7932 26296
rect 6963 26265 6975 26268
rect 6917 26259 6975 26265
rect 7466 26228 7472 26240
rect 7427 26200 7472 26228
rect 7466 26188 7472 26200
rect 7524 26188 7530 26240
rect 7760 26228 7788 26268
rect 7926 26256 7932 26268
rect 7984 26256 7990 26308
rect 9766 26296 9772 26308
rect 9727 26268 9772 26296
rect 9766 26256 9772 26268
rect 9824 26256 9830 26308
rect 12066 26296 12072 26308
rect 12027 26268 12072 26296
rect 12066 26256 12072 26268
rect 12124 26256 12130 26308
rect 14458 26256 14464 26308
rect 14516 26296 14522 26308
rect 15102 26296 15108 26308
rect 14516 26268 15108 26296
rect 14516 26256 14522 26268
rect 15102 26256 15108 26268
rect 15160 26296 15166 26308
rect 15197 26299 15255 26305
rect 15197 26296 15209 26299
rect 15160 26268 15209 26296
rect 15160 26256 15166 26268
rect 15197 26265 15209 26268
rect 15243 26265 15255 26299
rect 15197 26259 15255 26265
rect 15654 26256 15660 26308
rect 15712 26296 15718 26308
rect 15764 26296 15792 26327
rect 15930 26324 15936 26336
rect 15988 26324 15994 26376
rect 16390 26364 16396 26376
rect 16351 26336 16396 26364
rect 16390 26324 16396 26336
rect 16448 26324 16454 26376
rect 16574 26364 16580 26376
rect 16535 26336 16580 26364
rect 16574 26324 16580 26336
rect 16632 26324 16638 26376
rect 16666 26324 16672 26376
rect 16724 26364 16730 26376
rect 16776 26364 16804 26404
rect 16960 26364 16988 26472
rect 17313 26435 17371 26441
rect 17313 26401 17325 26435
rect 17359 26432 17371 26435
rect 17402 26432 17408 26444
rect 17359 26404 17408 26432
rect 17359 26401 17371 26404
rect 17313 26395 17371 26401
rect 17402 26392 17408 26404
rect 17460 26392 17466 26444
rect 17586 26392 17592 26444
rect 17644 26432 17650 26444
rect 17773 26435 17831 26441
rect 17773 26432 17785 26435
rect 17644 26404 17785 26432
rect 17644 26392 17650 26404
rect 17773 26401 17785 26404
rect 17819 26401 17831 26435
rect 17773 26395 17831 26401
rect 17862 26392 17868 26444
rect 17920 26432 17926 26444
rect 17957 26435 18015 26441
rect 17957 26432 17969 26435
rect 17920 26404 17969 26432
rect 17920 26392 17926 26404
rect 17957 26401 17969 26404
rect 18003 26401 18015 26435
rect 18050 26432 18078 26472
rect 18230 26460 18236 26512
rect 18288 26500 18294 26512
rect 19610 26500 19616 26512
rect 18288 26472 19616 26500
rect 18288 26460 18294 26472
rect 19610 26460 19616 26472
rect 19668 26460 19674 26512
rect 19797 26503 19855 26509
rect 19797 26469 19809 26503
rect 19843 26500 19855 26503
rect 19843 26472 20300 26500
rect 19843 26469 19855 26472
rect 19797 26463 19855 26469
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 18050 26404 19901 26432
rect 17957 26395 18015 26401
rect 19889 26401 19901 26404
rect 19935 26401 19947 26435
rect 19889 26395 19947 26401
rect 16724 26336 16804 26364
rect 16856 26336 16988 26364
rect 16724 26324 16730 26336
rect 15838 26296 15844 26308
rect 15712 26268 15844 26296
rect 15712 26256 15718 26268
rect 15838 26256 15844 26268
rect 15896 26256 15902 26308
rect 16482 26256 16488 26308
rect 16540 26296 16546 26308
rect 16856 26296 16884 26336
rect 17034 26324 17040 26376
rect 17092 26364 17098 26376
rect 18049 26367 18107 26373
rect 17092 26336 17137 26364
rect 17092 26324 17098 26336
rect 18049 26333 18061 26367
rect 18095 26364 18107 26367
rect 18230 26364 18236 26376
rect 18095 26336 18236 26364
rect 18095 26333 18107 26336
rect 18049 26327 18107 26333
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18601 26367 18659 26373
rect 18601 26364 18613 26367
rect 18472 26336 18613 26364
rect 18472 26324 18478 26336
rect 18601 26333 18613 26336
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 18690 26324 18696 26376
rect 18748 26364 18754 26376
rect 19150 26364 19156 26376
rect 18748 26336 19156 26364
rect 18748 26324 18754 26336
rect 19150 26324 19156 26336
rect 19208 26324 19214 26376
rect 19702 26324 19708 26376
rect 19760 26364 19766 26376
rect 19978 26364 19984 26376
rect 19760 26336 19984 26364
rect 19760 26324 19766 26336
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 20070 26324 20076 26376
rect 20128 26364 20134 26376
rect 20272 26364 20300 26472
rect 20622 26460 20628 26512
rect 20680 26500 20686 26512
rect 20717 26503 20775 26509
rect 20717 26500 20729 26503
rect 20680 26472 20729 26500
rect 20680 26460 20686 26472
rect 20717 26469 20729 26472
rect 20763 26469 20775 26503
rect 20717 26463 20775 26469
rect 20346 26392 20352 26444
rect 20404 26432 20410 26444
rect 20916 26432 20944 26531
rect 21008 26441 21036 26540
rect 22002 26528 22008 26540
rect 22060 26528 22066 26580
rect 25038 26568 25044 26580
rect 23032 26540 25044 26568
rect 21174 26460 21180 26512
rect 21232 26500 21238 26512
rect 23032 26500 23060 26540
rect 25038 26528 25044 26540
rect 25096 26568 25102 26580
rect 25590 26568 25596 26580
rect 25096 26540 25596 26568
rect 25096 26528 25102 26540
rect 25590 26528 25596 26540
rect 25648 26568 25654 26580
rect 28902 26568 28908 26580
rect 25648 26540 27936 26568
rect 25648 26528 25654 26540
rect 21232 26472 21864 26500
rect 21232 26460 21238 26472
rect 21836 26441 21864 26472
rect 21928 26472 23060 26500
rect 20404 26404 20944 26432
rect 20993 26435 21051 26441
rect 20404 26392 20410 26404
rect 20993 26401 21005 26435
rect 21039 26401 21051 26435
rect 20993 26395 21051 26401
rect 21821 26435 21879 26441
rect 21821 26401 21833 26435
rect 21867 26401 21879 26435
rect 21821 26395 21879 26401
rect 21174 26364 21180 26376
rect 20128 26336 20173 26364
rect 20272 26358 20392 26364
rect 20548 26358 21180 26364
rect 20272 26336 21180 26358
rect 20128 26324 20134 26336
rect 20364 26330 20576 26336
rect 21174 26324 21180 26336
rect 21232 26324 21238 26376
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26364 21327 26367
rect 21928 26364 21956 26472
rect 23106 26460 23112 26512
rect 23164 26460 23170 26512
rect 23474 26500 23480 26512
rect 23296 26472 23480 26500
rect 22186 26392 22192 26444
rect 22244 26392 22250 26444
rect 22554 26392 22560 26444
rect 22612 26392 22618 26444
rect 23124 26432 23152 26460
rect 23124 26404 23244 26432
rect 21315 26336 21956 26364
rect 21991 26367 22049 26373
rect 21315 26333 21327 26336
rect 21269 26327 21327 26333
rect 21991 26333 22003 26367
rect 22037 26364 22049 26367
rect 22204 26364 22232 26392
rect 22037 26336 22232 26364
rect 22572 26364 22600 26392
rect 23216 26373 23244 26404
rect 23109 26367 23167 26373
rect 23109 26364 23121 26367
rect 22572 26336 23121 26364
rect 22037 26333 22049 26336
rect 21991 26327 22049 26333
rect 23109 26333 23121 26336
rect 23155 26333 23167 26367
rect 23109 26327 23167 26333
rect 23201 26367 23259 26373
rect 23201 26333 23213 26367
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 16540 26268 16884 26296
rect 16540 26256 16546 26268
rect 17402 26256 17408 26308
rect 17460 26296 17466 26308
rect 19886 26296 19892 26308
rect 17460 26268 19892 26296
rect 17460 26256 17466 26268
rect 19886 26256 19892 26268
rect 19944 26256 19950 26308
rect 20257 26299 20315 26305
rect 20257 26265 20269 26299
rect 20303 26296 20315 26299
rect 22554 26296 22560 26308
rect 20303 26268 22560 26296
rect 20303 26265 20315 26268
rect 20257 26259 20315 26265
rect 22554 26256 22560 26268
rect 22612 26256 22618 26308
rect 23296 26296 23324 26472
rect 23474 26460 23480 26472
rect 23532 26500 23538 26512
rect 23532 26472 25452 26500
rect 23532 26460 23538 26472
rect 23382 26392 23388 26444
rect 23440 26392 23446 26444
rect 25317 26435 25375 26441
rect 25317 26432 25329 26435
rect 23676 26404 25329 26432
rect 23400 26305 23428 26392
rect 23566 26364 23572 26376
rect 23527 26336 23572 26364
rect 23566 26324 23572 26336
rect 23624 26324 23630 26376
rect 22664 26268 23324 26296
rect 23385 26299 23443 26305
rect 12342 26228 12348 26240
rect 7760 26200 12348 26228
rect 12342 26188 12348 26200
rect 12400 26188 12406 26240
rect 12710 26188 12716 26240
rect 12768 26228 12774 26240
rect 13630 26228 13636 26240
rect 12768 26200 13636 26228
rect 12768 26188 12774 26200
rect 13630 26188 13636 26200
rect 13688 26188 13694 26240
rect 16577 26231 16635 26237
rect 16577 26197 16589 26231
rect 16623 26228 16635 26231
rect 17034 26228 17040 26240
rect 16623 26200 17040 26228
rect 16623 26197 16635 26200
rect 16577 26191 16635 26197
rect 17034 26188 17040 26200
rect 17092 26188 17098 26240
rect 17126 26188 17132 26240
rect 17184 26228 17190 26240
rect 17773 26231 17831 26237
rect 17773 26228 17785 26231
rect 17184 26200 17785 26228
rect 17184 26188 17190 26200
rect 17773 26197 17785 26200
rect 17819 26197 17831 26231
rect 17773 26191 17831 26197
rect 18138 26188 18144 26240
rect 18196 26228 18202 26240
rect 18598 26228 18604 26240
rect 18196 26200 18604 26228
rect 18196 26188 18202 26200
rect 18598 26188 18604 26200
rect 18656 26188 18662 26240
rect 19058 26188 19064 26240
rect 19116 26228 19122 26240
rect 21358 26228 21364 26240
rect 19116 26200 21364 26228
rect 19116 26188 19122 26200
rect 21358 26188 21364 26200
rect 21416 26188 21422 26240
rect 21910 26188 21916 26240
rect 21968 26228 21974 26240
rect 22281 26231 22339 26237
rect 22281 26228 22293 26231
rect 21968 26200 22293 26228
rect 21968 26188 21974 26200
rect 22281 26197 22293 26200
rect 22327 26197 22339 26231
rect 22281 26191 22339 26197
rect 22370 26188 22376 26240
rect 22428 26228 22434 26240
rect 22664 26228 22692 26268
rect 23385 26265 23397 26299
rect 23431 26265 23443 26299
rect 23385 26259 23443 26265
rect 23474 26256 23480 26308
rect 23532 26296 23538 26308
rect 23532 26268 23577 26296
rect 23532 26256 23538 26268
rect 22428 26200 22692 26228
rect 22428 26188 22434 26200
rect 22738 26188 22744 26240
rect 22796 26228 22802 26240
rect 23676 26228 23704 26404
rect 25317 26401 25329 26404
rect 25363 26401 25375 26435
rect 25424 26432 25452 26472
rect 25682 26460 25688 26512
rect 25740 26500 25746 26512
rect 25777 26503 25835 26509
rect 25777 26500 25789 26503
rect 25740 26472 25789 26500
rect 25740 26460 25746 26472
rect 25777 26469 25789 26472
rect 25823 26469 25835 26503
rect 25777 26463 25835 26469
rect 26418 26460 26424 26512
rect 26476 26460 26482 26512
rect 26694 26460 26700 26512
rect 26752 26500 26758 26512
rect 26752 26472 27325 26500
rect 26752 26460 26758 26472
rect 25866 26432 25872 26444
rect 25424 26404 25872 26432
rect 25317 26395 25375 26401
rect 25866 26392 25872 26404
rect 25924 26432 25930 26444
rect 26053 26435 26111 26441
rect 26053 26432 26065 26435
rect 25924 26404 26065 26432
rect 25924 26392 25930 26404
rect 26053 26401 26065 26404
rect 26099 26401 26111 26435
rect 26436 26432 26464 26460
rect 26436 26404 27108 26432
rect 26053 26395 26111 26401
rect 27080 26376 27108 26404
rect 23842 26324 23848 26376
rect 23900 26324 23906 26376
rect 23934 26324 23940 26376
rect 23992 26364 23998 26376
rect 24857 26367 24915 26373
rect 24857 26364 24869 26367
rect 23992 26336 24869 26364
rect 23992 26324 23998 26336
rect 24857 26333 24869 26336
rect 24903 26333 24915 26367
rect 24857 26327 24915 26333
rect 25041 26367 25099 26373
rect 25041 26333 25053 26367
rect 25087 26364 25099 26367
rect 25130 26364 25136 26376
rect 25087 26336 25136 26364
rect 25087 26333 25099 26336
rect 25041 26327 25099 26333
rect 25130 26324 25136 26336
rect 25188 26324 25194 26376
rect 25225 26367 25283 26373
rect 25225 26333 25237 26367
rect 25271 26364 25283 26367
rect 25271 26361 25452 26364
rect 25271 26336 25636 26361
rect 25271 26333 25283 26336
rect 25424 26333 25636 26336
rect 25225 26327 25283 26333
rect 22796 26200 23704 26228
rect 23753 26231 23811 26237
rect 22796 26188 22802 26200
rect 23753 26197 23765 26231
rect 23799 26228 23811 26231
rect 23860 26228 23888 26324
rect 24578 26296 24584 26308
rect 24539 26268 24584 26296
rect 24578 26256 24584 26268
rect 24636 26256 24642 26308
rect 23799 26200 23888 26228
rect 23799 26197 23811 26200
rect 23753 26191 23811 26197
rect 24670 26188 24676 26240
rect 24728 26228 24734 26240
rect 24949 26231 25007 26237
rect 24949 26228 24961 26231
rect 24728 26200 24961 26228
rect 24728 26188 24734 26200
rect 24949 26197 24961 26200
rect 24995 26197 25007 26231
rect 25608 26228 25636 26333
rect 25682 26324 25688 26376
rect 25740 26364 25746 26376
rect 25961 26367 26019 26373
rect 25961 26364 25973 26367
rect 25740 26336 25973 26364
rect 25740 26324 25746 26336
rect 25961 26333 25973 26336
rect 26007 26333 26019 26367
rect 26142 26364 26148 26376
rect 26103 26336 26148 26364
rect 25961 26327 26019 26333
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 26237 26367 26295 26373
rect 26237 26333 26249 26367
rect 26283 26333 26295 26367
rect 26418 26364 26424 26376
rect 26379 26336 26424 26364
rect 26237 26327 26295 26333
rect 26252 26296 26280 26327
rect 26418 26324 26424 26336
rect 26476 26324 26482 26376
rect 26602 26324 26608 26376
rect 26660 26364 26666 26376
rect 26881 26367 26939 26373
rect 26881 26364 26893 26367
rect 26660 26336 26893 26364
rect 26660 26324 26666 26336
rect 26881 26333 26893 26336
rect 26927 26333 26939 26367
rect 27062 26364 27068 26376
rect 27023 26336 27068 26364
rect 26881 26327 26939 26333
rect 27062 26324 27068 26336
rect 27120 26324 27126 26376
rect 27154 26324 27160 26376
rect 27212 26364 27218 26376
rect 27297 26373 27325 26472
rect 27522 26432 27528 26444
rect 27483 26404 27528 26432
rect 27522 26392 27528 26404
rect 27580 26392 27586 26444
rect 27706 26392 27712 26444
rect 27764 26392 27770 26444
rect 27908 26432 27936 26540
rect 28000 26540 28908 26568
rect 28000 26509 28028 26540
rect 28902 26528 28908 26540
rect 28960 26528 28966 26580
rect 29362 26528 29368 26580
rect 29420 26568 29426 26580
rect 29733 26571 29791 26577
rect 29733 26568 29745 26571
rect 29420 26540 29745 26568
rect 29420 26528 29426 26540
rect 29733 26537 29745 26540
rect 29779 26537 29791 26571
rect 30926 26568 30932 26580
rect 30887 26540 30932 26568
rect 29733 26531 29791 26537
rect 30926 26528 30932 26540
rect 30984 26528 30990 26580
rect 27985 26503 28043 26509
rect 27985 26469 27997 26503
rect 28031 26469 28043 26503
rect 27985 26463 28043 26469
rect 28258 26460 28264 26512
rect 28316 26460 28322 26512
rect 28994 26460 29000 26512
rect 29052 26500 29058 26512
rect 29546 26500 29552 26512
rect 29052 26472 29552 26500
rect 29052 26460 29058 26472
rect 29546 26460 29552 26472
rect 29604 26460 29610 26512
rect 29822 26460 29828 26512
rect 29880 26500 29886 26512
rect 30098 26500 30104 26512
rect 29880 26472 30104 26500
rect 29880 26460 29886 26472
rect 30098 26460 30104 26472
rect 30156 26460 30162 26512
rect 30653 26503 30711 26509
rect 30653 26469 30665 26503
rect 30699 26500 30711 26503
rect 30834 26500 30840 26512
rect 30699 26472 30840 26500
rect 30699 26469 30711 26472
rect 30653 26463 30711 26469
rect 30834 26460 30840 26472
rect 30892 26460 30898 26512
rect 28074 26432 28080 26444
rect 27908 26404 28080 26432
rect 28074 26392 28080 26404
rect 28132 26392 28138 26444
rect 27295 26367 27353 26373
rect 27212 26336 27257 26364
rect 27212 26324 27218 26336
rect 27295 26333 27307 26367
rect 27341 26333 27353 26367
rect 27724 26364 27752 26392
rect 27890 26364 27896 26376
rect 27724 26336 27896 26364
rect 27295 26327 27353 26333
rect 27890 26324 27896 26336
rect 27948 26324 27954 26376
rect 28166 26364 28172 26376
rect 28127 26336 28172 26364
rect 28166 26324 28172 26336
rect 28224 26324 28230 26376
rect 28276 26373 28304 26460
rect 31202 26432 31208 26444
rect 30300 26404 31208 26432
rect 28261 26367 28319 26373
rect 28261 26333 28273 26367
rect 28307 26333 28319 26367
rect 28261 26327 28319 26333
rect 28353 26367 28411 26373
rect 28353 26333 28365 26367
rect 28399 26364 28411 26367
rect 28718 26364 28724 26376
rect 28399 26336 28724 26364
rect 28399 26333 28411 26336
rect 28353 26327 28411 26333
rect 28718 26324 28724 26336
rect 28776 26324 28782 26376
rect 28994 26364 29000 26376
rect 28955 26336 29000 26364
rect 28994 26324 29000 26336
rect 29052 26324 29058 26376
rect 29086 26324 29092 26376
rect 29144 26364 29150 26376
rect 29144 26336 29189 26364
rect 29144 26324 29150 26336
rect 29362 26324 29368 26376
rect 29420 26364 29426 26376
rect 29917 26367 29975 26373
rect 29917 26364 29929 26367
rect 29420 26336 29929 26364
rect 29420 26324 29426 26336
rect 29917 26333 29929 26336
rect 29963 26333 29975 26367
rect 29917 26327 29975 26333
rect 30193 26367 30251 26373
rect 30193 26333 30205 26367
rect 30239 26364 30251 26367
rect 30300 26364 30328 26404
rect 31202 26392 31208 26404
rect 31260 26392 31266 26444
rect 30834 26364 30840 26376
rect 30239 26336 30328 26364
rect 30795 26336 30840 26364
rect 30239 26333 30251 26336
rect 30193 26327 30251 26333
rect 27982 26296 27988 26308
rect 26252 26268 27988 26296
rect 27982 26256 27988 26268
rect 28040 26256 28046 26308
rect 28537 26299 28595 26305
rect 28537 26265 28549 26299
rect 28583 26296 28595 26299
rect 29822 26296 29828 26308
rect 28583 26268 29828 26296
rect 28583 26265 28595 26268
rect 28537 26259 28595 26265
rect 29822 26256 29828 26268
rect 29880 26256 29886 26308
rect 29932 26296 29960 26327
rect 30834 26324 30840 26336
rect 30892 26324 30898 26376
rect 31021 26367 31079 26373
rect 31021 26333 31033 26367
rect 31067 26364 31079 26367
rect 31478 26364 31484 26376
rect 31067 26336 31484 26364
rect 31067 26333 31079 26336
rect 31021 26327 31079 26333
rect 31478 26324 31484 26336
rect 31536 26324 31542 26376
rect 29932 26268 30880 26296
rect 30852 26240 30880 26268
rect 31846 26256 31852 26308
rect 31904 26296 31910 26308
rect 31904 26268 32260 26296
rect 31904 26256 31910 26268
rect 25774 26228 25780 26240
rect 25608 26200 25780 26228
rect 24949 26191 25007 26197
rect 25774 26188 25780 26200
rect 25832 26228 25838 26240
rect 29086 26228 29092 26240
rect 25832 26200 29092 26228
rect 25832 26188 25838 26200
rect 29086 26188 29092 26200
rect 29144 26228 29150 26240
rect 30101 26231 30159 26237
rect 30101 26228 30113 26231
rect 29144 26200 30113 26228
rect 29144 26188 29150 26200
rect 30101 26197 30113 26200
rect 30147 26197 30159 26231
rect 30101 26191 30159 26197
rect 30834 26188 30840 26240
rect 30892 26188 30898 26240
rect 30926 26188 30932 26240
rect 30984 26228 30990 26240
rect 31662 26228 31668 26240
rect 30984 26200 31668 26228
rect 30984 26188 30990 26200
rect 31662 26188 31668 26200
rect 31720 26188 31726 26240
rect 31754 26188 31760 26240
rect 31812 26228 31818 26240
rect 31812 26200 32168 26228
rect 31812 26188 31818 26200
rect 32140 26172 32168 26200
rect 1104 26138 31992 26160
rect 1104 26086 8632 26138
rect 8684 26086 8696 26138
rect 8748 26086 8760 26138
rect 8812 26086 8824 26138
rect 8876 26086 8888 26138
rect 8940 26086 16314 26138
rect 16366 26086 16378 26138
rect 16430 26086 16442 26138
rect 16494 26086 16506 26138
rect 16558 26086 16570 26138
rect 16622 26086 23996 26138
rect 24048 26086 24060 26138
rect 24112 26086 24124 26138
rect 24176 26086 24188 26138
rect 24240 26086 24252 26138
rect 24304 26086 31678 26138
rect 31730 26086 31742 26138
rect 31794 26086 31806 26138
rect 31858 26086 31870 26138
rect 31922 26086 31934 26138
rect 31986 26086 31992 26138
rect 32122 26120 32128 26172
rect 32180 26120 32186 26172
rect 1104 26064 31992 26086
rect 5445 26027 5503 26033
rect 5445 25993 5457 26027
rect 5491 26024 5503 26027
rect 7926 26024 7932 26036
rect 5491 25996 7932 26024
rect 5491 25993 5503 25996
rect 5445 25987 5503 25993
rect 7926 25984 7932 25996
rect 7984 26024 7990 26036
rect 11882 26024 11888 26036
rect 7984 25996 11888 26024
rect 7984 25984 7990 25996
rect 11882 25984 11888 25996
rect 11940 26024 11946 26036
rect 12161 26027 12219 26033
rect 12161 26024 12173 26027
rect 11940 25996 12173 26024
rect 11940 25984 11946 25996
rect 12161 25993 12173 25996
rect 12207 26024 12219 26027
rect 13722 26024 13728 26036
rect 12207 25996 13728 26024
rect 12207 25993 12219 25996
rect 12161 25987 12219 25993
rect 8941 25959 8999 25965
rect 8941 25925 8953 25959
rect 8987 25956 8999 25959
rect 11146 25956 11152 25968
rect 8987 25928 9674 25956
rect 11059 25928 11152 25956
rect 8987 25925 8999 25928
rect 8941 25919 8999 25925
rect 9646 25888 9674 25928
rect 11146 25916 11152 25928
rect 11204 25956 11210 25968
rect 11422 25956 11428 25968
rect 11204 25928 11428 25956
rect 11204 25916 11210 25928
rect 11422 25916 11428 25928
rect 11480 25916 11486 25968
rect 13538 25888 13544 25900
rect 9646 25860 13544 25888
rect 13538 25848 13544 25860
rect 13596 25848 13602 25900
rect 8570 25780 8576 25832
rect 8628 25820 8634 25832
rect 9493 25823 9551 25829
rect 9493 25820 9505 25823
rect 8628 25792 9505 25820
rect 8628 25780 8634 25792
rect 9493 25789 9505 25792
rect 9539 25820 9551 25823
rect 10045 25823 10103 25829
rect 10045 25820 10057 25823
rect 9539 25792 10057 25820
rect 9539 25789 9551 25792
rect 9493 25783 9551 25789
rect 10045 25789 10057 25792
rect 10091 25820 10103 25823
rect 10594 25820 10600 25832
rect 10091 25792 10600 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10594 25780 10600 25792
rect 10652 25780 10658 25832
rect 12158 25780 12164 25832
rect 12216 25820 12222 25832
rect 13078 25820 13084 25832
rect 12216 25792 13084 25820
rect 12216 25780 12222 25792
rect 13078 25780 13084 25792
rect 13136 25820 13142 25832
rect 13173 25823 13231 25829
rect 13173 25820 13185 25823
rect 13136 25792 13185 25820
rect 13136 25780 13142 25792
rect 13173 25789 13185 25792
rect 13219 25789 13231 25823
rect 13648 25820 13676 25996
rect 13722 25984 13728 25996
rect 13780 25984 13786 26036
rect 13817 26027 13875 26033
rect 13817 25993 13829 26027
rect 13863 26024 13875 26027
rect 13906 26024 13912 26036
rect 13863 25996 13912 26024
rect 13863 25993 13875 25996
rect 13817 25987 13875 25993
rect 13906 25984 13912 25996
rect 13964 25984 13970 26036
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 18690 26024 18696 26036
rect 16540 25996 18696 26024
rect 16540 25984 16546 25996
rect 18690 25984 18696 25996
rect 18748 25984 18754 26036
rect 22097 26027 22155 26033
rect 22097 26024 22109 26027
rect 19168 25996 22109 26024
rect 17497 25959 17555 25965
rect 13740 25928 17448 25956
rect 13740 25900 13768 25928
rect 13722 25848 13728 25900
rect 13780 25848 13786 25900
rect 14826 25888 14832 25900
rect 14787 25860 14832 25888
rect 14826 25848 14832 25860
rect 14884 25848 14890 25900
rect 15010 25888 15016 25900
rect 14971 25860 15016 25888
rect 15010 25848 15016 25860
rect 15068 25848 15074 25900
rect 15286 25848 15292 25900
rect 15344 25888 15350 25900
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 15344 25860 15485 25888
rect 15344 25848 15350 25860
rect 15473 25857 15485 25860
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25888 16175 25891
rect 16206 25888 16212 25900
rect 16163 25860 16212 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 16206 25848 16212 25860
rect 16264 25848 16270 25900
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25888 16359 25891
rect 16390 25888 16396 25900
rect 16347 25860 16396 25888
rect 16347 25857 16359 25860
rect 16301 25851 16359 25857
rect 16390 25848 16396 25860
rect 16448 25848 16454 25900
rect 16850 25848 16856 25900
rect 16908 25888 16914 25900
rect 17313 25891 17371 25897
rect 17313 25888 17325 25891
rect 16908 25860 17325 25888
rect 16908 25848 16914 25860
rect 17313 25857 17325 25860
rect 17359 25857 17371 25891
rect 17313 25851 17371 25857
rect 13906 25820 13912 25832
rect 13648 25792 13912 25820
rect 13173 25783 13231 25789
rect 13906 25780 13912 25792
rect 13964 25780 13970 25832
rect 15565 25823 15623 25829
rect 15565 25789 15577 25823
rect 15611 25820 15623 25823
rect 16666 25820 16672 25832
rect 15611 25792 16672 25820
rect 15611 25789 15623 25792
rect 15565 25783 15623 25789
rect 16666 25780 16672 25792
rect 16724 25780 16730 25832
rect 16758 25780 16764 25832
rect 16816 25820 16822 25832
rect 16942 25820 16948 25832
rect 16816 25792 16948 25820
rect 16816 25780 16822 25792
rect 16942 25780 16948 25792
rect 17000 25780 17006 25832
rect 5997 25755 6055 25761
rect 5997 25721 6009 25755
rect 6043 25752 6055 25755
rect 7650 25752 7656 25764
rect 6043 25724 7656 25752
rect 6043 25721 6055 25724
rect 5997 25715 6055 25721
rect 7650 25712 7656 25724
rect 7708 25712 7714 25764
rect 7837 25755 7895 25761
rect 7837 25721 7849 25755
rect 7883 25752 7895 25755
rect 9306 25752 9312 25764
rect 7883 25724 9312 25752
rect 7883 25721 7895 25724
rect 7837 25715 7895 25721
rect 9306 25712 9312 25724
rect 9364 25712 9370 25764
rect 11790 25712 11796 25764
rect 11848 25752 11854 25764
rect 14366 25752 14372 25764
rect 11848 25724 14372 25752
rect 11848 25712 11854 25724
rect 14366 25712 14372 25724
rect 14424 25712 14430 25764
rect 15013 25755 15071 25761
rect 15013 25721 15025 25755
rect 15059 25752 15071 25755
rect 17218 25752 17224 25764
rect 15059 25724 17224 25752
rect 15059 25721 15071 25724
rect 15013 25715 15071 25721
rect 17218 25712 17224 25724
rect 17276 25712 17282 25764
rect 17420 25752 17448 25928
rect 17497 25925 17509 25959
rect 17543 25956 17555 25959
rect 18230 25956 18236 25968
rect 17543 25928 18236 25956
rect 17543 25925 17555 25928
rect 17497 25919 17555 25925
rect 18230 25916 18236 25928
rect 18288 25916 18294 25968
rect 19168 25956 19196 25996
rect 22097 25993 22109 25996
rect 22143 25993 22155 26027
rect 22097 25987 22155 25993
rect 22281 26027 22339 26033
rect 22281 25993 22293 26027
rect 22327 25993 22339 26027
rect 22281 25987 22339 25993
rect 21358 25956 21364 25968
rect 18800 25928 19196 25956
rect 19536 25928 21364 25956
rect 17586 25848 17592 25900
rect 17644 25888 17650 25900
rect 18141 25894 18199 25897
rect 17972 25891 18199 25894
rect 17972 25888 18153 25891
rect 17644 25866 18153 25888
rect 17644 25860 18000 25866
rect 17644 25848 17650 25860
rect 18141 25857 18153 25866
rect 18187 25857 18199 25891
rect 18141 25851 18199 25857
rect 18325 25891 18383 25897
rect 18325 25857 18337 25891
rect 18371 25888 18383 25891
rect 18414 25888 18420 25900
rect 18371 25860 18420 25888
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 18414 25848 18420 25860
rect 18472 25848 18478 25900
rect 18230 25780 18236 25832
rect 18288 25820 18294 25832
rect 18800 25820 18828 25928
rect 18874 25848 18880 25900
rect 18932 25888 18938 25900
rect 19153 25894 19211 25897
rect 19076 25891 19211 25894
rect 19076 25888 19165 25891
rect 18932 25866 19165 25888
rect 18932 25860 19104 25866
rect 18932 25848 18938 25860
rect 19153 25857 19165 25866
rect 19199 25857 19211 25891
rect 19249 25858 19255 25910
rect 19307 25898 19313 25910
rect 19307 25888 19403 25898
rect 19441 25891 19499 25897
rect 19441 25888 19453 25891
rect 19307 25870 19453 25888
rect 19307 25858 19313 25870
rect 19375 25860 19453 25870
rect 19153 25851 19211 25857
rect 19441 25857 19453 25860
rect 19487 25857 19499 25891
rect 19441 25851 19499 25857
rect 18288 25792 18828 25820
rect 18969 25823 19027 25829
rect 18288 25780 18294 25792
rect 18969 25789 18981 25823
rect 19015 25820 19027 25823
rect 19058 25820 19064 25832
rect 19015 25792 19064 25820
rect 19015 25789 19027 25792
rect 18969 25783 19027 25789
rect 19058 25780 19064 25792
rect 19116 25780 19122 25832
rect 19536 25820 19564 25928
rect 19610 25848 19616 25900
rect 19668 25888 19674 25900
rect 20070 25888 20076 25900
rect 19668 25860 19932 25888
rect 20031 25860 20076 25888
rect 19668 25848 19674 25860
rect 19702 25820 19708 25832
rect 19168 25792 19564 25820
rect 19619 25792 19708 25820
rect 18509 25755 18567 25761
rect 17420 25724 18460 25752
rect 6733 25687 6791 25693
rect 6733 25653 6745 25687
rect 6779 25684 6791 25687
rect 7285 25687 7343 25693
rect 7285 25684 7297 25687
rect 6779 25656 7297 25684
rect 6779 25653 6791 25656
rect 6733 25647 6791 25653
rect 7285 25653 7297 25656
rect 7331 25684 7343 25687
rect 7466 25684 7472 25696
rect 7331 25656 7472 25684
rect 7331 25653 7343 25656
rect 7285 25647 7343 25653
rect 7466 25644 7472 25656
rect 7524 25644 7530 25696
rect 8110 25644 8116 25696
rect 8168 25684 8174 25696
rect 8389 25687 8447 25693
rect 8389 25684 8401 25687
rect 8168 25656 8401 25684
rect 8168 25644 8174 25656
rect 8389 25653 8401 25656
rect 8435 25684 8447 25687
rect 10597 25687 10655 25693
rect 10597 25684 10609 25687
rect 8435 25656 10609 25684
rect 8435 25653 8447 25656
rect 8389 25647 8447 25653
rect 10597 25653 10609 25656
rect 10643 25684 10655 25687
rect 12158 25684 12164 25696
rect 10643 25656 12164 25684
rect 10643 25653 10655 25656
rect 10597 25647 10655 25653
rect 12158 25644 12164 25656
rect 12216 25644 12222 25696
rect 12713 25687 12771 25693
rect 12713 25653 12725 25687
rect 12759 25684 12771 25687
rect 13446 25684 13452 25696
rect 12759 25656 13452 25684
rect 12759 25653 12771 25656
rect 12713 25647 12771 25653
rect 13446 25644 13452 25656
rect 13504 25644 13510 25696
rect 14274 25684 14280 25696
rect 14235 25656 14280 25684
rect 14274 25644 14280 25656
rect 14332 25644 14338 25696
rect 14642 25644 14648 25696
rect 14700 25684 14706 25696
rect 16209 25687 16267 25693
rect 16209 25684 16221 25687
rect 14700 25656 16221 25684
rect 14700 25644 14706 25656
rect 16209 25653 16221 25656
rect 16255 25653 16267 25687
rect 16209 25647 16267 25653
rect 16390 25644 16396 25696
rect 16448 25684 16454 25696
rect 17402 25684 17408 25696
rect 16448 25656 17408 25684
rect 16448 25644 16454 25656
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 17678 25684 17684 25696
rect 17639 25656 17684 25684
rect 17678 25644 17684 25656
rect 17736 25644 17742 25696
rect 17862 25644 17868 25696
rect 17920 25684 17926 25696
rect 18230 25684 18236 25696
rect 17920 25656 18236 25684
rect 17920 25644 17926 25656
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 18432 25684 18460 25724
rect 18509 25721 18521 25755
rect 18555 25752 18567 25755
rect 18598 25752 18604 25764
rect 18555 25724 18604 25752
rect 18555 25721 18567 25724
rect 18509 25715 18567 25721
rect 18598 25712 18604 25724
rect 18656 25712 18662 25764
rect 19168 25684 19196 25792
rect 19242 25712 19248 25764
rect 19300 25752 19306 25764
rect 19619 25752 19647 25792
rect 19702 25780 19708 25792
rect 19760 25780 19766 25832
rect 19904 25829 19932 25860
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20180 25897 20208 25928
rect 21358 25916 21364 25928
rect 21416 25916 21422 25968
rect 21726 25916 21732 25968
rect 21784 25956 21790 25968
rect 22296 25956 22324 25987
rect 22738 25984 22744 26036
rect 22796 26024 22802 26036
rect 23293 26027 23351 26033
rect 23293 26024 23305 26027
rect 22796 25996 23305 26024
rect 22796 25984 22802 25996
rect 23293 25993 23305 25996
rect 23339 25993 23351 26027
rect 25038 26024 25044 26036
rect 23293 25987 23351 25993
rect 23388 25996 25044 26024
rect 23388 25956 23416 25996
rect 25038 25984 25044 25996
rect 25096 25984 25102 26036
rect 25590 25984 25596 26036
rect 25648 26024 25654 26036
rect 25777 26027 25835 26033
rect 25777 26024 25789 26027
rect 25648 25996 25789 26024
rect 25648 25984 25654 25996
rect 25777 25993 25789 25996
rect 25823 25993 25835 26027
rect 25777 25987 25835 25993
rect 25869 26027 25927 26033
rect 25869 25993 25881 26027
rect 25915 26024 25927 26027
rect 28902 26024 28908 26036
rect 25915 25996 28908 26024
rect 25915 25993 25927 25996
rect 25869 25987 25927 25993
rect 28902 25984 28908 25996
rect 28960 25984 28966 26036
rect 29178 25984 29184 26036
rect 29236 26024 29242 26036
rect 29273 26027 29331 26033
rect 29273 26024 29285 26027
rect 29236 25996 29285 26024
rect 29236 25984 29242 25996
rect 29273 25993 29285 25996
rect 29319 25993 29331 26027
rect 30374 26024 30380 26036
rect 29273 25987 29331 25993
rect 29564 25996 30380 26024
rect 21784 25928 22324 25956
rect 23032 25928 23416 25956
rect 21784 25916 21790 25928
rect 20165 25891 20223 25897
rect 20165 25857 20177 25891
rect 20211 25857 20223 25891
rect 20165 25851 20223 25857
rect 20254 25848 20260 25900
rect 20312 25888 20318 25900
rect 20312 25860 20357 25888
rect 20312 25848 20318 25860
rect 20438 25848 20444 25900
rect 20496 25888 20502 25900
rect 20901 25891 20959 25897
rect 20901 25888 20913 25891
rect 20496 25860 20913 25888
rect 20496 25848 20502 25860
rect 20901 25857 20913 25860
rect 20947 25857 20959 25891
rect 20901 25851 20959 25857
rect 21100 25860 22094 25888
rect 19889 25823 19947 25829
rect 19889 25789 19901 25823
rect 19935 25789 19947 25823
rect 19889 25783 19947 25789
rect 20349 25823 20407 25829
rect 20349 25789 20361 25823
rect 20395 25820 20407 25823
rect 21100 25820 21128 25860
rect 20395 25792 21128 25820
rect 21177 25823 21235 25829
rect 20395 25789 20407 25792
rect 20349 25783 20407 25789
rect 21177 25789 21189 25823
rect 21223 25789 21235 25823
rect 21177 25783 21235 25789
rect 20438 25752 20444 25764
rect 19300 25724 19647 25752
rect 19719 25724 20444 25752
rect 19300 25712 19306 25724
rect 18432 25656 19196 25684
rect 19337 25687 19395 25693
rect 19337 25653 19349 25687
rect 19383 25684 19395 25687
rect 19426 25684 19432 25696
rect 19383 25656 19432 25684
rect 19383 25653 19395 25656
rect 19337 25647 19395 25653
rect 19426 25644 19432 25656
rect 19484 25644 19490 25696
rect 19518 25644 19524 25696
rect 19576 25684 19582 25696
rect 19719 25684 19747 25724
rect 20438 25712 20444 25724
rect 20496 25712 20502 25764
rect 20622 25712 20628 25764
rect 20680 25752 20686 25764
rect 20806 25752 20812 25764
rect 20680 25724 20812 25752
rect 20680 25712 20686 25724
rect 20806 25712 20812 25724
rect 20864 25712 20870 25764
rect 19576 25656 19747 25684
rect 19576 25644 19582 25656
rect 19794 25644 19800 25696
rect 19852 25684 19858 25696
rect 21192 25684 21220 25783
rect 21266 25780 21272 25832
rect 21324 25820 21330 25832
rect 21726 25820 21732 25832
rect 21324 25792 21732 25820
rect 21324 25780 21330 25792
rect 21726 25780 21732 25792
rect 21784 25780 21790 25832
rect 22066 25820 22094 25860
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22278 25891 22336 25897
rect 22278 25888 22290 25891
rect 22244 25860 22290 25888
rect 22244 25848 22250 25860
rect 22278 25857 22290 25860
rect 22324 25888 22336 25891
rect 23032 25888 23060 25928
rect 24486 25916 24492 25968
rect 24544 25956 24550 25968
rect 24765 25959 24823 25965
rect 24765 25956 24777 25959
rect 24544 25928 24777 25956
rect 24544 25916 24550 25928
rect 24765 25925 24777 25928
rect 24811 25925 24823 25959
rect 24765 25919 24823 25925
rect 25682 25916 25688 25968
rect 25740 25956 25746 25968
rect 26510 25956 26516 25968
rect 25740 25928 26516 25956
rect 25740 25916 25746 25928
rect 26510 25916 26516 25928
rect 26568 25916 26574 25968
rect 27706 25956 27712 25968
rect 27172 25928 27712 25956
rect 22324 25860 23060 25888
rect 22324 25857 22336 25860
rect 22278 25851 22336 25857
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 23164 25860 23690 25888
rect 23164 25848 23170 25860
rect 26050 25848 26056 25900
rect 26108 25888 26114 25900
rect 27062 25888 27068 25900
rect 26108 25860 27068 25888
rect 26108 25848 26114 25860
rect 27062 25848 27068 25860
rect 27120 25848 27126 25900
rect 27172 25897 27200 25928
rect 27706 25916 27712 25928
rect 27764 25916 27770 25968
rect 27801 25959 27859 25965
rect 27801 25925 27813 25959
rect 27847 25956 27859 25959
rect 29564 25956 29592 25996
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 30742 26024 30748 26036
rect 30703 25996 30748 26024
rect 30742 25984 30748 25996
rect 30800 25984 30806 26036
rect 27847 25928 29592 25956
rect 27847 25925 27859 25928
rect 27801 25919 27859 25925
rect 29638 25916 29644 25968
rect 29696 25956 29702 25968
rect 29696 25928 30328 25956
rect 29696 25916 29702 25928
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27341 25891 27399 25897
rect 27341 25888 27353 25891
rect 27157 25851 27215 25857
rect 27264 25860 27353 25888
rect 22066 25792 22508 25820
rect 21453 25755 21511 25761
rect 21453 25721 21465 25755
rect 21499 25752 21511 25755
rect 22370 25752 22376 25764
rect 21499 25724 22376 25752
rect 21499 25721 21511 25724
rect 21453 25715 21511 25721
rect 22370 25712 22376 25724
rect 22428 25712 22434 25764
rect 19852 25656 21220 25684
rect 21269 25687 21327 25693
rect 19852 25644 19858 25656
rect 21269 25653 21281 25687
rect 21315 25684 21327 25687
rect 21726 25684 21732 25696
rect 21315 25656 21732 25684
rect 21315 25653 21327 25656
rect 21269 25647 21327 25653
rect 21726 25644 21732 25656
rect 21784 25644 21790 25696
rect 21910 25644 21916 25696
rect 21968 25684 21974 25696
rect 22186 25684 22192 25696
rect 21968 25656 22192 25684
rect 21968 25644 21974 25656
rect 22186 25644 22192 25656
rect 22244 25644 22250 25696
rect 22480 25684 22508 25792
rect 22554 25780 22560 25832
rect 22612 25820 22618 25832
rect 22735 25823 22793 25829
rect 22735 25820 22747 25823
rect 22612 25792 22747 25820
rect 22612 25780 22618 25792
rect 22735 25789 22747 25792
rect 22781 25789 22793 25823
rect 24026 25820 24032 25832
rect 22735 25783 22793 25789
rect 23768 25792 24032 25820
rect 22649 25755 22707 25761
rect 22649 25721 22661 25755
rect 22695 25752 22707 25755
rect 23768 25752 23796 25792
rect 24026 25780 24032 25792
rect 24084 25780 24090 25832
rect 24762 25780 24768 25832
rect 24820 25820 24826 25832
rect 25041 25823 25099 25829
rect 25041 25820 25053 25823
rect 24820 25792 25053 25820
rect 24820 25780 24826 25792
rect 25041 25789 25053 25792
rect 25087 25789 25099 25823
rect 25041 25783 25099 25789
rect 25685 25823 25743 25829
rect 25685 25789 25697 25823
rect 25731 25820 25743 25823
rect 25958 25820 25964 25832
rect 25731 25792 25964 25820
rect 25731 25789 25743 25792
rect 25685 25783 25743 25789
rect 25958 25780 25964 25792
rect 26016 25780 26022 25832
rect 26142 25780 26148 25832
rect 26200 25820 26206 25832
rect 26510 25820 26516 25832
rect 26200 25792 26516 25820
rect 26200 25780 26206 25792
rect 26510 25780 26516 25792
rect 26568 25780 26574 25832
rect 27264 25820 27292 25860
rect 27341 25857 27353 25860
rect 27387 25857 27399 25891
rect 27341 25851 27399 25857
rect 27433 25891 27491 25897
rect 27433 25857 27445 25891
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 27172 25792 27292 25820
rect 27448 25820 27476 25851
rect 27522 25848 27528 25900
rect 27580 25888 27586 25900
rect 28629 25891 28687 25897
rect 28629 25888 28641 25891
rect 27580 25860 27625 25888
rect 27724 25860 28641 25888
rect 27580 25848 27586 25860
rect 27724 25832 27752 25860
rect 28629 25857 28641 25860
rect 28675 25888 28687 25891
rect 28810 25888 28816 25900
rect 28675 25860 28816 25888
rect 28675 25857 28687 25860
rect 28629 25851 28687 25857
rect 28810 25848 28816 25860
rect 28868 25848 28874 25900
rect 29457 25891 29515 25897
rect 29457 25857 29469 25891
rect 29503 25857 29515 25891
rect 29457 25851 29515 25857
rect 29549 25891 29607 25897
rect 29549 25857 29561 25891
rect 29595 25857 29607 25891
rect 29822 25888 29828 25900
rect 29783 25860 29828 25888
rect 29549 25851 29607 25857
rect 27614 25820 27620 25832
rect 27448 25792 27620 25820
rect 27172 25764 27200 25792
rect 27614 25780 27620 25792
rect 27672 25780 27678 25832
rect 27706 25780 27712 25832
rect 27764 25780 27770 25832
rect 28721 25823 28779 25829
rect 28721 25789 28733 25823
rect 28767 25820 28779 25823
rect 29178 25820 29184 25832
rect 28767 25792 29184 25820
rect 28767 25789 28779 25792
rect 28721 25783 28779 25789
rect 29178 25780 29184 25792
rect 29236 25780 29242 25832
rect 22695 25724 23796 25752
rect 22695 25721 22707 25724
rect 22649 25715 22707 25721
rect 25866 25712 25872 25764
rect 25924 25752 25930 25764
rect 26237 25755 26295 25761
rect 26237 25752 26249 25755
rect 25924 25724 26249 25752
rect 25924 25712 25930 25724
rect 26237 25721 26249 25724
rect 26283 25721 26295 25755
rect 26237 25715 26295 25721
rect 27154 25712 27160 25764
rect 27212 25712 27218 25764
rect 27430 25712 27436 25764
rect 27488 25752 27494 25764
rect 27798 25752 27804 25764
rect 27488 25724 27804 25752
rect 27488 25712 27494 25724
rect 27798 25712 27804 25724
rect 27856 25712 27862 25764
rect 28261 25755 28319 25761
rect 28261 25721 28273 25755
rect 28307 25721 28319 25755
rect 28261 25715 28319 25721
rect 24670 25684 24676 25696
rect 22480 25656 24676 25684
rect 24670 25644 24676 25656
rect 24728 25644 24734 25696
rect 25406 25644 25412 25696
rect 25464 25684 25470 25696
rect 25958 25684 25964 25696
rect 25464 25656 25964 25684
rect 25464 25644 25470 25656
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 26142 25644 26148 25696
rect 26200 25684 26206 25696
rect 28276 25684 28304 25715
rect 28350 25712 28356 25764
rect 28408 25752 28414 25764
rect 29270 25752 29276 25764
rect 28408 25724 29276 25752
rect 28408 25712 28414 25724
rect 29270 25712 29276 25724
rect 29328 25712 29334 25764
rect 26200 25656 28304 25684
rect 29472 25684 29500 25851
rect 29564 25752 29592 25851
rect 29822 25848 29828 25860
rect 29880 25848 29886 25900
rect 30300 25897 30328 25928
rect 30285 25891 30343 25897
rect 30285 25857 30297 25891
rect 30331 25857 30343 25891
rect 30285 25851 30343 25857
rect 30374 25848 30380 25900
rect 30432 25888 30438 25900
rect 30561 25891 30619 25897
rect 30432 25860 30477 25888
rect 30432 25848 30438 25860
rect 30561 25857 30573 25891
rect 30607 25888 30619 25891
rect 30926 25888 30932 25900
rect 30607 25860 30932 25888
rect 30607 25857 30619 25860
rect 30561 25851 30619 25857
rect 30926 25848 30932 25860
rect 30984 25848 30990 25900
rect 32232 25888 32260 26268
rect 31128 25860 32260 25888
rect 29730 25820 29736 25832
rect 29691 25792 29736 25820
rect 29730 25780 29736 25792
rect 29788 25780 29794 25832
rect 31128 25820 31156 25860
rect 30392 25792 31156 25820
rect 29638 25752 29644 25764
rect 29564 25724 29644 25752
rect 29638 25712 29644 25724
rect 29696 25712 29702 25764
rect 30392 25684 30420 25792
rect 31202 25780 31208 25832
rect 31260 25780 31266 25832
rect 30926 25712 30932 25764
rect 30984 25752 30990 25764
rect 31220 25752 31248 25780
rect 30984 25724 31248 25752
rect 30984 25712 30990 25724
rect 29472 25656 30420 25684
rect 26200 25644 26206 25656
rect 30466 25644 30472 25696
rect 30524 25684 30530 25696
rect 30742 25684 30748 25696
rect 30524 25656 30748 25684
rect 30524 25644 30530 25656
rect 30742 25644 30748 25656
rect 30800 25644 30806 25696
rect 31202 25684 31208 25696
rect 31163 25656 31208 25684
rect 31202 25644 31208 25656
rect 31260 25644 31266 25696
rect 1104 25594 31832 25616
rect 1104 25542 4791 25594
rect 4843 25542 4855 25594
rect 4907 25542 4919 25594
rect 4971 25542 4983 25594
rect 5035 25542 5047 25594
rect 5099 25542 12473 25594
rect 12525 25542 12537 25594
rect 12589 25542 12601 25594
rect 12653 25542 12665 25594
rect 12717 25542 12729 25594
rect 12781 25542 20155 25594
rect 20207 25542 20219 25594
rect 20271 25542 20283 25594
rect 20335 25542 20347 25594
rect 20399 25542 20411 25594
rect 20463 25542 27837 25594
rect 27889 25542 27901 25594
rect 27953 25542 27965 25594
rect 28017 25542 28029 25594
rect 28081 25542 28093 25594
rect 28145 25542 31832 25594
rect 1104 25520 31832 25542
rect 5261 25483 5319 25489
rect 5261 25449 5273 25483
rect 5307 25480 5319 25483
rect 6270 25480 6276 25492
rect 5307 25452 6276 25480
rect 5307 25449 5319 25452
rect 5261 25443 5319 25449
rect 6270 25440 6276 25452
rect 6328 25440 6334 25492
rect 6362 25440 6368 25492
rect 6420 25480 6426 25492
rect 7377 25483 7435 25489
rect 7377 25480 7389 25483
rect 6420 25452 7389 25480
rect 6420 25440 6426 25452
rect 7377 25449 7389 25452
rect 7423 25449 7435 25483
rect 7377 25443 7435 25449
rect 8021 25483 8079 25489
rect 8021 25449 8033 25483
rect 8067 25480 8079 25483
rect 8478 25480 8484 25492
rect 8067 25452 8484 25480
rect 8067 25449 8079 25452
rect 8021 25443 8079 25449
rect 8478 25440 8484 25452
rect 8536 25440 8542 25492
rect 10321 25483 10379 25489
rect 10321 25449 10333 25483
rect 10367 25480 10379 25483
rect 11238 25480 11244 25492
rect 10367 25452 11244 25480
rect 10367 25449 10379 25452
rect 10321 25443 10379 25449
rect 11238 25440 11244 25452
rect 11296 25480 11302 25492
rect 11606 25480 11612 25492
rect 11296 25452 11612 25480
rect 11296 25440 11302 25452
rect 11606 25440 11612 25452
rect 11664 25440 11670 25492
rect 11882 25480 11888 25492
rect 11843 25452 11888 25480
rect 11882 25440 11888 25452
rect 11940 25440 11946 25492
rect 13630 25480 13636 25492
rect 13591 25452 13636 25480
rect 13630 25440 13636 25452
rect 13688 25440 13694 25492
rect 14458 25480 14464 25492
rect 13740 25452 14464 25480
rect 6288 25412 6316 25440
rect 6822 25412 6828 25424
rect 6288 25384 6828 25412
rect 6822 25372 6828 25384
rect 6880 25372 6886 25424
rect 7466 25372 7472 25424
rect 7524 25412 7530 25424
rect 9769 25415 9827 25421
rect 9769 25412 9781 25415
rect 7524 25384 9781 25412
rect 7524 25372 7530 25384
rect 9769 25381 9781 25384
rect 9815 25412 9827 25415
rect 12802 25412 12808 25424
rect 9815 25384 12808 25412
rect 9815 25381 9827 25384
rect 9769 25375 9827 25381
rect 12802 25372 12808 25384
rect 12860 25372 12866 25424
rect 8573 25347 8631 25353
rect 8573 25313 8585 25347
rect 8619 25344 8631 25347
rect 9030 25344 9036 25356
rect 8619 25316 9036 25344
rect 8619 25313 8631 25316
rect 8573 25307 8631 25313
rect 9030 25304 9036 25316
rect 9088 25344 9094 25356
rect 11606 25344 11612 25356
rect 9088 25316 11612 25344
rect 9088 25304 9094 25316
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 13740 25344 13768 25452
rect 14458 25440 14464 25452
rect 14516 25440 14522 25492
rect 14737 25483 14795 25489
rect 14737 25449 14749 25483
rect 14783 25449 14795 25483
rect 14737 25443 14795 25449
rect 13906 25372 13912 25424
rect 13964 25372 13970 25424
rect 14274 25372 14280 25424
rect 14332 25412 14338 25424
rect 14752 25412 14780 25443
rect 15194 25440 15200 25492
rect 15252 25480 15258 25492
rect 15289 25483 15347 25489
rect 15289 25480 15301 25483
rect 15252 25452 15301 25480
rect 15252 25440 15258 25452
rect 15289 25449 15301 25452
rect 15335 25449 15347 25483
rect 16117 25483 16175 25489
rect 16117 25480 16129 25483
rect 15289 25443 15347 25449
rect 15948 25452 16129 25480
rect 15948 25424 15976 25452
rect 16117 25449 16129 25452
rect 16163 25449 16175 25483
rect 16758 25480 16764 25492
rect 16719 25452 16764 25480
rect 16117 25443 16175 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 17126 25480 17132 25492
rect 17087 25452 17132 25480
rect 17126 25440 17132 25452
rect 17184 25440 17190 25492
rect 17218 25440 17224 25492
rect 17276 25480 17282 25492
rect 17494 25480 17500 25492
rect 17276 25452 17500 25480
rect 17276 25440 17282 25452
rect 17494 25440 17500 25452
rect 17552 25440 17558 25492
rect 17770 25440 17776 25492
rect 17828 25480 17834 25492
rect 18414 25480 18420 25492
rect 17828 25452 18420 25480
rect 17828 25440 17834 25452
rect 18414 25440 18420 25452
rect 18472 25480 18478 25492
rect 18877 25483 18935 25489
rect 18877 25480 18889 25483
rect 18472 25452 18889 25480
rect 18472 25440 18478 25452
rect 18877 25449 18889 25452
rect 18923 25449 18935 25483
rect 20162 25480 20168 25492
rect 18877 25443 18935 25449
rect 18984 25452 20168 25480
rect 14332 25384 15693 25412
rect 14332 25372 14338 25384
rect 13556 25316 13768 25344
rect 13924 25344 13952 25372
rect 14734 25344 14740 25356
rect 13924 25316 14740 25344
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 11790 25276 11796 25288
rect 6963 25248 11796 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 13170 25236 13176 25288
rect 13228 25236 13234 25288
rect 13556 25285 13584 25316
rect 14734 25304 14740 25316
rect 14792 25344 14798 25356
rect 14792 25316 15424 25344
rect 14792 25304 14798 25316
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 13630 25236 13636 25288
rect 13688 25236 13694 25288
rect 14458 25236 14464 25288
rect 14516 25276 14522 25288
rect 14645 25279 14703 25285
rect 14645 25276 14657 25279
rect 14516 25248 14657 25276
rect 14516 25236 14522 25248
rect 14645 25245 14657 25248
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 14829 25279 14887 25285
rect 14829 25245 14841 25279
rect 14875 25245 14887 25279
rect 15277 25279 15335 25285
rect 15277 25276 15289 25279
rect 14829 25239 14887 25245
rect 15212 25248 15289 25276
rect 9217 25211 9275 25217
rect 9217 25177 9229 25211
rect 9263 25208 9275 25211
rect 10594 25208 10600 25220
rect 9263 25180 10600 25208
rect 9263 25177 9275 25180
rect 9217 25171 9275 25177
rect 10594 25168 10600 25180
rect 10652 25168 10658 25220
rect 12894 25168 12900 25220
rect 12952 25208 12958 25220
rect 13188 25208 13216 25236
rect 13648 25208 13676 25236
rect 14844 25208 14872 25239
rect 12952 25180 13584 25208
rect 13648 25180 14872 25208
rect 12952 25168 12958 25180
rect 5810 25140 5816 25152
rect 5771 25112 5816 25140
rect 5810 25100 5816 25112
rect 5868 25100 5874 25152
rect 9858 25100 9864 25152
rect 9916 25140 9922 25152
rect 10781 25143 10839 25149
rect 10781 25140 10793 25143
rect 9916 25112 10793 25140
rect 9916 25100 9922 25112
rect 10781 25109 10793 25112
rect 10827 25109 10839 25143
rect 11422 25140 11428 25152
rect 11383 25112 11428 25140
rect 10781 25103 10839 25109
rect 11422 25100 11428 25112
rect 11480 25100 11486 25152
rect 11790 25100 11796 25152
rect 11848 25140 11854 25152
rect 12437 25143 12495 25149
rect 12437 25140 12449 25143
rect 11848 25112 12449 25140
rect 11848 25100 11854 25112
rect 12437 25109 12449 25112
rect 12483 25109 12495 25143
rect 12437 25103 12495 25109
rect 13081 25143 13139 25149
rect 13081 25109 13093 25143
rect 13127 25140 13139 25143
rect 13170 25140 13176 25152
rect 13127 25112 13176 25140
rect 13127 25109 13139 25112
rect 13081 25103 13139 25109
rect 13170 25100 13176 25112
rect 13228 25100 13234 25152
rect 13556 25140 13584 25180
rect 15212 25152 15240 25248
rect 15277 25245 15289 25248
rect 15323 25245 15335 25279
rect 15277 25239 15335 25245
rect 15396 25208 15424 25316
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25276 15531 25279
rect 15562 25276 15568 25288
rect 15519 25248 15568 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 15562 25236 15568 25248
rect 15620 25236 15626 25288
rect 15665 25276 15693 25384
rect 15930 25372 15936 25424
rect 15988 25372 15994 25424
rect 16301 25415 16359 25421
rect 16301 25381 16313 25415
rect 16347 25412 16359 25415
rect 16482 25412 16488 25424
rect 16347 25384 16488 25412
rect 16347 25381 16359 25384
rect 16301 25375 16359 25381
rect 16482 25372 16488 25384
rect 16540 25372 16546 25424
rect 16574 25372 16580 25424
rect 16632 25412 16638 25424
rect 17310 25412 17316 25424
rect 16632 25384 17316 25412
rect 16632 25372 16638 25384
rect 17310 25372 17316 25384
rect 17368 25372 17374 25424
rect 16206 25304 16212 25356
rect 16264 25344 16270 25356
rect 17788 25344 17816 25440
rect 18984 25412 19012 25452
rect 20162 25440 20168 25452
rect 20220 25480 20226 25492
rect 20349 25483 20407 25489
rect 20349 25480 20361 25483
rect 20220 25452 20361 25480
rect 20220 25440 20226 25452
rect 20349 25449 20361 25452
rect 20395 25449 20407 25483
rect 21174 25480 21180 25492
rect 21135 25452 21180 25480
rect 20349 25443 20407 25449
rect 21174 25440 21180 25452
rect 21232 25440 21238 25492
rect 21284 25452 21494 25480
rect 16264 25316 16712 25344
rect 16264 25304 16270 25316
rect 15665 25248 16574 25276
rect 15933 25211 15991 25217
rect 15933 25208 15945 25211
rect 15396 25180 15945 25208
rect 15933 25177 15945 25180
rect 15979 25177 15991 25211
rect 15933 25171 15991 25177
rect 13630 25140 13636 25152
rect 13556 25112 13636 25140
rect 13630 25100 13636 25112
rect 13688 25100 13694 25152
rect 15194 25100 15200 25152
rect 15252 25100 15258 25152
rect 15654 25100 15660 25152
rect 15712 25140 15718 25152
rect 16133 25143 16191 25149
rect 16133 25140 16145 25143
rect 15712 25112 16145 25140
rect 15712 25100 15718 25112
rect 16133 25109 16145 25112
rect 16179 25109 16191 25143
rect 16546 25140 16574 25248
rect 16684 25208 16712 25316
rect 16776 25316 17816 25344
rect 17906 25384 19012 25412
rect 19267 25384 19938 25412
rect 16776 25285 16804 25316
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25245 16819 25279
rect 16761 25239 16819 25245
rect 16945 25279 17003 25285
rect 16945 25245 16957 25279
rect 16991 25276 17003 25279
rect 17310 25276 17316 25288
rect 16991 25248 17316 25276
rect 16991 25245 17003 25248
rect 16945 25239 17003 25245
rect 17310 25236 17316 25248
rect 17368 25236 17374 25288
rect 17494 25236 17500 25288
rect 17552 25276 17558 25288
rect 17589 25279 17647 25285
rect 17589 25276 17601 25279
rect 17552 25248 17601 25276
rect 17552 25236 17558 25248
rect 17589 25245 17601 25248
rect 17635 25245 17647 25279
rect 17906 25278 17934 25384
rect 19150 25344 19156 25356
rect 17880 25276 17934 25278
rect 17589 25239 17647 25245
rect 17788 25250 17934 25276
rect 17972 25316 19156 25344
rect 17788 25248 17908 25250
rect 17788 25217 17816 25248
rect 17773 25211 17831 25217
rect 17773 25208 17785 25211
rect 16684 25180 17785 25208
rect 17773 25177 17785 25180
rect 17819 25177 17831 25211
rect 17773 25171 17831 25177
rect 17862 25168 17868 25220
rect 17920 25208 17926 25220
rect 17972 25208 18000 25316
rect 19150 25304 19156 25316
rect 19208 25304 19214 25356
rect 18322 25236 18328 25288
rect 18380 25276 18386 25288
rect 18417 25279 18475 25285
rect 18417 25276 18429 25279
rect 18380 25248 18429 25276
rect 18380 25236 18386 25248
rect 18417 25245 18429 25248
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18506 25236 18512 25288
rect 18564 25285 18570 25288
rect 18564 25279 18593 25285
rect 18581 25245 18593 25279
rect 18564 25239 18593 25245
rect 18564 25236 18570 25239
rect 18782 25236 18788 25288
rect 18840 25276 18846 25288
rect 19267 25276 19295 25384
rect 19334 25304 19340 25356
rect 19392 25344 19398 25356
rect 19632 25347 19690 25353
rect 19632 25344 19644 25347
rect 19392 25316 19644 25344
rect 19392 25304 19398 25316
rect 19632 25313 19644 25316
rect 19678 25313 19690 25347
rect 19910 25344 19938 25384
rect 19978 25372 19984 25424
rect 20036 25412 20042 25424
rect 20438 25412 20444 25424
rect 20036 25384 20444 25412
rect 20036 25372 20042 25384
rect 20438 25372 20444 25384
rect 20496 25372 20502 25424
rect 20530 25372 20536 25424
rect 20588 25412 20594 25424
rect 21284 25412 21312 25452
rect 20588 25384 21312 25412
rect 20588 25372 20594 25384
rect 21358 25372 21364 25424
rect 21416 25372 21422 25424
rect 21466 25412 21494 25452
rect 21542 25440 21548 25492
rect 21600 25480 21606 25492
rect 23658 25480 23664 25492
rect 21600 25452 23664 25480
rect 21600 25440 21606 25452
rect 23658 25440 23664 25452
rect 23716 25440 23722 25492
rect 23934 25440 23940 25492
rect 23992 25480 23998 25492
rect 24029 25483 24087 25489
rect 24029 25480 24041 25483
rect 23992 25452 24041 25480
rect 23992 25440 23998 25452
rect 24029 25449 24041 25452
rect 24075 25449 24087 25483
rect 24029 25443 24087 25449
rect 24118 25440 24124 25492
rect 24176 25480 24182 25492
rect 24854 25480 24860 25492
rect 24176 25452 24860 25480
rect 24176 25440 24182 25452
rect 24854 25440 24860 25452
rect 24912 25440 24918 25492
rect 24946 25440 24952 25492
rect 25004 25480 25010 25492
rect 25004 25452 26262 25480
rect 25004 25440 25010 25452
rect 21466 25384 21588 25412
rect 21266 25344 21272 25356
rect 19910 25316 21272 25344
rect 19632 25307 19690 25313
rect 21266 25304 21272 25316
rect 21324 25304 21330 25356
rect 21376 25344 21404 25372
rect 21453 25347 21511 25353
rect 21453 25344 21465 25347
rect 21376 25316 21465 25344
rect 21453 25313 21465 25316
rect 21499 25313 21511 25347
rect 21560 25344 21588 25384
rect 22002 25372 22008 25424
rect 22060 25412 22066 25424
rect 22278 25412 22284 25424
rect 22060 25384 22284 25412
rect 22060 25372 22066 25384
rect 22278 25372 22284 25384
rect 22336 25372 22342 25424
rect 23750 25372 23756 25424
rect 23808 25412 23814 25424
rect 24578 25412 24584 25424
rect 23808 25384 24584 25412
rect 23808 25372 23814 25384
rect 24578 25372 24584 25384
rect 24636 25372 24642 25424
rect 25958 25372 25964 25424
rect 26016 25412 26022 25424
rect 26234 25412 26262 25452
rect 26418 25440 26424 25492
rect 26476 25480 26482 25492
rect 26881 25483 26939 25489
rect 26881 25480 26893 25483
rect 26476 25452 26893 25480
rect 26476 25440 26482 25452
rect 26881 25449 26893 25452
rect 26927 25449 26939 25483
rect 27982 25480 27988 25492
rect 26881 25443 26939 25449
rect 26977 25452 27988 25480
rect 26977 25412 27005 25452
rect 27982 25440 27988 25452
rect 28040 25440 28046 25492
rect 28445 25483 28503 25489
rect 28445 25449 28457 25483
rect 28491 25480 28503 25483
rect 29638 25480 29644 25492
rect 28491 25452 29644 25480
rect 28491 25449 28503 25452
rect 28445 25443 28503 25449
rect 29638 25440 29644 25452
rect 29696 25440 29702 25492
rect 29730 25440 29736 25492
rect 29788 25480 29794 25492
rect 29917 25483 29975 25489
rect 29917 25480 29929 25483
rect 29788 25452 29929 25480
rect 29788 25440 29794 25452
rect 29917 25449 29929 25452
rect 29963 25480 29975 25483
rect 30926 25480 30932 25492
rect 29963 25452 30696 25480
rect 30887 25452 30932 25480
rect 29963 25449 29975 25452
rect 29917 25443 29975 25449
rect 26016 25384 26197 25412
rect 26234 25384 27005 25412
rect 26016 25372 26022 25384
rect 22557 25347 22615 25353
rect 22557 25344 22569 25347
rect 21560 25316 22569 25344
rect 21453 25307 21511 25313
rect 22557 25313 22569 25316
rect 22603 25313 22615 25347
rect 22557 25307 22615 25313
rect 22646 25304 22652 25356
rect 22704 25344 22710 25356
rect 23106 25344 23112 25356
rect 22704 25316 23112 25344
rect 22704 25304 22710 25316
rect 23106 25304 23112 25316
rect 23164 25304 23170 25356
rect 23198 25304 23204 25356
rect 23256 25344 23262 25356
rect 24857 25347 24915 25353
rect 24857 25344 24869 25347
rect 23256 25316 24869 25344
rect 23256 25304 23262 25316
rect 24857 25313 24869 25316
rect 24903 25313 24915 25347
rect 24857 25307 24915 25313
rect 25222 25304 25228 25356
rect 25280 25344 25286 25356
rect 26169 25344 26197 25384
rect 27062 25372 27068 25424
rect 27120 25372 27126 25424
rect 27246 25372 27252 25424
rect 27304 25412 27310 25424
rect 28629 25415 28687 25421
rect 27304 25384 28580 25412
rect 27304 25372 27310 25384
rect 27080 25344 27108 25372
rect 25280 25316 26092 25344
rect 26169 25316 27420 25344
rect 25280 25304 25286 25316
rect 19426 25276 19432 25288
rect 18840 25248 19295 25276
rect 19387 25248 19432 25276
rect 18840 25236 18846 25248
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 19518 25236 19524 25288
rect 19576 25276 19582 25288
rect 20346 25276 20352 25288
rect 19576 25248 19621 25276
rect 20307 25248 20352 25276
rect 19576 25236 19582 25248
rect 20346 25236 20352 25248
rect 20404 25236 20410 25288
rect 20717 25279 20775 25285
rect 20717 25245 20729 25279
rect 20763 25276 20775 25279
rect 20763 25248 20852 25276
rect 20763 25245 20775 25248
rect 20717 25239 20775 25245
rect 17920 25180 18000 25208
rect 17920 25168 17926 25180
rect 18230 25168 18236 25220
rect 18288 25208 18294 25220
rect 18288 25180 18920 25208
rect 18288 25168 18294 25180
rect 16758 25140 16764 25152
rect 16546 25112 16764 25140
rect 16133 25103 16191 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 17402 25100 17408 25152
rect 17460 25140 17466 25152
rect 17957 25143 18015 25149
rect 17957 25140 17969 25143
rect 17460 25112 17969 25140
rect 17460 25100 17466 25112
rect 17957 25109 17969 25112
rect 18003 25109 18015 25143
rect 17957 25103 18015 25109
rect 18046 25100 18052 25152
rect 18104 25140 18110 25152
rect 18598 25140 18604 25152
rect 18104 25112 18604 25140
rect 18104 25100 18110 25112
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 18693 25143 18751 25149
rect 18693 25109 18705 25143
rect 18739 25140 18751 25143
rect 18782 25140 18788 25152
rect 18739 25112 18788 25140
rect 18739 25109 18751 25112
rect 18693 25103 18751 25109
rect 18782 25100 18788 25112
rect 18840 25100 18846 25152
rect 18892 25140 18920 25180
rect 19334 25168 19340 25220
rect 19392 25208 19398 25220
rect 19610 25208 19616 25220
rect 19392 25180 19616 25208
rect 19392 25168 19398 25180
rect 19610 25168 19616 25180
rect 19668 25208 19674 25220
rect 19705 25211 19763 25217
rect 19705 25208 19717 25211
rect 19668 25180 19717 25208
rect 19668 25168 19674 25180
rect 19705 25177 19717 25180
rect 19751 25177 19763 25211
rect 19705 25171 19763 25177
rect 19886 25168 19892 25220
rect 19944 25208 19950 25220
rect 20530 25208 20536 25220
rect 19944 25180 20536 25208
rect 19944 25168 19950 25180
rect 20530 25168 20536 25180
rect 20588 25168 20594 25220
rect 20165 25143 20223 25149
rect 20165 25140 20177 25143
rect 18892 25112 20177 25140
rect 20165 25109 20177 25112
rect 20211 25109 20223 25143
rect 20165 25103 20223 25109
rect 20714 25100 20720 25152
rect 20772 25140 20778 25152
rect 20824 25140 20852 25248
rect 20898 25236 20904 25288
rect 20956 25276 20962 25288
rect 21361 25279 21419 25285
rect 21361 25276 21373 25279
rect 20956 25248 21373 25276
rect 20956 25236 20962 25248
rect 21361 25245 21373 25248
rect 21407 25245 21419 25279
rect 21545 25279 21603 25285
rect 21545 25276 21557 25279
rect 21361 25239 21419 25245
rect 21468 25248 21557 25276
rect 20990 25168 20996 25220
rect 21048 25208 21054 25220
rect 21468 25208 21496 25248
rect 21545 25245 21557 25248
rect 21591 25245 21603 25279
rect 21545 25239 21603 25245
rect 21637 25279 21695 25285
rect 21637 25245 21649 25279
rect 21683 25245 21695 25279
rect 21637 25239 21695 25245
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25245 21879 25279
rect 22278 25276 22284 25288
rect 22239 25248 22284 25276
rect 21821 25239 21879 25245
rect 21652 25208 21680 25239
rect 21048 25180 21496 25208
rect 21560 25180 21680 25208
rect 21836 25208 21864 25239
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 24302 25276 24308 25288
rect 23690 25248 24308 25276
rect 24302 25236 24308 25248
rect 24360 25236 24366 25288
rect 24578 25276 24584 25288
rect 24539 25248 24584 25276
rect 24578 25236 24584 25248
rect 24636 25236 24642 25288
rect 26064 25276 26092 25316
rect 26064 25248 26556 25276
rect 22646 25208 22652 25220
rect 21836 25180 22652 25208
rect 21048 25168 21054 25180
rect 21376 25152 21404 25180
rect 21560 25152 21588 25180
rect 22646 25168 22652 25180
rect 22704 25168 22710 25220
rect 23828 25180 25346 25208
rect 20772 25112 20852 25140
rect 20772 25100 20778 25112
rect 21358 25100 21364 25152
rect 21416 25100 21422 25152
rect 21542 25100 21548 25152
rect 21600 25100 21606 25152
rect 22002 25100 22008 25152
rect 22060 25140 22066 25152
rect 23198 25140 23204 25152
rect 22060 25112 23204 25140
rect 22060 25100 22066 25112
rect 23198 25100 23204 25112
rect 23256 25100 23262 25152
rect 23566 25100 23572 25152
rect 23624 25140 23630 25152
rect 23828 25140 23856 25180
rect 23624 25112 23856 25140
rect 23624 25100 23630 25112
rect 24210 25100 24216 25152
rect 24268 25140 24274 25152
rect 24854 25140 24860 25152
rect 24268 25112 24860 25140
rect 24268 25100 24274 25112
rect 24854 25100 24860 25112
rect 24912 25100 24918 25152
rect 25130 25100 25136 25152
rect 25188 25140 25194 25152
rect 26329 25143 26387 25149
rect 26329 25140 26341 25143
rect 25188 25112 26341 25140
rect 25188 25100 25194 25112
rect 26329 25109 26341 25112
rect 26375 25140 26387 25143
rect 26418 25140 26424 25152
rect 26375 25112 26424 25140
rect 26375 25109 26387 25112
rect 26329 25103 26387 25109
rect 26418 25100 26424 25112
rect 26476 25100 26482 25152
rect 26528 25140 26556 25248
rect 26970 25236 26976 25288
rect 27028 25285 27034 25288
rect 27028 25279 27077 25285
rect 27028 25245 27031 25279
rect 27065 25245 27077 25279
rect 27154 25276 27160 25288
rect 27115 25248 27160 25276
rect 27028 25239 27077 25245
rect 27028 25236 27034 25239
rect 27154 25236 27160 25248
rect 27212 25236 27218 25288
rect 27246 25236 27252 25288
rect 27304 25276 27310 25288
rect 27392 25285 27420 25316
rect 27798 25304 27804 25356
rect 27856 25344 27862 25356
rect 28261 25347 28319 25353
rect 28261 25344 28273 25347
rect 27856 25316 28273 25344
rect 27856 25304 27862 25316
rect 28261 25313 28273 25316
rect 28307 25313 28319 25347
rect 28552 25344 28580 25384
rect 28629 25381 28641 25415
rect 28675 25412 28687 25415
rect 30558 25412 30564 25424
rect 28675 25384 30564 25412
rect 28675 25381 28687 25384
rect 28629 25375 28687 25381
rect 30558 25372 30564 25384
rect 30616 25372 30622 25424
rect 30374 25344 30380 25356
rect 28552 25316 30380 25344
rect 28261 25307 28319 25313
rect 30374 25304 30380 25316
rect 30432 25304 30438 25356
rect 27377 25279 27435 25285
rect 27304 25248 27349 25276
rect 27304 25236 27310 25248
rect 27377 25245 27389 25279
rect 27423 25245 27435 25279
rect 27377 25239 27435 25245
rect 27525 25279 27583 25285
rect 27525 25245 27537 25279
rect 27571 25276 27583 25279
rect 27706 25276 27712 25288
rect 27571 25248 27712 25276
rect 27571 25245 27583 25248
rect 27525 25239 27583 25245
rect 27706 25236 27712 25248
rect 27764 25236 27770 25288
rect 27985 25279 28043 25285
rect 27985 25245 27997 25279
rect 28031 25276 28043 25279
rect 28166 25276 28172 25288
rect 28031 25248 28172 25276
rect 28031 25245 28043 25248
rect 27985 25239 28043 25245
rect 28166 25236 28172 25248
rect 28224 25236 28230 25288
rect 28445 25279 28503 25285
rect 28445 25245 28457 25279
rect 28491 25245 28503 25279
rect 28445 25239 28503 25245
rect 26694 25168 26700 25220
rect 26752 25208 26758 25220
rect 28258 25208 28264 25220
rect 26752 25180 28264 25208
rect 26752 25168 26758 25180
rect 28258 25168 28264 25180
rect 28316 25208 28322 25220
rect 28460 25208 28488 25239
rect 28810 25236 28816 25288
rect 28868 25276 28874 25288
rect 29822 25276 29828 25288
rect 28868 25248 29828 25276
rect 28868 25236 28874 25248
rect 29822 25236 29828 25248
rect 29880 25276 29886 25288
rect 29917 25279 29975 25285
rect 29917 25276 29929 25279
rect 29880 25248 29929 25276
rect 29880 25236 29886 25248
rect 29917 25245 29929 25248
rect 29963 25245 29975 25279
rect 29917 25239 29975 25245
rect 30098 25236 30104 25288
rect 30156 25276 30162 25288
rect 30285 25279 30343 25285
rect 30285 25276 30297 25279
rect 30156 25248 30297 25276
rect 30156 25236 30162 25248
rect 30285 25245 30297 25248
rect 30331 25245 30343 25279
rect 30285 25239 30343 25245
rect 30558 25236 30564 25288
rect 30616 25276 30622 25288
rect 30668 25276 30696 25452
rect 30926 25440 30932 25452
rect 30984 25440 30990 25492
rect 30834 25372 30840 25424
rect 30892 25412 30898 25424
rect 31297 25415 31355 25421
rect 31297 25412 31309 25415
rect 30892 25384 31309 25412
rect 30892 25372 30898 25384
rect 31297 25381 31309 25384
rect 31343 25381 31355 25415
rect 31297 25375 31355 25381
rect 30616 25248 30696 25276
rect 30616 25236 30622 25248
rect 29178 25208 29184 25220
rect 28316 25180 28488 25208
rect 29139 25180 29184 25208
rect 28316 25168 28322 25180
rect 29178 25168 29184 25180
rect 29236 25168 29242 25220
rect 29288 25180 30788 25208
rect 29288 25140 29316 25180
rect 29730 25140 29736 25152
rect 26528 25112 29316 25140
rect 29691 25112 29736 25140
rect 29730 25100 29736 25112
rect 29788 25100 29794 25152
rect 30760 25149 30788 25180
rect 30745 25143 30803 25149
rect 30745 25109 30757 25143
rect 30791 25109 30803 25143
rect 30745 25103 30803 25109
rect 30834 25100 30840 25152
rect 30892 25140 30898 25152
rect 30929 25143 30987 25149
rect 30929 25140 30941 25143
rect 30892 25112 30941 25140
rect 30892 25100 30898 25112
rect 30929 25109 30941 25112
rect 30975 25109 30987 25143
rect 30929 25103 30987 25109
rect 1104 25050 31992 25072
rect 1104 24998 8632 25050
rect 8684 24998 8696 25050
rect 8748 24998 8760 25050
rect 8812 24998 8824 25050
rect 8876 24998 8888 25050
rect 8940 24998 16314 25050
rect 16366 24998 16378 25050
rect 16430 24998 16442 25050
rect 16494 24998 16506 25050
rect 16558 24998 16570 25050
rect 16622 24998 23996 25050
rect 24048 24998 24060 25050
rect 24112 24998 24124 25050
rect 24176 24998 24188 25050
rect 24240 24998 24252 25050
rect 24304 24998 31678 25050
rect 31730 24998 31742 25050
rect 31794 24998 31806 25050
rect 31858 24998 31870 25050
rect 31922 24998 31934 25050
rect 31986 24998 31992 25050
rect 1104 24976 31992 24998
rect 10045 24939 10103 24945
rect 10045 24905 10057 24939
rect 10091 24936 10103 24939
rect 11422 24936 11428 24948
rect 10091 24908 11428 24936
rect 10091 24905 10103 24908
rect 10045 24899 10103 24905
rect 11422 24896 11428 24908
rect 11480 24896 11486 24948
rect 12069 24939 12127 24945
rect 12069 24905 12081 24939
rect 12115 24936 12127 24939
rect 12158 24936 12164 24948
rect 12115 24908 12164 24936
rect 12115 24905 12127 24908
rect 12069 24899 12127 24905
rect 12158 24896 12164 24908
rect 12216 24896 12222 24948
rect 13173 24939 13231 24945
rect 13173 24905 13185 24939
rect 13219 24936 13231 24939
rect 13354 24936 13360 24948
rect 13219 24908 13360 24936
rect 13219 24905 13231 24908
rect 13173 24899 13231 24905
rect 13354 24896 13360 24908
rect 13412 24896 13418 24948
rect 14734 24896 14740 24948
rect 14792 24936 14798 24948
rect 14792 24908 15608 24936
rect 14792 24896 14798 24908
rect 4246 24828 4252 24880
rect 4304 24868 4310 24880
rect 12894 24868 12900 24880
rect 4304 24840 11100 24868
rect 4304 24828 4310 24840
rect 4893 24803 4951 24809
rect 4893 24769 4905 24803
rect 4939 24800 4951 24803
rect 5166 24800 5172 24812
rect 4939 24772 5172 24800
rect 4939 24769 4951 24772
rect 4893 24763 4951 24769
rect 5166 24760 5172 24772
rect 5224 24760 5230 24812
rect 5445 24803 5503 24809
rect 5445 24769 5457 24803
rect 5491 24800 5503 24803
rect 8386 24800 8392 24812
rect 5491 24772 8392 24800
rect 5491 24769 5503 24772
rect 5445 24763 5503 24769
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 9306 24760 9312 24812
rect 9364 24800 9370 24812
rect 9401 24803 9459 24809
rect 9401 24800 9413 24803
rect 9364 24772 9413 24800
rect 9364 24760 9370 24772
rect 9401 24769 9413 24772
rect 9447 24769 9459 24803
rect 9401 24763 9459 24769
rect 9582 24760 9588 24812
rect 9640 24800 9646 24812
rect 11072 24800 11100 24840
rect 11532 24840 12900 24868
rect 11532 24800 11560 24840
rect 12894 24828 12900 24840
rect 12952 24828 12958 24880
rect 14826 24868 14832 24880
rect 13280 24840 14832 24868
rect 13280 24812 13308 24840
rect 14826 24828 14832 24840
rect 14884 24868 14890 24880
rect 15105 24871 15163 24877
rect 15105 24868 15117 24871
rect 14884 24840 15117 24868
rect 14884 24828 14890 24840
rect 15105 24837 15117 24840
rect 15151 24837 15163 24871
rect 15378 24868 15384 24880
rect 15105 24831 15163 24837
rect 15228 24840 15384 24868
rect 9640 24772 11008 24800
rect 11072 24772 11560 24800
rect 9640 24760 9646 24772
rect 4338 24692 4344 24744
rect 4396 24732 4402 24744
rect 7285 24735 7343 24741
rect 7285 24732 7297 24735
rect 4396 24704 7297 24732
rect 4396 24692 4402 24704
rect 7285 24701 7297 24704
rect 7331 24732 7343 24735
rect 10226 24732 10232 24744
rect 7331 24704 10232 24732
rect 7331 24701 7343 24704
rect 7285 24695 7343 24701
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 10980 24732 11008 24772
rect 12710 24760 12716 24812
rect 12768 24800 12774 24812
rect 13081 24803 13139 24809
rect 13081 24800 13093 24803
rect 12768 24772 13093 24800
rect 12768 24760 12774 24772
rect 13081 24769 13093 24772
rect 13127 24769 13139 24803
rect 13262 24800 13268 24812
rect 13223 24772 13268 24800
rect 13081 24763 13139 24769
rect 13262 24760 13268 24772
rect 13320 24760 13326 24812
rect 13722 24800 13728 24812
rect 13683 24772 13728 24800
rect 13722 24760 13728 24772
rect 13780 24760 13786 24812
rect 14274 24760 14280 24812
rect 14332 24800 14338 24812
rect 14369 24803 14427 24809
rect 14369 24800 14381 24803
rect 14332 24772 14381 24800
rect 14332 24760 14338 24772
rect 14369 24769 14381 24772
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 14461 24803 14519 24809
rect 14461 24769 14473 24803
rect 14507 24769 14519 24803
rect 14461 24763 14519 24769
rect 14655 24803 14713 24809
rect 14655 24769 14667 24803
rect 14701 24800 14713 24803
rect 15228 24800 15256 24840
rect 15378 24828 15384 24840
rect 15436 24828 15442 24880
rect 15580 24868 15608 24908
rect 15654 24896 15660 24948
rect 15712 24936 15718 24948
rect 20162 24936 20168 24948
rect 15712 24908 20168 24936
rect 15712 24896 15718 24908
rect 20162 24896 20168 24908
rect 20220 24896 20226 24948
rect 20530 24896 20536 24948
rect 20588 24936 20594 24948
rect 20990 24936 20996 24948
rect 20588 24908 20996 24936
rect 20588 24896 20594 24908
rect 20990 24896 20996 24908
rect 21048 24896 21054 24948
rect 21177 24939 21235 24945
rect 21177 24905 21189 24939
rect 21223 24936 21235 24939
rect 21910 24936 21916 24948
rect 21223 24908 21916 24936
rect 21223 24905 21235 24908
rect 21177 24899 21235 24905
rect 15930 24868 15936 24880
rect 15580 24840 15700 24868
rect 15891 24840 15936 24868
rect 14701 24772 15256 24800
rect 15289 24803 15347 24809
rect 14701 24769 14713 24772
rect 14655 24763 14713 24769
rect 15289 24769 15301 24803
rect 15335 24800 15347 24803
rect 15562 24800 15568 24812
rect 15335 24772 15568 24800
rect 15335 24769 15347 24772
rect 15289 24763 15347 24769
rect 11057 24735 11115 24741
rect 11057 24732 11069 24735
rect 10980 24704 11069 24732
rect 11057 24701 11069 24704
rect 11103 24732 11115 24735
rect 12894 24732 12900 24744
rect 11103 24704 12900 24732
rect 11103 24701 11115 24704
rect 11057 24695 11115 24701
rect 12894 24692 12900 24704
rect 12952 24692 12958 24744
rect 12986 24692 12992 24744
rect 13044 24732 13050 24744
rect 13354 24732 13360 24744
rect 13044 24704 13360 24732
rect 13044 24692 13050 24704
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 13817 24735 13875 24741
rect 13817 24701 13829 24735
rect 13863 24732 13875 24735
rect 14476 24732 14504 24763
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 13863 24704 14504 24732
rect 14572 24735 14630 24741
rect 13863 24701 13875 24704
rect 13817 24695 13875 24701
rect 14572 24701 14584 24735
rect 14618 24732 14630 24735
rect 15378 24732 15384 24744
rect 14618 24704 15384 24732
rect 14618 24701 14630 24704
rect 14572 24695 14630 24701
rect 15378 24692 15384 24704
rect 15436 24692 15442 24744
rect 15473 24735 15531 24741
rect 15473 24701 15485 24735
rect 15519 24732 15531 24735
rect 15672 24732 15700 24840
rect 15930 24828 15936 24840
rect 15988 24828 15994 24880
rect 16114 24828 16120 24880
rect 16172 24877 16178 24880
rect 16172 24871 16207 24877
rect 16195 24837 16207 24871
rect 16172 24831 16207 24837
rect 16172 24828 16178 24831
rect 16574 24828 16580 24880
rect 16632 24868 16638 24880
rect 16945 24871 17003 24877
rect 16945 24868 16957 24871
rect 16632 24840 16957 24868
rect 16632 24828 16638 24840
rect 16945 24837 16957 24840
rect 16991 24868 17003 24871
rect 17770 24868 17776 24880
rect 16991 24840 17776 24868
rect 16991 24837 17003 24840
rect 16945 24831 17003 24837
rect 17770 24828 17776 24840
rect 17828 24828 17834 24880
rect 18782 24868 18788 24880
rect 17880 24840 18788 24868
rect 15948 24800 15976 24828
rect 16758 24800 16764 24812
rect 15948 24772 16764 24800
rect 16758 24760 16764 24772
rect 16816 24760 16822 24812
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24800 17187 24803
rect 17218 24800 17224 24812
rect 17175 24772 17224 24800
rect 17175 24769 17187 24772
rect 17129 24763 17187 24769
rect 17218 24760 17224 24772
rect 17276 24760 17282 24812
rect 15519 24704 15700 24732
rect 16776 24732 16804 24760
rect 17880 24741 17908 24840
rect 18782 24828 18788 24840
rect 18840 24828 18846 24880
rect 18892 24840 19196 24868
rect 17957 24803 18015 24809
rect 17957 24769 17969 24803
rect 18003 24800 18015 24803
rect 18046 24800 18052 24812
rect 18003 24772 18052 24800
rect 18003 24769 18015 24772
rect 17957 24763 18015 24769
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 18598 24800 18604 24812
rect 18196 24772 18604 24800
rect 18196 24760 18202 24772
rect 18598 24760 18604 24772
rect 18656 24800 18662 24812
rect 18892 24800 18920 24840
rect 18656 24772 18920 24800
rect 18656 24760 18662 24772
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19168 24809 19196 24840
rect 19242 24828 19248 24880
rect 19300 24868 19306 24880
rect 19300 24840 20024 24868
rect 19300 24828 19306 24840
rect 19153 24803 19211 24809
rect 19024 24772 19069 24800
rect 19024 24760 19030 24772
rect 19153 24769 19165 24803
rect 19199 24800 19211 24803
rect 19794 24800 19800 24812
rect 19199 24772 19800 24800
rect 19199 24769 19211 24772
rect 19153 24763 19211 24769
rect 19794 24760 19800 24772
rect 19852 24760 19858 24812
rect 19996 24809 20024 24840
rect 20070 24828 20076 24880
rect 20128 24868 20134 24880
rect 21192 24868 21220 24899
rect 21910 24896 21916 24908
rect 21968 24896 21974 24948
rect 22278 24896 22284 24948
rect 22336 24936 22342 24948
rect 24578 24936 24584 24948
rect 22336 24908 24584 24936
rect 22336 24896 22342 24908
rect 24578 24896 24584 24908
rect 24636 24896 24642 24948
rect 24946 24896 24952 24948
rect 25004 24936 25010 24948
rect 26510 24936 26516 24948
rect 25004 24908 26516 24936
rect 25004 24896 25010 24908
rect 26510 24896 26516 24908
rect 26568 24896 26574 24948
rect 26605 24939 26663 24945
rect 26605 24905 26617 24939
rect 26651 24936 26663 24939
rect 26694 24936 26700 24948
rect 26651 24908 26700 24936
rect 26651 24905 26663 24908
rect 26605 24899 26663 24905
rect 26694 24896 26700 24908
rect 26752 24896 26758 24948
rect 26903 24908 27568 24936
rect 20128 24840 21220 24868
rect 21361 24871 21419 24877
rect 20128 24828 20134 24840
rect 21361 24837 21373 24871
rect 21407 24868 21419 24871
rect 23566 24868 23572 24880
rect 21407 24840 23572 24868
rect 21407 24837 21419 24840
rect 21361 24831 21419 24837
rect 19981 24803 20039 24809
rect 19981 24769 19993 24803
rect 20027 24769 20039 24803
rect 21376 24800 21404 24831
rect 23566 24828 23572 24840
rect 23624 24828 23630 24880
rect 23842 24828 23848 24880
rect 23900 24868 23906 24880
rect 23900 24840 24058 24868
rect 23900 24828 23906 24840
rect 25038 24828 25044 24880
rect 25096 24868 25102 24880
rect 26786 24868 26792 24880
rect 25096 24840 26092 24868
rect 25096 24828 25102 24840
rect 22005 24803 22063 24809
rect 22005 24800 22017 24803
rect 19981 24763 20039 24769
rect 20067 24772 21404 24800
rect 21560 24772 22017 24800
rect 17865 24735 17923 24741
rect 16776 24704 17816 24732
rect 15519 24701 15531 24704
rect 15473 24695 15531 24701
rect 5994 24664 6000 24676
rect 5955 24636 6000 24664
rect 5994 24624 6000 24636
rect 6052 24624 6058 24676
rect 6733 24667 6791 24673
rect 6733 24633 6745 24667
rect 6779 24664 6791 24667
rect 8389 24667 8447 24673
rect 6779 24636 8340 24664
rect 6779 24633 6791 24636
rect 6733 24627 6791 24633
rect 7742 24596 7748 24608
rect 7703 24568 7748 24596
rect 7742 24556 7748 24568
rect 7800 24556 7806 24608
rect 8312 24596 8340 24636
rect 8389 24633 8401 24667
rect 8435 24664 8447 24667
rect 9766 24664 9772 24676
rect 8435 24636 9772 24664
rect 8435 24633 8447 24636
rect 8389 24627 8447 24633
rect 9766 24624 9772 24636
rect 9824 24664 9830 24676
rect 12529 24667 12587 24673
rect 12529 24664 12541 24667
rect 9824 24636 12541 24664
rect 9824 24624 9830 24636
rect 12529 24633 12541 24636
rect 12575 24664 12587 24667
rect 14734 24664 14740 24676
rect 12575 24636 14740 24664
rect 12575 24633 12587 24636
rect 12529 24627 12587 24633
rect 14734 24624 14740 24636
rect 14792 24624 14798 24676
rect 15930 24624 15936 24676
rect 15988 24664 15994 24676
rect 16301 24667 16359 24673
rect 16301 24664 16313 24667
rect 15988 24636 16313 24664
rect 15988 24624 15994 24636
rect 16301 24633 16313 24636
rect 16347 24633 16359 24667
rect 16301 24627 16359 24633
rect 16482 24624 16488 24676
rect 16540 24664 16546 24676
rect 17402 24664 17408 24676
rect 16540 24636 17408 24664
rect 16540 24624 16546 24636
rect 17402 24624 17408 24636
rect 17460 24624 17466 24676
rect 17788 24664 17816 24704
rect 17865 24701 17877 24735
rect 17911 24701 17923 24735
rect 18874 24732 18880 24744
rect 17865 24695 17923 24701
rect 17972 24704 18782 24732
rect 18835 24704 18880 24732
rect 17972 24664 18000 24704
rect 17788 24636 18000 24664
rect 18046 24624 18052 24676
rect 18104 24664 18110 24676
rect 18754 24664 18782 24704
rect 18874 24692 18880 24704
rect 18932 24692 18938 24744
rect 19061 24735 19119 24741
rect 19061 24701 19073 24735
rect 19107 24732 19119 24735
rect 19702 24732 19708 24744
rect 19107 24704 19708 24732
rect 19107 24701 19119 24704
rect 19061 24695 19119 24701
rect 19076 24664 19104 24695
rect 19702 24692 19708 24704
rect 19760 24692 19766 24744
rect 19889 24735 19947 24741
rect 19889 24732 19901 24735
rect 19805 24704 19901 24732
rect 18104 24636 18352 24664
rect 18754 24636 19104 24664
rect 18104 24624 18110 24636
rect 8478 24596 8484 24608
rect 8312 24568 8484 24596
rect 8478 24556 8484 24568
rect 8536 24556 8542 24608
rect 8938 24596 8944 24608
rect 8851 24568 8944 24596
rect 8938 24556 8944 24568
rect 8996 24596 9002 24608
rect 9674 24596 9680 24608
rect 8996 24568 9680 24596
rect 8996 24556 9002 24568
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 10226 24556 10232 24608
rect 10284 24596 10290 24608
rect 10597 24599 10655 24605
rect 10597 24596 10609 24599
rect 10284 24568 10609 24596
rect 10284 24556 10290 24568
rect 10597 24565 10609 24568
rect 10643 24596 10655 24599
rect 11054 24596 11060 24608
rect 10643 24568 11060 24596
rect 10643 24565 10655 24568
rect 10597 24559 10655 24565
rect 11054 24556 11060 24568
rect 11112 24556 11118 24608
rect 11882 24556 11888 24608
rect 11940 24596 11946 24608
rect 12250 24596 12256 24608
rect 11940 24568 12256 24596
rect 11940 24556 11946 24568
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 14458 24556 14464 24608
rect 14516 24596 14522 24608
rect 16022 24596 16028 24608
rect 14516 24568 16028 24596
rect 14516 24556 14522 24568
rect 16022 24556 16028 24568
rect 16080 24556 16086 24608
rect 16117 24599 16175 24605
rect 16117 24565 16129 24599
rect 16163 24596 16175 24599
rect 16850 24596 16856 24608
rect 16163 24568 16856 24596
rect 16163 24565 16175 24568
rect 16117 24559 16175 24565
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 17313 24599 17371 24605
rect 17313 24565 17325 24599
rect 17359 24596 17371 24599
rect 17586 24596 17592 24608
rect 17359 24568 17592 24596
rect 17359 24565 17371 24568
rect 17313 24559 17371 24565
rect 17586 24556 17592 24568
rect 17644 24556 17650 24608
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 18012 24568 18245 24596
rect 18012 24556 18018 24568
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 18324 24596 18352 24636
rect 19242 24624 19248 24676
rect 19300 24664 19306 24676
rect 19805 24664 19833 24704
rect 19889 24701 19901 24704
rect 19935 24701 19947 24735
rect 20067 24732 20095 24772
rect 21560 24744 21588 24772
rect 22005 24769 22017 24772
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 22152 24772 22201 24800
rect 22152 24760 22158 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 22281 24803 22339 24809
rect 22281 24769 22293 24803
rect 22327 24769 22339 24803
rect 22281 24763 22339 24769
rect 22373 24803 22431 24809
rect 22373 24769 22385 24803
rect 22419 24769 22431 24803
rect 25590 24800 25596 24812
rect 25551 24772 25596 24800
rect 22373 24763 22431 24769
rect 19889 24695 19947 24701
rect 19996 24704 20095 24732
rect 19996 24664 20024 24704
rect 20162 24692 20168 24744
rect 20220 24732 20226 24744
rect 20809 24735 20867 24741
rect 20809 24732 20821 24735
rect 20220 24704 20821 24732
rect 20220 24692 20226 24704
rect 20809 24701 20821 24704
rect 20855 24701 20867 24735
rect 20809 24695 20867 24701
rect 20993 24735 21051 24741
rect 20993 24701 21005 24735
rect 21039 24701 21051 24735
rect 20993 24695 21051 24701
rect 19300 24636 19833 24664
rect 19910 24636 20024 24664
rect 21008 24664 21036 24695
rect 21082 24692 21088 24744
rect 21140 24732 21146 24744
rect 21453 24735 21511 24741
rect 21140 24704 21185 24732
rect 21140 24692 21146 24704
rect 21453 24701 21465 24735
rect 21499 24701 21511 24735
rect 21453 24695 21511 24701
rect 21266 24664 21272 24676
rect 21008 24636 21272 24664
rect 19300 24624 19306 24636
rect 19150 24596 19156 24608
rect 18324 24568 19156 24596
rect 18233 24559 18291 24565
rect 19150 24556 19156 24568
rect 19208 24556 19214 24608
rect 19337 24599 19395 24605
rect 19337 24565 19349 24599
rect 19383 24596 19395 24599
rect 19702 24596 19708 24608
rect 19383 24568 19708 24596
rect 19383 24565 19395 24568
rect 19337 24559 19395 24565
rect 19702 24556 19708 24568
rect 19760 24556 19766 24608
rect 19794 24556 19800 24608
rect 19852 24596 19858 24608
rect 19910 24596 19938 24636
rect 21266 24624 21272 24636
rect 21324 24624 21330 24676
rect 21468 24664 21496 24695
rect 21542 24692 21548 24744
rect 21600 24692 21606 24744
rect 21818 24692 21824 24744
rect 21876 24732 21882 24744
rect 22296 24732 22324 24763
rect 21876 24704 22324 24732
rect 22388 24732 22416 24763
rect 25590 24760 25596 24772
rect 25648 24760 25654 24812
rect 25866 24800 25872 24812
rect 25827 24772 25872 24800
rect 25866 24760 25872 24772
rect 25924 24760 25930 24812
rect 25961 24803 26019 24809
rect 25961 24769 25973 24803
rect 26007 24769 26019 24803
rect 25961 24763 26019 24769
rect 23014 24732 23020 24744
rect 22388 24704 23020 24732
rect 21876 24692 21882 24704
rect 23014 24692 23020 24704
rect 23072 24692 23078 24744
rect 23106 24692 23112 24744
rect 23164 24732 23170 24744
rect 23293 24735 23351 24741
rect 23293 24732 23305 24735
rect 23164 24704 23305 24732
rect 23164 24692 23170 24704
rect 23293 24701 23305 24704
rect 23339 24701 23351 24735
rect 23569 24735 23627 24741
rect 23569 24732 23581 24735
rect 23293 24695 23351 24701
rect 23400 24704 23581 24732
rect 21468 24636 22784 24664
rect 19852 24568 19938 24596
rect 20257 24599 20315 24605
rect 19852 24556 19858 24568
rect 20257 24565 20269 24599
rect 20303 24596 20315 24599
rect 21818 24596 21824 24608
rect 20303 24568 21824 24596
rect 20303 24565 20315 24568
rect 20257 24559 20315 24565
rect 21818 24556 21824 24568
rect 21876 24596 21882 24608
rect 22462 24596 22468 24608
rect 21876 24568 22468 24596
rect 21876 24556 21882 24568
rect 22462 24556 22468 24568
rect 22520 24556 22526 24608
rect 22646 24596 22652 24608
rect 22607 24568 22652 24596
rect 22646 24556 22652 24568
rect 22704 24556 22710 24608
rect 22756 24596 22784 24636
rect 22922 24624 22928 24676
rect 22980 24664 22986 24676
rect 23400 24664 23428 24704
rect 23569 24701 23581 24704
rect 23615 24701 23627 24735
rect 23569 24695 23627 24701
rect 25038 24692 25044 24744
rect 25096 24732 25102 24744
rect 25976 24732 26004 24763
rect 25096 24704 26004 24732
rect 26064 24732 26092 24840
rect 26344 24840 26792 24868
rect 26344 24809 26372 24840
rect 26786 24828 26792 24840
rect 26844 24828 26850 24880
rect 26329 24803 26387 24809
rect 26329 24769 26341 24803
rect 26375 24800 26387 24803
rect 26510 24800 26516 24812
rect 26375 24772 26516 24800
rect 26375 24769 26387 24772
rect 26329 24763 26387 24769
rect 26510 24760 26516 24772
rect 26568 24760 26574 24812
rect 26605 24803 26663 24809
rect 26605 24769 26617 24803
rect 26651 24800 26663 24803
rect 26903 24800 26931 24908
rect 26970 24828 26976 24880
rect 27028 24868 27034 24880
rect 27222 24868 27228 24880
rect 27028 24840 27228 24868
rect 27028 24828 27034 24840
rect 27222 24828 27228 24840
rect 27280 24868 27286 24880
rect 27406 24871 27464 24877
rect 27406 24868 27418 24871
rect 27280 24840 27418 24868
rect 27280 24828 27286 24840
rect 27406 24837 27418 24840
rect 27452 24837 27464 24871
rect 27540 24868 27568 24908
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 28810 24936 28816 24948
rect 27672 24908 28816 24936
rect 27672 24896 27678 24908
rect 28810 24896 28816 24908
rect 28868 24896 28874 24948
rect 29086 24896 29092 24948
rect 29144 24936 29150 24948
rect 29733 24939 29791 24945
rect 29733 24936 29745 24939
rect 29144 24908 29745 24936
rect 29144 24896 29150 24908
rect 29733 24905 29745 24908
rect 29779 24936 29791 24939
rect 30834 24936 30840 24948
rect 29779 24908 30840 24936
rect 29779 24905 29791 24908
rect 29733 24899 29791 24905
rect 30834 24896 30840 24908
rect 30892 24896 30898 24948
rect 31110 24868 31116 24880
rect 27540 24840 31116 24868
rect 27406 24831 27464 24837
rect 31110 24828 31116 24840
rect 31168 24868 31174 24880
rect 31478 24868 31484 24880
rect 31168 24840 31484 24868
rect 31168 24828 31174 24840
rect 31478 24828 31484 24840
rect 31536 24828 31542 24880
rect 27062 24800 27068 24812
rect 26651 24772 27068 24800
rect 26651 24769 26663 24772
rect 26605 24763 26663 24769
rect 27062 24760 27068 24772
rect 27120 24760 27126 24812
rect 27310 24803 27368 24809
rect 27310 24769 27322 24803
rect 27356 24769 27368 24803
rect 27310 24763 27368 24769
rect 27325 24732 27353 24763
rect 27706 24760 27712 24812
rect 27764 24800 27770 24812
rect 27801 24803 27859 24809
rect 27801 24800 27813 24803
rect 27764 24772 27813 24800
rect 27764 24760 27770 24772
rect 27801 24769 27813 24772
rect 27847 24800 27859 24803
rect 28166 24800 28172 24812
rect 27847 24772 28172 24800
rect 27847 24769 27859 24772
rect 27801 24763 27859 24769
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 28442 24760 28448 24812
rect 28500 24800 28506 24812
rect 28537 24803 28595 24809
rect 28537 24800 28549 24803
rect 28500 24772 28549 24800
rect 28500 24760 28506 24772
rect 28537 24769 28549 24772
rect 28583 24769 28595 24803
rect 28537 24763 28595 24769
rect 28629 24803 28687 24809
rect 28629 24769 28641 24803
rect 28675 24769 28687 24803
rect 28629 24763 28687 24769
rect 26064 24704 27910 24732
rect 25096 24692 25102 24704
rect 22980 24636 23428 24664
rect 22980 24624 22986 24636
rect 24670 24624 24676 24676
rect 24728 24664 24734 24676
rect 27882 24664 27910 24704
rect 27982 24692 27988 24744
rect 28040 24732 28046 24744
rect 28644 24732 28672 24763
rect 28718 24760 28724 24812
rect 28776 24800 28782 24812
rect 28905 24803 28963 24809
rect 28776 24772 28821 24800
rect 28776 24760 28782 24772
rect 28905 24769 28917 24803
rect 28951 24800 28963 24803
rect 29270 24800 29276 24812
rect 28951 24772 29276 24800
rect 28951 24769 28963 24772
rect 28905 24763 28963 24769
rect 29270 24760 29276 24772
rect 29328 24760 29334 24812
rect 29641 24803 29699 24809
rect 29641 24769 29653 24803
rect 29687 24800 29699 24803
rect 29730 24800 29736 24812
rect 29687 24772 29736 24800
rect 29687 24769 29699 24772
rect 29641 24763 29699 24769
rect 29730 24760 29736 24772
rect 29788 24760 29794 24812
rect 29822 24760 29828 24812
rect 29880 24809 29886 24812
rect 29880 24803 29908 24809
rect 29896 24769 29908 24803
rect 29880 24763 29908 24769
rect 29880 24760 29886 24763
rect 30374 24760 30380 24812
rect 30432 24800 30438 24812
rect 30469 24803 30527 24809
rect 30469 24800 30481 24803
rect 30432 24772 30481 24800
rect 30432 24760 30438 24772
rect 30469 24769 30481 24772
rect 30515 24769 30527 24803
rect 30469 24763 30527 24769
rect 30653 24803 30711 24809
rect 30653 24769 30665 24803
rect 30699 24769 30711 24803
rect 30653 24763 30711 24769
rect 28040 24704 28672 24732
rect 29365 24735 29423 24741
rect 28040 24692 28046 24704
rect 29365 24701 29377 24735
rect 29411 24732 29423 24735
rect 30006 24732 30012 24744
rect 29411 24704 30012 24732
rect 29411 24701 29423 24704
rect 29365 24695 29423 24701
rect 30006 24692 30012 24704
rect 30064 24692 30070 24744
rect 30668 24732 30696 24763
rect 30742 24760 30748 24812
rect 30800 24800 30806 24812
rect 30800 24772 30845 24800
rect 30800 24760 30806 24772
rect 30926 24760 30932 24812
rect 30984 24800 30990 24812
rect 32214 24800 32220 24812
rect 30984 24772 32220 24800
rect 30984 24760 30990 24772
rect 32214 24760 32220 24772
rect 32272 24760 32278 24812
rect 32490 24732 32496 24744
rect 30668 24704 32496 24732
rect 29730 24664 29736 24676
rect 24728 24636 27844 24664
rect 27882 24636 29736 24664
rect 24728 24624 24734 24636
rect 24302 24596 24308 24608
rect 22756 24568 24308 24596
rect 24302 24556 24308 24568
rect 24360 24556 24366 24608
rect 25038 24596 25044 24608
rect 24999 24568 25044 24596
rect 25038 24556 25044 24568
rect 25096 24556 25102 24608
rect 25774 24556 25780 24608
rect 25832 24596 25838 24608
rect 27157 24599 27215 24605
rect 27157 24596 27169 24599
rect 25832 24568 27169 24596
rect 25832 24556 25838 24568
rect 27157 24565 27169 24568
rect 27203 24565 27215 24599
rect 27157 24559 27215 24565
rect 27246 24556 27252 24608
rect 27304 24596 27310 24608
rect 27522 24596 27528 24608
rect 27304 24568 27528 24596
rect 27304 24556 27310 24568
rect 27522 24556 27528 24568
rect 27580 24556 27586 24608
rect 27706 24596 27712 24608
rect 27667 24568 27712 24596
rect 27706 24556 27712 24568
rect 27764 24556 27770 24608
rect 27816 24596 27844 24636
rect 29730 24624 29736 24636
rect 29788 24664 29794 24676
rect 30668 24664 30696 24704
rect 32490 24692 32496 24704
rect 32548 24692 32554 24744
rect 30834 24664 30840 24676
rect 29788 24636 30696 24664
rect 30795 24636 30840 24664
rect 29788 24624 29794 24636
rect 30834 24624 30840 24636
rect 30892 24624 30898 24676
rect 28261 24599 28319 24605
rect 28261 24596 28273 24599
rect 27816 24568 28273 24596
rect 28261 24565 28273 24568
rect 28307 24565 28319 24599
rect 28261 24559 28319 24565
rect 28442 24556 28448 24608
rect 28500 24596 28506 24608
rect 29270 24596 29276 24608
rect 28500 24568 29276 24596
rect 28500 24556 28506 24568
rect 29270 24556 29276 24568
rect 29328 24556 29334 24608
rect 30009 24599 30067 24605
rect 30009 24565 30021 24599
rect 30055 24596 30067 24599
rect 32582 24596 32588 24608
rect 30055 24568 32588 24596
rect 30055 24565 30067 24568
rect 30009 24559 30067 24565
rect 32582 24556 32588 24568
rect 32640 24556 32646 24608
rect 1104 24506 31832 24528
rect 1104 24454 4791 24506
rect 4843 24454 4855 24506
rect 4907 24454 4919 24506
rect 4971 24454 4983 24506
rect 5035 24454 5047 24506
rect 5099 24454 12473 24506
rect 12525 24454 12537 24506
rect 12589 24454 12601 24506
rect 12653 24454 12665 24506
rect 12717 24454 12729 24506
rect 12781 24454 20155 24506
rect 20207 24454 20219 24506
rect 20271 24454 20283 24506
rect 20335 24454 20347 24506
rect 20399 24454 20411 24506
rect 20463 24454 27837 24506
rect 27889 24454 27901 24506
rect 27953 24454 27965 24506
rect 28017 24454 28029 24506
rect 28081 24454 28093 24506
rect 28145 24454 31832 24506
rect 1104 24432 31832 24454
rect 4154 24392 4160 24404
rect 4115 24364 4160 24392
rect 4154 24352 4160 24364
rect 4212 24352 4218 24404
rect 6914 24352 6920 24404
rect 6972 24392 6978 24404
rect 7929 24395 7987 24401
rect 7929 24392 7941 24395
rect 6972 24364 7941 24392
rect 6972 24352 6978 24364
rect 7929 24361 7941 24364
rect 7975 24361 7987 24395
rect 7929 24355 7987 24361
rect 8478 24352 8484 24404
rect 8536 24392 8542 24404
rect 10226 24392 10232 24404
rect 8536 24364 10232 24392
rect 8536 24352 8542 24364
rect 10226 24352 10232 24364
rect 10284 24352 10290 24404
rect 11790 24352 11796 24404
rect 11848 24392 11854 24404
rect 11848 24364 14688 24392
rect 11848 24352 11854 24364
rect 5810 24324 5816 24336
rect 5723 24296 5816 24324
rect 5810 24284 5816 24296
rect 5868 24324 5874 24336
rect 12897 24327 12955 24333
rect 5868 24296 12848 24324
rect 5868 24284 5874 24296
rect 5261 24259 5319 24265
rect 5261 24225 5273 24259
rect 5307 24256 5319 24259
rect 8938 24256 8944 24268
rect 5307 24228 8944 24256
rect 5307 24225 5319 24228
rect 5261 24219 5319 24225
rect 8938 24216 8944 24228
rect 8996 24216 9002 24268
rect 9582 24216 9588 24268
rect 9640 24216 9646 24268
rect 9674 24216 9680 24268
rect 9732 24256 9738 24268
rect 10226 24256 10232 24268
rect 9732 24228 10232 24256
rect 9732 24216 9738 24228
rect 10226 24216 10232 24228
rect 10284 24256 10290 24268
rect 10284 24228 11744 24256
rect 10284 24216 10290 24228
rect 9600 24188 9628 24216
rect 11716 24200 11744 24228
rect 11882 24216 11888 24268
rect 11940 24256 11946 24268
rect 12345 24259 12403 24265
rect 12345 24256 12357 24259
rect 11940 24228 12357 24256
rect 11940 24216 11946 24228
rect 12345 24225 12357 24228
rect 12391 24256 12403 24259
rect 12820 24256 12848 24296
rect 12897 24293 12909 24327
rect 12943 24324 12955 24327
rect 13538 24324 13544 24336
rect 12943 24296 13544 24324
rect 12943 24293 12955 24296
rect 12897 24287 12955 24293
rect 13538 24284 13544 24296
rect 13596 24284 13602 24336
rect 13906 24284 13912 24336
rect 13964 24284 13970 24336
rect 14660 24324 14688 24364
rect 14734 24352 14740 24404
rect 14792 24392 14798 24404
rect 14792 24364 14837 24392
rect 14792 24352 14798 24364
rect 15010 24352 15016 24404
rect 15068 24392 15074 24404
rect 15105 24395 15163 24401
rect 15105 24392 15117 24395
rect 15068 24364 15117 24392
rect 15068 24352 15074 24364
rect 15105 24361 15117 24364
rect 15151 24361 15163 24395
rect 15746 24392 15752 24404
rect 15105 24355 15163 24361
rect 15196 24364 15752 24392
rect 15196 24324 15224 24364
rect 15746 24352 15752 24364
rect 15804 24352 15810 24404
rect 15930 24352 15936 24404
rect 15988 24392 15994 24404
rect 18325 24395 18383 24401
rect 15988 24364 18091 24392
rect 15988 24352 15994 24364
rect 14660 24296 15224 24324
rect 16206 24284 16212 24336
rect 16264 24324 16270 24336
rect 16485 24327 16543 24333
rect 16485 24324 16497 24327
rect 16264 24296 16497 24324
rect 16264 24284 16270 24296
rect 16485 24293 16497 24296
rect 16531 24293 16543 24327
rect 16485 24287 16543 24293
rect 16853 24327 16911 24333
rect 16853 24293 16865 24327
rect 16899 24324 16911 24327
rect 18063 24324 18091 24364
rect 18325 24361 18337 24395
rect 18371 24392 18383 24395
rect 18414 24392 18420 24404
rect 18371 24364 18420 24392
rect 18371 24361 18383 24364
rect 18325 24355 18383 24361
rect 18414 24352 18420 24364
rect 18472 24352 18478 24404
rect 20346 24392 20352 24404
rect 18524 24364 20352 24392
rect 18524 24324 18552 24364
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 21450 24392 21456 24404
rect 20548 24364 21456 24392
rect 18690 24324 18696 24336
rect 16899 24296 18000 24324
rect 18063 24296 18552 24324
rect 18651 24296 18696 24324
rect 16899 24293 16911 24296
rect 16853 24287 16911 24293
rect 13722 24256 13728 24268
rect 12391 24228 12674 24256
rect 12820 24228 13032 24256
rect 12391 24225 12403 24228
rect 12345 24219 12403 24225
rect 10134 24188 10140 24200
rect 6288 24160 9628 24188
rect 10095 24160 10140 24188
rect 4709 24123 4767 24129
rect 4709 24089 4721 24123
rect 4755 24120 4767 24123
rect 5902 24120 5908 24132
rect 4755 24092 5908 24120
rect 4755 24089 4767 24092
rect 4709 24083 4767 24089
rect 5902 24080 5908 24092
rect 5960 24080 5966 24132
rect 5626 24012 5632 24064
rect 5684 24052 5690 24064
rect 6288 24061 6316 24160
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 11698 24148 11704 24200
rect 11756 24188 11762 24200
rect 12253 24191 12311 24197
rect 12253 24188 12265 24191
rect 11756 24160 12265 24188
rect 11756 24148 11762 24160
rect 12253 24157 12265 24160
rect 12299 24157 12311 24191
rect 12253 24151 12311 24157
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 12646 24188 12674 24228
rect 12897 24191 12955 24197
rect 12897 24188 12909 24191
rect 12492 24160 12537 24188
rect 12646 24160 12909 24188
rect 12492 24148 12498 24160
rect 12897 24157 12909 24160
rect 12943 24157 12955 24191
rect 12897 24151 12955 24157
rect 6914 24120 6920 24132
rect 6875 24092 6920 24120
rect 6914 24080 6920 24092
rect 6972 24080 6978 24132
rect 7650 24080 7656 24132
rect 7708 24120 7714 24132
rect 8478 24120 8484 24132
rect 7708 24092 8484 24120
rect 7708 24080 7714 24092
rect 8478 24080 8484 24092
rect 8536 24080 8542 24132
rect 9582 24080 9588 24132
rect 9640 24120 9646 24132
rect 13004 24120 13032 24228
rect 13096 24228 13728 24256
rect 13096 24197 13124 24228
rect 13722 24216 13728 24228
rect 13780 24216 13786 24268
rect 13924 24256 13952 24284
rect 16390 24256 16396 24268
rect 13924 24228 14780 24256
rect 16351 24228 16396 24256
rect 13081 24191 13139 24197
rect 13081 24157 13093 24191
rect 13127 24157 13139 24191
rect 13081 24151 13139 24157
rect 13354 24148 13360 24200
rect 13412 24188 13418 24200
rect 13541 24191 13599 24197
rect 13541 24188 13553 24191
rect 13412 24160 13553 24188
rect 13412 24148 13418 24160
rect 13541 24157 13553 24160
rect 13587 24188 13599 24191
rect 13906 24188 13912 24200
rect 13587 24160 13912 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14752 24197 14780 24228
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 16758 24216 16764 24268
rect 16816 24256 16822 24268
rect 17589 24259 17647 24265
rect 17589 24256 17601 24259
rect 16816 24228 17601 24256
rect 16816 24216 16822 24228
rect 17589 24225 17601 24228
rect 17635 24225 17647 24259
rect 17972 24256 18000 24296
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 19150 24284 19156 24336
rect 19208 24324 19214 24336
rect 20548 24324 20576 24364
rect 21450 24352 21456 24364
rect 21508 24352 21514 24404
rect 21563 24395 21621 24401
rect 21563 24361 21575 24395
rect 21609 24392 21621 24395
rect 21726 24392 21732 24404
rect 21609 24364 21732 24392
rect 21609 24361 21621 24364
rect 21563 24355 21621 24361
rect 21726 24352 21732 24364
rect 21784 24352 21790 24404
rect 22922 24392 22928 24404
rect 21836 24364 22928 24392
rect 21836 24336 21864 24364
rect 22922 24352 22928 24364
rect 22980 24352 22986 24404
rect 24029 24395 24087 24401
rect 24029 24361 24041 24395
rect 24075 24392 24087 24395
rect 24394 24392 24400 24404
rect 24075 24364 24400 24392
rect 24075 24361 24087 24364
rect 24029 24355 24087 24361
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 25038 24352 25044 24404
rect 25096 24392 25102 24404
rect 26694 24392 26700 24404
rect 25096 24364 26700 24392
rect 25096 24352 25102 24364
rect 26694 24352 26700 24364
rect 26752 24352 26758 24404
rect 27614 24392 27620 24404
rect 26988 24364 27620 24392
rect 19208 24296 20576 24324
rect 19208 24284 19214 24296
rect 21818 24284 21824 24336
rect 21876 24284 21882 24336
rect 22066 24296 22416 24324
rect 22066 24256 22094 24296
rect 22278 24256 22284 24268
rect 17589 24219 17647 24225
rect 17696 24228 17908 24256
rect 17972 24228 22094 24256
rect 22239 24228 22284 24256
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24157 14887 24191
rect 14829 24151 14887 24157
rect 14936 24160 15700 24188
rect 13998 24120 14004 24132
rect 9640 24092 12940 24120
rect 13004 24092 14004 24120
rect 9640 24080 9646 24092
rect 6273 24055 6331 24061
rect 6273 24052 6285 24055
rect 5684 24024 6285 24052
rect 5684 24012 5690 24024
rect 6273 24021 6285 24024
rect 6319 24021 6331 24055
rect 6273 24015 6331 24021
rect 7469 24055 7527 24061
rect 7469 24021 7481 24055
rect 7515 24052 7527 24055
rect 7742 24052 7748 24064
rect 7515 24024 7748 24052
rect 7515 24021 7527 24024
rect 7469 24015 7527 24021
rect 7742 24012 7748 24024
rect 7800 24012 7806 24064
rect 9398 24012 9404 24064
rect 9456 24052 9462 24064
rect 9493 24055 9551 24061
rect 9493 24052 9505 24055
rect 9456 24024 9505 24052
rect 9456 24012 9462 24024
rect 9493 24021 9505 24024
rect 9539 24021 9551 24055
rect 9493 24015 9551 24021
rect 10689 24055 10747 24061
rect 10689 24021 10701 24055
rect 10735 24052 10747 24055
rect 10962 24052 10968 24064
rect 10735 24024 10968 24052
rect 10735 24021 10747 24024
rect 10689 24015 10747 24021
rect 10962 24012 10968 24024
rect 11020 24012 11026 24064
rect 11241 24055 11299 24061
rect 11241 24021 11253 24055
rect 11287 24052 11299 24055
rect 11793 24055 11851 24061
rect 11793 24052 11805 24055
rect 11287 24024 11805 24052
rect 11287 24021 11299 24024
rect 11241 24015 11299 24021
rect 11793 24021 11805 24024
rect 11839 24052 11851 24055
rect 12250 24052 12256 24064
rect 11839 24024 12256 24052
rect 11839 24021 11851 24024
rect 11793 24015 11851 24021
rect 12250 24012 12256 24024
rect 12308 24012 12314 24064
rect 12912 24052 12940 24092
rect 13998 24080 14004 24092
rect 14056 24120 14062 24132
rect 14274 24120 14280 24132
rect 14056 24092 14280 24120
rect 14056 24080 14062 24092
rect 14274 24080 14280 24092
rect 14332 24080 14338 24132
rect 14366 24080 14372 24132
rect 14424 24120 14430 24132
rect 14844 24120 14872 24151
rect 14424 24092 14872 24120
rect 14424 24080 14430 24092
rect 13354 24052 13360 24064
rect 12912 24024 13360 24052
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 13633 24055 13691 24061
rect 13633 24021 13645 24055
rect 13679 24052 13691 24055
rect 13906 24052 13912 24064
rect 13679 24024 13912 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 14090 24012 14096 24064
rect 14148 24052 14154 24064
rect 14936 24052 14964 24160
rect 15672 24132 15700 24160
rect 16298 24148 16304 24200
rect 16356 24188 16362 24200
rect 16669 24191 16727 24197
rect 16669 24188 16681 24191
rect 16356 24160 16681 24188
rect 16356 24148 16362 24160
rect 16669 24157 16681 24160
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 16850 24148 16856 24200
rect 16908 24188 16914 24200
rect 17310 24188 17316 24200
rect 16908 24160 17316 24188
rect 16908 24148 16914 24160
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 17494 24188 17500 24200
rect 17455 24160 17500 24188
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 17696 24197 17724 24228
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 15562 24120 15568 24132
rect 15523 24092 15568 24120
rect 15562 24080 15568 24092
rect 15620 24080 15626 24132
rect 15654 24080 15660 24132
rect 15712 24120 15718 24132
rect 15765 24123 15823 24129
rect 15765 24120 15777 24123
rect 15712 24092 15777 24120
rect 15712 24080 15718 24092
rect 15765 24089 15777 24092
rect 15811 24089 15823 24123
rect 15765 24083 15823 24089
rect 16942 24080 16948 24132
rect 17000 24120 17006 24132
rect 17696 24120 17724 24151
rect 17000 24092 17724 24120
rect 17000 24080 17006 24092
rect 14148 24024 14964 24052
rect 14148 24012 14154 24024
rect 15010 24012 15016 24064
rect 15068 24052 15074 24064
rect 15933 24055 15991 24061
rect 15933 24052 15945 24055
rect 15068 24024 15945 24052
rect 15068 24012 15074 24024
rect 15933 24021 15945 24024
rect 15979 24021 15991 24055
rect 15933 24015 15991 24021
rect 16666 24012 16672 24064
rect 16724 24052 16730 24064
rect 17313 24055 17371 24061
rect 17313 24052 17325 24055
rect 16724 24024 17325 24052
rect 16724 24012 16730 24024
rect 17313 24021 17325 24024
rect 17359 24021 17371 24055
rect 17313 24015 17371 24021
rect 17402 24012 17408 24064
rect 17460 24052 17466 24064
rect 17788 24052 17816 24151
rect 17880 24120 17908 24228
rect 22278 24216 22284 24228
rect 22336 24216 22342 24268
rect 22388 24256 22416 24296
rect 23566 24284 23572 24336
rect 23624 24324 23630 24336
rect 24486 24324 24492 24336
rect 23624 24296 24492 24324
rect 23624 24284 23630 24296
rect 24486 24284 24492 24296
rect 24544 24284 24550 24336
rect 25866 24284 25872 24336
rect 25924 24324 25930 24336
rect 26329 24327 26387 24333
rect 26329 24324 26341 24327
rect 25924 24296 26341 24324
rect 25924 24284 25930 24296
rect 26329 24293 26341 24296
rect 26375 24324 26387 24327
rect 26988 24324 27016 24364
rect 27614 24352 27620 24364
rect 27672 24352 27678 24404
rect 28258 24352 28264 24404
rect 28316 24392 28322 24404
rect 28629 24395 28687 24401
rect 28629 24392 28641 24395
rect 28316 24364 28641 24392
rect 28316 24352 28322 24364
rect 28629 24361 28641 24364
rect 28675 24361 28687 24395
rect 28629 24355 28687 24361
rect 26375 24296 27016 24324
rect 28644 24324 28672 24355
rect 28902 24352 28908 24404
rect 28960 24392 28966 24404
rect 30377 24395 30435 24401
rect 30377 24392 30389 24395
rect 28960 24364 30389 24392
rect 28960 24352 28966 24364
rect 30377 24361 30389 24364
rect 30423 24361 30435 24395
rect 31018 24392 31024 24404
rect 30979 24364 31024 24392
rect 30377 24355 30435 24361
rect 31018 24352 31024 24364
rect 31076 24352 31082 24404
rect 29178 24324 29184 24336
rect 28644 24296 28948 24324
rect 29091 24296 29184 24324
rect 26375 24293 26387 24296
rect 26329 24287 26387 24293
rect 28920 24268 28948 24296
rect 29178 24284 29184 24296
rect 29236 24324 29242 24336
rect 29914 24324 29920 24336
rect 29236 24296 29920 24324
rect 29236 24284 29242 24296
rect 29914 24284 29920 24296
rect 29972 24324 29978 24336
rect 31202 24324 31208 24336
rect 29972 24296 31208 24324
rect 29972 24284 29978 24296
rect 31202 24284 31208 24296
rect 31260 24284 31266 24336
rect 22557 24259 22615 24265
rect 22557 24256 22569 24259
rect 22388 24228 22569 24256
rect 22557 24225 22569 24228
rect 22603 24225 22615 24259
rect 22557 24219 22615 24225
rect 22922 24216 22928 24268
rect 22980 24256 22986 24268
rect 24857 24259 24915 24265
rect 24857 24256 24869 24259
rect 22980 24228 24869 24256
rect 22980 24216 22986 24228
rect 24857 24225 24869 24228
rect 24903 24225 24915 24259
rect 24857 24219 24915 24225
rect 25406 24216 25412 24268
rect 25464 24256 25470 24268
rect 28718 24256 28724 24268
rect 25464 24228 28724 24256
rect 25464 24216 25470 24228
rect 28718 24216 28724 24228
rect 28776 24216 28782 24268
rect 28902 24216 28908 24268
rect 28960 24216 28966 24268
rect 29638 24216 29644 24268
rect 29696 24256 29702 24268
rect 31018 24256 31024 24268
rect 29696 24228 30144 24256
rect 30979 24228 31024 24256
rect 29696 24216 29702 24228
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 18138 24188 18144 24200
rect 18012 24160 18144 24188
rect 18012 24148 18018 24160
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18322 24148 18328 24200
rect 18380 24188 18386 24200
rect 18509 24191 18567 24197
rect 18509 24188 18521 24191
rect 18380 24160 18521 24188
rect 18380 24148 18386 24160
rect 18509 24157 18521 24160
rect 18555 24157 18567 24191
rect 18509 24151 18567 24157
rect 18598 24148 18604 24200
rect 18656 24188 18662 24200
rect 18785 24191 18843 24197
rect 18656 24160 18701 24188
rect 18656 24148 18662 24160
rect 18785 24157 18797 24191
rect 18831 24188 18843 24191
rect 18874 24188 18880 24200
rect 18831 24160 18880 24188
rect 18831 24157 18843 24160
rect 18785 24151 18843 24157
rect 18874 24148 18880 24160
rect 18932 24148 18938 24200
rect 18966 24148 18972 24200
rect 19024 24188 19030 24200
rect 19334 24188 19340 24200
rect 19024 24160 19340 24188
rect 19024 24148 19030 24160
rect 19334 24148 19340 24160
rect 19392 24148 19398 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19518 24188 19524 24200
rect 19475 24160 19524 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 19978 24188 19984 24200
rect 19659 24160 19984 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 19978 24148 19984 24160
rect 20036 24148 20042 24200
rect 20070 24148 20076 24200
rect 20128 24188 20134 24200
rect 20254 24188 20260 24200
rect 20128 24160 20260 24188
rect 20128 24148 20134 24160
rect 20254 24148 20260 24160
rect 20312 24148 20318 24200
rect 21821 24191 21879 24197
rect 21821 24157 21833 24191
rect 21867 24188 21879 24191
rect 22094 24188 22100 24200
rect 21867 24160 22100 24188
rect 21867 24157 21879 24160
rect 21821 24151 21879 24157
rect 22094 24148 22100 24160
rect 22152 24148 22158 24200
rect 23658 24148 23664 24200
rect 23716 24148 23722 24200
rect 24578 24188 24584 24200
rect 24491 24160 24584 24188
rect 24578 24148 24584 24160
rect 24636 24148 24642 24200
rect 25958 24148 25964 24200
rect 26016 24148 26022 24200
rect 26881 24191 26939 24197
rect 26881 24188 26893 24191
rect 26159 24160 26893 24188
rect 17880 24092 20116 24120
rect 17460 24024 17816 24052
rect 17460 24012 17466 24024
rect 17862 24012 17868 24064
rect 17920 24052 17926 24064
rect 19242 24052 19248 24064
rect 17920 24024 19248 24052
rect 17920 24012 17926 24024
rect 19242 24012 19248 24024
rect 19300 24012 19306 24064
rect 19334 24012 19340 24064
rect 19392 24052 19398 24064
rect 19429 24055 19487 24061
rect 19429 24052 19441 24055
rect 19392 24024 19441 24052
rect 19392 24012 19398 24024
rect 19429 24021 19441 24024
rect 19475 24021 19487 24055
rect 19429 24015 19487 24021
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 19886 24052 19892 24064
rect 19760 24024 19892 24052
rect 19760 24012 19766 24024
rect 19886 24012 19892 24024
rect 19944 24012 19950 24064
rect 20088 24061 20116 24092
rect 21082 24080 21088 24132
rect 21140 24080 21146 24132
rect 21266 24080 21272 24132
rect 21324 24120 21330 24132
rect 22830 24120 22836 24132
rect 21324 24092 22836 24120
rect 21324 24080 21330 24092
rect 22830 24080 22836 24092
rect 22888 24080 22894 24132
rect 24596 24120 24624 24148
rect 24596 24092 25084 24120
rect 25056 24064 25084 24092
rect 20073 24055 20131 24061
rect 20073 24021 20085 24055
rect 20119 24052 20131 24055
rect 23566 24052 23572 24064
rect 20119 24024 23572 24052
rect 20119 24021 20131 24024
rect 20073 24015 20131 24021
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 25038 24012 25044 24064
rect 25096 24052 25102 24064
rect 26159 24052 26187 24160
rect 26881 24157 26893 24160
rect 26927 24157 26939 24191
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 26881 24151 26939 24157
rect 28644 24160 29745 24188
rect 27157 24123 27215 24129
rect 27157 24089 27169 24123
rect 27203 24089 27215 24123
rect 28534 24120 28540 24132
rect 28382 24092 28540 24120
rect 27157 24083 27215 24089
rect 25096 24024 26187 24052
rect 25096 24012 25102 24024
rect 26234 24012 26240 24064
rect 26292 24052 26298 24064
rect 27172 24052 27200 24083
rect 28534 24080 28540 24092
rect 28592 24080 28598 24132
rect 26292 24024 27200 24052
rect 26292 24012 26298 24024
rect 27798 24012 27804 24064
rect 27856 24052 27862 24064
rect 28644 24052 28672 24160
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 29822 24148 29828 24200
rect 29880 24188 29886 24200
rect 30116 24197 30144 24228
rect 31018 24216 31024 24228
rect 31076 24216 31082 24268
rect 29917 24191 29975 24197
rect 29917 24188 29929 24191
rect 29880 24160 29929 24188
rect 29880 24148 29886 24160
rect 29917 24157 29929 24160
rect 29963 24157 29975 24191
rect 29917 24151 29975 24157
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 30101 24191 30159 24197
rect 30101 24157 30113 24191
rect 30147 24157 30159 24191
rect 30101 24151 30159 24157
rect 29178 24080 29184 24132
rect 29236 24120 29242 24132
rect 29454 24120 29460 24132
rect 29236 24092 29460 24120
rect 29236 24080 29242 24092
rect 29454 24080 29460 24092
rect 29512 24080 29518 24132
rect 30024 24120 30052 24151
rect 30742 24148 30748 24200
rect 30800 24188 30806 24200
rect 31113 24191 31171 24197
rect 31113 24188 31125 24191
rect 30800 24160 31125 24188
rect 30800 24148 30806 24160
rect 31113 24157 31125 24160
rect 31159 24157 31171 24191
rect 31113 24151 31171 24157
rect 30834 24120 30840 24132
rect 29840 24092 30052 24120
rect 30795 24092 30840 24120
rect 29840 24064 29868 24092
rect 30834 24080 30840 24092
rect 30892 24080 30898 24132
rect 27856 24024 28672 24052
rect 27856 24012 27862 24024
rect 28718 24012 28724 24064
rect 28776 24052 28782 24064
rect 29730 24052 29736 24064
rect 28776 24024 29736 24052
rect 28776 24012 28782 24024
rect 29730 24012 29736 24024
rect 29788 24012 29794 24064
rect 29822 24012 29828 24064
rect 29880 24012 29886 24064
rect 31297 24055 31355 24061
rect 31297 24021 31309 24055
rect 31343 24052 31355 24055
rect 31570 24052 31576 24064
rect 31343 24024 31576 24052
rect 31343 24021 31355 24024
rect 31297 24015 31355 24021
rect 31570 24012 31576 24024
rect 31628 24012 31634 24064
rect 1104 23962 31992 23984
rect 1104 23910 8632 23962
rect 8684 23910 8696 23962
rect 8748 23910 8760 23962
rect 8812 23910 8824 23962
rect 8876 23910 8888 23962
rect 8940 23910 16314 23962
rect 16366 23910 16378 23962
rect 16430 23910 16442 23962
rect 16494 23910 16506 23962
rect 16558 23910 16570 23962
rect 16622 23910 23996 23962
rect 24048 23910 24060 23962
rect 24112 23910 24124 23962
rect 24176 23910 24188 23962
rect 24240 23910 24252 23962
rect 24304 23910 31678 23962
rect 31730 23910 31742 23962
rect 31794 23910 31806 23962
rect 31858 23910 31870 23962
rect 31922 23910 31934 23962
rect 31986 23910 31992 23962
rect 1104 23888 31992 23910
rect 4338 23848 4344 23860
rect 4299 23820 4344 23848
rect 4338 23808 4344 23820
rect 4396 23808 4402 23860
rect 7006 23808 7012 23860
rect 7064 23848 7070 23860
rect 7282 23848 7288 23860
rect 7064 23820 7288 23848
rect 7064 23808 7070 23820
rect 7282 23808 7288 23820
rect 7340 23848 7346 23860
rect 9398 23848 9404 23860
rect 7340 23820 9404 23848
rect 7340 23808 7346 23820
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 9493 23851 9551 23857
rect 9493 23817 9505 23851
rect 9539 23848 9551 23851
rect 10870 23848 10876 23860
rect 9539 23820 10876 23848
rect 9539 23817 9551 23820
rect 9493 23811 9551 23817
rect 10870 23808 10876 23820
rect 10928 23848 10934 23860
rect 12158 23848 12164 23860
rect 10928 23820 12020 23848
rect 12119 23820 12164 23848
rect 10928 23808 10934 23820
rect 6733 23783 6791 23789
rect 6733 23749 6745 23783
rect 6779 23780 6791 23783
rect 10502 23780 10508 23792
rect 6779 23752 10508 23780
rect 6779 23749 6791 23752
rect 6733 23743 6791 23749
rect 10502 23740 10508 23752
rect 10560 23740 10566 23792
rect 11146 23740 11152 23792
rect 11204 23780 11210 23792
rect 11992 23780 12020 23820
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 14385 23851 14443 23857
rect 14385 23848 14397 23851
rect 12360 23820 14397 23848
rect 12360 23780 12388 23820
rect 14385 23817 14397 23820
rect 14431 23817 14443 23851
rect 15378 23848 15384 23860
rect 15339 23820 15384 23848
rect 14385 23811 14443 23817
rect 15378 23808 15384 23820
rect 15436 23808 15442 23860
rect 15470 23808 15476 23860
rect 15528 23848 15534 23860
rect 20622 23848 20628 23860
rect 15528 23820 18368 23848
rect 15528 23808 15534 23820
rect 18340 23792 18368 23820
rect 19444 23820 20628 23848
rect 14090 23780 14096 23792
rect 11204 23752 11560 23780
rect 11992 23752 12388 23780
rect 12728 23752 14096 23780
rect 11204 23740 11210 23752
rect 4893 23715 4951 23721
rect 4893 23681 4905 23715
rect 4939 23712 4951 23715
rect 10410 23712 10416 23724
rect 4939 23684 10416 23712
rect 4939 23681 4951 23684
rect 4893 23675 4951 23681
rect 10410 23672 10416 23684
rect 10468 23672 10474 23724
rect 11054 23672 11060 23724
rect 11112 23712 11118 23724
rect 11422 23712 11428 23724
rect 11112 23684 11428 23712
rect 11112 23672 11118 23684
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11532 23712 11560 23752
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 11532 23684 12173 23712
rect 12161 23681 12173 23684
rect 12207 23681 12219 23715
rect 12342 23712 12348 23724
rect 12303 23684 12348 23712
rect 12161 23675 12219 23681
rect 12342 23672 12348 23684
rect 12400 23672 12406 23724
rect 1578 23644 1584 23656
rect 1539 23616 1584 23644
rect 1578 23604 1584 23616
rect 1636 23604 1642 23656
rect 5445 23647 5503 23653
rect 5445 23613 5457 23647
rect 5491 23644 5503 23647
rect 5997 23647 6055 23653
rect 5997 23644 6009 23647
rect 5491 23616 6009 23644
rect 5491 23613 5503 23616
rect 5445 23607 5503 23613
rect 5997 23613 6009 23616
rect 6043 23644 6055 23647
rect 7098 23644 7104 23656
rect 6043 23616 7104 23644
rect 6043 23613 6055 23616
rect 5997 23607 6055 23613
rect 7098 23604 7104 23616
rect 7156 23644 7162 23656
rect 9950 23644 9956 23656
rect 7156 23616 9956 23644
rect 7156 23604 7162 23616
rect 9950 23604 9956 23616
rect 10008 23604 10014 23656
rect 11146 23604 11152 23656
rect 11204 23644 11210 23656
rect 12728 23644 12756 23752
rect 14090 23740 14096 23752
rect 14148 23740 14154 23792
rect 14185 23783 14243 23789
rect 14185 23749 14197 23783
rect 14231 23780 14243 23783
rect 14274 23780 14280 23792
rect 14231 23752 14280 23780
rect 14231 23749 14243 23752
rect 14185 23743 14243 23749
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 14550 23740 14556 23792
rect 14608 23780 14614 23792
rect 15013 23783 15071 23789
rect 15013 23780 15025 23783
rect 14608 23752 15025 23780
rect 14608 23740 14614 23752
rect 15013 23749 15025 23752
rect 15059 23749 15071 23783
rect 15013 23743 15071 23749
rect 15229 23783 15287 23789
rect 15229 23749 15241 23783
rect 15275 23780 15287 23783
rect 15654 23780 15660 23792
rect 15275 23752 15660 23780
rect 15275 23749 15287 23752
rect 15229 23743 15287 23749
rect 15654 23740 15660 23752
rect 15712 23740 15718 23792
rect 16666 23780 16672 23792
rect 15948 23752 16672 23780
rect 12805 23715 12863 23721
rect 12805 23681 12817 23715
rect 12851 23681 12863 23715
rect 13446 23712 13452 23724
rect 13359 23684 13452 23712
rect 12805 23675 12863 23681
rect 11204 23616 12756 23644
rect 11204 23604 11210 23616
rect 5350 23536 5356 23588
rect 5408 23576 5414 23588
rect 8389 23579 8447 23585
rect 5408 23548 8340 23576
rect 5408 23536 5414 23548
rect 7834 23508 7840 23520
rect 7795 23480 7840 23508
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 8312 23508 8340 23548
rect 8389 23545 8401 23579
rect 8435 23576 8447 23579
rect 9582 23576 9588 23588
rect 8435 23548 9588 23576
rect 8435 23545 8447 23548
rect 8389 23539 8447 23545
rect 9582 23536 9588 23548
rect 9640 23536 9646 23588
rect 12820 23576 12848 23675
rect 13446 23672 13452 23684
rect 13504 23712 13510 23724
rect 14366 23712 14372 23724
rect 13504 23684 14372 23712
rect 13504 23672 13510 23684
rect 14366 23672 14372 23684
rect 14424 23672 14430 23724
rect 15102 23712 15108 23724
rect 14752 23684 15108 23712
rect 14752 23656 14780 23684
rect 15102 23672 15108 23684
rect 15160 23672 15166 23724
rect 15838 23712 15844 23724
rect 15799 23684 15844 23712
rect 15838 23672 15844 23684
rect 15896 23672 15902 23724
rect 15948 23721 15976 23752
rect 16666 23740 16672 23752
rect 16724 23740 16730 23792
rect 16850 23740 16856 23792
rect 16908 23780 16914 23792
rect 17773 23783 17831 23789
rect 16908 23752 17540 23780
rect 16908 23740 16914 23752
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23681 15991 23715
rect 16114 23712 16120 23724
rect 16075 23684 16120 23712
rect 15933 23675 15991 23681
rect 16114 23672 16120 23684
rect 16172 23672 16178 23724
rect 16206 23672 16212 23724
rect 16264 23712 16270 23724
rect 16264 23684 17080 23712
rect 16264 23672 16270 23684
rect 13354 23604 13360 23656
rect 13412 23644 13418 23656
rect 13725 23647 13783 23653
rect 13725 23644 13737 23647
rect 13412 23616 13737 23644
rect 13412 23604 13418 23616
rect 13725 23613 13737 23616
rect 13771 23644 13783 23647
rect 14734 23644 14740 23656
rect 13771 23616 14740 23644
rect 13771 23613 13783 23616
rect 13725 23607 13783 23613
rect 14734 23604 14740 23616
rect 14792 23604 14798 23656
rect 16758 23644 16764 23656
rect 15166 23616 16764 23644
rect 15166 23588 15194 23616
rect 16758 23604 16764 23616
rect 16816 23604 16822 23656
rect 17052 23644 17080 23684
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 17221 23715 17279 23721
rect 17221 23712 17233 23715
rect 17184 23684 17233 23712
rect 17184 23672 17190 23684
rect 17221 23681 17233 23684
rect 17267 23681 17279 23715
rect 17221 23675 17279 23681
rect 17310 23672 17316 23724
rect 17368 23712 17374 23724
rect 17512 23721 17540 23752
rect 17773 23749 17785 23783
rect 17819 23780 17831 23783
rect 18138 23780 18144 23792
rect 17819 23752 18144 23780
rect 17819 23749 17831 23752
rect 17773 23743 17831 23749
rect 18138 23740 18144 23752
rect 18196 23740 18202 23792
rect 18322 23740 18328 23792
rect 18380 23740 18386 23792
rect 19150 23780 19156 23792
rect 18527 23752 19156 23780
rect 17497 23715 17555 23721
rect 17368 23684 17413 23712
rect 17368 23672 17374 23684
rect 17497 23681 17509 23715
rect 17543 23681 17555 23715
rect 17497 23675 17555 23681
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23712 17647 23715
rect 17678 23712 17684 23724
rect 17635 23684 17684 23712
rect 17635 23681 17647 23684
rect 17589 23675 17647 23681
rect 17678 23672 17684 23684
rect 17736 23672 17742 23724
rect 18414 23712 18420 23724
rect 17788 23684 18420 23712
rect 17788 23644 17816 23684
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 18527 23644 18555 23752
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 19444 23780 19472 23820
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 21266 23808 21272 23860
rect 21324 23848 21330 23860
rect 21542 23848 21548 23860
rect 21324 23820 21548 23848
rect 21324 23808 21330 23820
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22370 23808 22376 23860
rect 22428 23848 22434 23860
rect 26878 23848 26884 23860
rect 22428 23820 26884 23848
rect 22428 23808 22434 23820
rect 26878 23808 26884 23820
rect 26936 23808 26942 23860
rect 27246 23808 27252 23860
rect 27304 23848 27310 23860
rect 27304 23820 27449 23848
rect 27304 23808 27310 23820
rect 19794 23780 19800 23792
rect 19260 23752 19472 23780
rect 19719 23752 19800 23780
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 18785 23715 18843 23721
rect 18656 23684 18701 23712
rect 18656 23672 18662 23684
rect 18785 23681 18797 23715
rect 18831 23712 18843 23715
rect 19260 23712 19288 23752
rect 19429 23715 19487 23721
rect 19429 23712 19441 23715
rect 18831 23684 19288 23712
rect 19352 23684 19441 23712
rect 18831 23681 18843 23684
rect 18785 23675 18843 23681
rect 19168 23656 19196 23684
rect 17052 23616 17816 23644
rect 17906 23616 18555 23644
rect 18693 23647 18751 23653
rect 14274 23576 14280 23588
rect 12820 23548 14280 23576
rect 14274 23536 14280 23548
rect 14332 23536 14338 23588
rect 14553 23579 14611 23585
rect 14553 23545 14565 23579
rect 14599 23576 14611 23579
rect 14826 23576 14832 23588
rect 14599 23548 14832 23576
rect 14599 23545 14611 23548
rect 14553 23539 14611 23545
rect 14826 23536 14832 23548
rect 14884 23536 14890 23588
rect 15102 23536 15108 23588
rect 15160 23548 15194 23588
rect 15160 23536 15166 23548
rect 15286 23536 15292 23588
rect 15344 23576 15350 23588
rect 16114 23576 16120 23588
rect 15344 23548 16120 23576
rect 15344 23536 15350 23548
rect 16114 23536 16120 23548
rect 16172 23536 16178 23588
rect 16224 23548 16528 23576
rect 8846 23508 8852 23520
rect 8312 23480 8852 23508
rect 8846 23468 8852 23480
rect 8904 23468 8910 23520
rect 10594 23508 10600 23520
rect 10555 23480 10600 23508
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 11057 23511 11115 23517
rect 11057 23508 11069 23511
rect 10836 23480 11069 23508
rect 10836 23468 10842 23480
rect 11057 23477 11069 23480
rect 11103 23508 11115 23511
rect 11974 23508 11980 23520
rect 11103 23480 11980 23508
rect 11103 23477 11115 23480
rect 11057 23471 11115 23477
rect 11974 23468 11980 23480
rect 12032 23468 12038 23520
rect 12158 23468 12164 23520
rect 12216 23508 12222 23520
rect 12434 23508 12440 23520
rect 12216 23480 12440 23508
rect 12216 23468 12222 23480
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 12986 23508 12992 23520
rect 12947 23480 12992 23508
rect 12986 23468 12992 23480
rect 13044 23468 13050 23520
rect 13538 23508 13544 23520
rect 13499 23480 13544 23508
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 13630 23468 13636 23520
rect 13688 23508 13694 23520
rect 13688 23480 13733 23508
rect 13688 23468 13694 23480
rect 13906 23468 13912 23520
rect 13964 23508 13970 23520
rect 14090 23508 14096 23520
rect 13964 23480 14096 23508
rect 13964 23468 13970 23480
rect 14090 23468 14096 23480
rect 14148 23468 14154 23520
rect 14182 23468 14188 23520
rect 14240 23508 14246 23520
rect 14369 23511 14427 23517
rect 14369 23508 14381 23511
rect 14240 23480 14381 23508
rect 14240 23468 14246 23480
rect 14369 23477 14381 23480
rect 14415 23477 14427 23511
rect 14369 23471 14427 23477
rect 15197 23511 15255 23517
rect 15197 23477 15209 23511
rect 15243 23508 15255 23511
rect 16224 23508 16252 23548
rect 15243 23480 16252 23508
rect 16301 23511 16359 23517
rect 15243 23477 15255 23480
rect 15197 23471 15255 23477
rect 16301 23477 16313 23511
rect 16347 23508 16359 23511
rect 16390 23508 16396 23520
rect 16347 23480 16396 23508
rect 16347 23477 16359 23480
rect 16301 23471 16359 23477
rect 16390 23468 16396 23480
rect 16448 23468 16454 23520
rect 16500 23508 16528 23548
rect 16574 23536 16580 23588
rect 16632 23576 16638 23588
rect 17906 23576 17934 23616
rect 18693 23613 18705 23647
rect 18739 23644 18751 23647
rect 19058 23644 19064 23656
rect 18739 23616 19064 23644
rect 18739 23613 18751 23616
rect 18693 23607 18751 23613
rect 19058 23604 19064 23616
rect 19116 23604 19122 23656
rect 19150 23604 19156 23656
rect 19208 23604 19214 23656
rect 19242 23604 19248 23656
rect 19300 23644 19306 23656
rect 19352 23644 19380 23684
rect 19429 23681 19441 23684
rect 19475 23681 19487 23715
rect 19429 23675 19487 23681
rect 19518 23672 19524 23724
rect 19576 23712 19582 23724
rect 19719 23721 19747 23752
rect 19794 23740 19800 23752
rect 19852 23740 19858 23792
rect 20990 23780 20996 23792
rect 19704 23715 19762 23721
rect 19576 23684 19621 23712
rect 19576 23672 19582 23684
rect 19704 23681 19716 23715
rect 19750 23681 19762 23715
rect 19892 23706 19898 23758
rect 19950 23706 19956 23758
rect 19996 23752 20484 23780
rect 19893 23703 19905 23706
rect 19939 23703 19951 23706
rect 19893 23697 19951 23703
rect 19704 23675 19762 23681
rect 19996 23644 20024 23752
rect 20349 23715 20407 23721
rect 20349 23712 20361 23715
rect 19300 23616 19380 23644
rect 19444 23616 20024 23644
rect 20088 23684 20361 23712
rect 19300 23604 19306 23616
rect 18138 23576 18144 23588
rect 16632 23548 17934 23576
rect 17972 23548 18144 23576
rect 16632 23536 16638 23548
rect 17972 23508 18000 23548
rect 18138 23536 18144 23548
rect 18196 23536 18202 23588
rect 18322 23536 18328 23588
rect 18380 23576 18386 23588
rect 19444 23576 19472 23616
rect 18380 23548 19472 23576
rect 19613 23579 19671 23585
rect 18380 23536 18386 23548
rect 19613 23545 19625 23579
rect 19659 23545 19671 23579
rect 19613 23539 19671 23545
rect 16500 23480 18000 23508
rect 18046 23468 18052 23520
rect 18104 23508 18110 23520
rect 19245 23511 19303 23517
rect 19245 23508 19257 23511
rect 18104 23480 19257 23508
rect 18104 23468 18110 23480
rect 19245 23477 19257 23480
rect 19291 23477 19303 23511
rect 19628 23508 19656 23539
rect 19794 23536 19800 23588
rect 19852 23576 19858 23588
rect 20088 23576 20116 23684
rect 20349 23681 20361 23684
rect 20395 23681 20407 23715
rect 20456 23712 20484 23752
rect 20640 23752 20852 23780
rect 20951 23752 20996 23780
rect 20640 23724 20668 23752
rect 20512 23715 20570 23721
rect 20512 23712 20524 23715
rect 20456 23684 20524 23712
rect 20349 23675 20407 23681
rect 20512 23681 20524 23684
rect 20558 23681 20570 23715
rect 20512 23675 20570 23681
rect 20612 23718 20670 23724
rect 20612 23684 20624 23718
rect 20658 23684 20670 23718
rect 20737 23715 20795 23721
rect 20737 23712 20749 23715
rect 20612 23678 20670 23684
rect 20732 23681 20749 23712
rect 20783 23681 20795 23715
rect 20824 23712 20852 23752
rect 20990 23740 20996 23752
rect 21048 23740 21054 23792
rect 21358 23740 21364 23792
rect 21416 23780 21422 23792
rect 21726 23780 21732 23792
rect 21416 23752 21732 23780
rect 21416 23740 21422 23752
rect 21726 23740 21732 23752
rect 21784 23740 21790 23792
rect 22922 23780 22928 23792
rect 21836 23752 22928 23780
rect 20824 23684 21496 23712
rect 20732 23675 20795 23681
rect 20732 23644 20760 23675
rect 21468 23656 21496 23684
rect 21082 23644 21088 23656
rect 20732 23616 21088 23644
rect 21082 23604 21088 23616
rect 21140 23604 21146 23656
rect 21450 23604 21456 23656
rect 21508 23604 21514 23656
rect 19852 23548 20116 23576
rect 19852 23536 19858 23548
rect 20254 23536 20260 23588
rect 20312 23576 20318 23588
rect 21836 23576 21864 23752
rect 22922 23740 22928 23752
rect 22980 23740 22986 23792
rect 23382 23780 23388 23792
rect 23216 23752 23388 23780
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23681 22063 23715
rect 22186 23712 22192 23724
rect 22147 23684 22192 23712
rect 22005 23675 22063 23681
rect 22020 23644 22048 23675
rect 22186 23672 22192 23684
rect 22244 23672 22250 23724
rect 22462 23712 22468 23724
rect 22423 23684 22468 23712
rect 22462 23672 22468 23684
rect 22520 23672 22526 23724
rect 23216 23721 23244 23752
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 23750 23740 23756 23792
rect 23808 23780 23814 23792
rect 23808 23752 23966 23780
rect 23808 23740 23814 23752
rect 24854 23740 24860 23792
rect 24912 23780 24918 23792
rect 25225 23783 25283 23789
rect 25225 23780 25237 23783
rect 24912 23752 25237 23780
rect 24912 23740 24918 23752
rect 25225 23749 25237 23752
rect 25271 23780 25283 23783
rect 25682 23780 25688 23792
rect 25271 23752 25688 23780
rect 25271 23749 25283 23752
rect 25225 23743 25283 23749
rect 25682 23740 25688 23752
rect 25740 23740 25746 23792
rect 25866 23740 25872 23792
rect 25924 23780 25930 23792
rect 26234 23780 26240 23792
rect 25924 23752 26240 23780
rect 25924 23740 25930 23752
rect 26234 23740 26240 23752
rect 26292 23740 26298 23792
rect 26786 23740 26792 23792
rect 26844 23780 26850 23792
rect 27421 23780 27449 23820
rect 27522 23808 27528 23860
rect 27580 23848 27586 23860
rect 27580 23820 28764 23848
rect 27580 23808 27586 23820
rect 28442 23780 28448 23792
rect 26844 23752 27384 23780
rect 27421 23752 27844 23780
rect 26844 23740 26850 23752
rect 23201 23715 23259 23721
rect 23201 23681 23213 23715
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 25498 23672 25504 23724
rect 25556 23712 25562 23724
rect 26050 23712 26056 23724
rect 25556 23684 26056 23712
rect 25556 23672 25562 23684
rect 26050 23672 26056 23684
rect 26108 23672 26114 23724
rect 26159 23684 26353 23712
rect 22738 23644 22744 23656
rect 22020 23616 22744 23644
rect 22738 23604 22744 23616
rect 22796 23604 22802 23656
rect 23474 23644 23480 23656
rect 23435 23616 23480 23644
rect 23474 23604 23480 23616
rect 23532 23604 23538 23656
rect 23566 23604 23572 23656
rect 23624 23644 23630 23656
rect 26159 23644 26187 23684
rect 23624 23616 26187 23644
rect 26237 23647 26295 23653
rect 23624 23604 23630 23616
rect 26237 23613 26249 23647
rect 26283 23613 26295 23647
rect 26237 23607 26295 23613
rect 20312 23548 21864 23576
rect 20312 23536 20318 23548
rect 21910 23536 21916 23588
rect 21968 23576 21974 23588
rect 22281 23579 22339 23585
rect 22281 23576 22293 23579
rect 21968 23548 22293 23576
rect 21968 23536 21974 23548
rect 22281 23545 22293 23548
rect 22327 23545 22339 23579
rect 22281 23539 22339 23545
rect 22646 23536 22652 23588
rect 22704 23576 22710 23588
rect 23198 23576 23204 23588
rect 22704 23548 23204 23576
rect 22704 23536 22710 23548
rect 23198 23536 23204 23548
rect 23256 23536 23262 23588
rect 26252 23576 26280 23607
rect 24826 23548 26280 23576
rect 26325 23576 26353 23684
rect 26970 23672 26976 23724
rect 27028 23712 27034 23724
rect 27356 23721 27384 23752
rect 27157 23715 27215 23721
rect 27157 23712 27169 23715
rect 27028 23684 27169 23712
rect 27028 23672 27034 23684
rect 27157 23681 27169 23684
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 27617 23715 27675 23721
rect 27617 23681 27629 23715
rect 27663 23712 27675 23715
rect 27706 23712 27712 23724
rect 27663 23684 27712 23712
rect 27663 23681 27675 23684
rect 27617 23675 27675 23681
rect 26510 23644 26516 23656
rect 26471 23616 26516 23644
rect 26510 23604 26516 23616
rect 26568 23604 26574 23656
rect 26694 23604 26700 23656
rect 26752 23644 26758 23656
rect 27632 23644 27660 23675
rect 27706 23672 27712 23684
rect 27764 23672 27770 23724
rect 26752 23616 27660 23644
rect 27816 23644 27844 23752
rect 27908 23752 28448 23780
rect 27908 23721 27936 23752
rect 28442 23740 28448 23752
rect 28500 23740 28506 23792
rect 27893 23715 27951 23721
rect 27893 23681 27905 23715
rect 27939 23681 27951 23715
rect 27893 23675 27951 23681
rect 27982 23672 27988 23724
rect 28040 23712 28046 23724
rect 28350 23712 28356 23724
rect 28040 23684 28356 23712
rect 28040 23672 28046 23684
rect 28350 23672 28356 23684
rect 28408 23672 28414 23724
rect 28534 23672 28540 23724
rect 28592 23712 28598 23724
rect 28736 23721 28764 23820
rect 29086 23808 29092 23860
rect 29144 23848 29150 23860
rect 29549 23851 29607 23857
rect 29549 23848 29561 23851
rect 29144 23820 29561 23848
rect 29144 23808 29150 23820
rect 29549 23817 29561 23820
rect 29595 23817 29607 23851
rect 29549 23811 29607 23817
rect 29638 23808 29644 23860
rect 29696 23848 29702 23860
rect 30190 23848 30196 23860
rect 29696 23820 30196 23848
rect 29696 23808 29702 23820
rect 30190 23808 30196 23820
rect 30248 23808 30254 23860
rect 30650 23848 30656 23860
rect 30611 23820 30656 23848
rect 30650 23808 30656 23820
rect 30708 23808 30714 23860
rect 31205 23783 31263 23789
rect 29748 23752 31156 23780
rect 28629 23715 28687 23721
rect 28629 23712 28641 23715
rect 28592 23684 28641 23712
rect 28592 23672 28598 23684
rect 28629 23681 28641 23684
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23681 28779 23715
rect 28721 23675 28779 23681
rect 28902 23672 28908 23724
rect 28960 23712 28966 23724
rect 28960 23684 29224 23712
rect 28960 23672 28966 23684
rect 28997 23647 29055 23653
rect 28997 23644 29009 23647
rect 27816 23616 29009 23644
rect 26752 23604 26758 23616
rect 28997 23613 29009 23616
rect 29043 23613 29055 23647
rect 28997 23607 29055 23613
rect 29089 23647 29147 23653
rect 29089 23613 29101 23647
rect 29135 23613 29147 23647
rect 29196 23644 29224 23684
rect 29546 23672 29552 23724
rect 29604 23712 29610 23724
rect 29748 23721 29776 23752
rect 29733 23715 29791 23721
rect 29733 23712 29745 23715
rect 29604 23684 29745 23712
rect 29604 23672 29610 23684
rect 29733 23681 29745 23684
rect 29779 23681 29791 23715
rect 30006 23712 30012 23724
rect 29967 23684 30012 23712
rect 29733 23675 29791 23681
rect 30006 23672 30012 23684
rect 30064 23672 30070 23724
rect 30193 23715 30251 23721
rect 30193 23681 30205 23715
rect 30239 23712 30251 23715
rect 30558 23712 30564 23724
rect 30239 23684 30564 23712
rect 30239 23681 30251 23684
rect 30193 23675 30251 23681
rect 30558 23672 30564 23684
rect 30616 23672 30622 23724
rect 30926 23712 30932 23724
rect 30887 23684 30932 23712
rect 30926 23672 30932 23684
rect 30984 23672 30990 23724
rect 31128 23712 31156 23752
rect 31205 23749 31217 23783
rect 31251 23780 31263 23783
rect 31386 23780 31392 23792
rect 31251 23752 31392 23780
rect 31251 23749 31263 23752
rect 31205 23743 31263 23749
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 32214 23712 32220 23724
rect 31128 23684 32220 23712
rect 32214 23672 32220 23684
rect 32272 23672 32278 23724
rect 30837 23647 30895 23653
rect 30837 23644 30849 23647
rect 29196 23616 30849 23644
rect 29089 23607 29147 23613
rect 30837 23613 30849 23616
rect 30883 23613 30895 23647
rect 31294 23644 31300 23656
rect 31255 23616 31300 23644
rect 30837 23607 30895 23613
rect 28445 23579 28503 23585
rect 28445 23576 28457 23579
rect 26325 23548 28457 23576
rect 21542 23508 21548 23520
rect 19628 23480 21548 23508
rect 19245 23471 19303 23477
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 22370 23508 22376 23520
rect 22331 23480 22376 23508
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 22738 23508 22744 23520
rect 22699 23480 22744 23508
rect 22738 23468 22744 23480
rect 22796 23468 22802 23520
rect 23106 23468 23112 23520
rect 23164 23508 23170 23520
rect 24118 23508 24124 23520
rect 23164 23480 24124 23508
rect 23164 23468 23170 23480
rect 24118 23468 24124 23480
rect 24176 23508 24182 23520
rect 24826 23508 24854 23548
rect 28445 23545 28457 23548
rect 28491 23545 28503 23579
rect 28445 23539 28503 23545
rect 28534 23536 28540 23588
rect 28592 23576 28598 23588
rect 28718 23576 28724 23588
rect 28592 23548 28724 23576
rect 28592 23536 28598 23548
rect 28718 23536 28724 23548
rect 28776 23536 28782 23588
rect 29104 23576 29132 23607
rect 31294 23604 31300 23616
rect 31352 23604 31358 23656
rect 31386 23604 31392 23656
rect 31444 23644 31450 23656
rect 32398 23644 32404 23656
rect 31444 23616 32404 23644
rect 31444 23604 31450 23616
rect 32398 23604 32404 23616
rect 32456 23604 32462 23656
rect 29454 23576 29460 23588
rect 29104 23548 29460 23576
rect 24176 23480 24854 23508
rect 24176 23468 24182 23480
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 25222 23508 25228 23520
rect 25096 23480 25228 23508
rect 25096 23468 25102 23480
rect 25222 23468 25228 23480
rect 25280 23468 25286 23520
rect 25314 23468 25320 23520
rect 25372 23508 25378 23520
rect 29104 23508 29132 23548
rect 29454 23536 29460 23548
rect 29512 23536 29518 23588
rect 29730 23536 29736 23588
rect 29788 23576 29794 23588
rect 30558 23576 30564 23588
rect 29788 23548 30564 23576
rect 29788 23536 29794 23548
rect 30558 23536 30564 23548
rect 30616 23536 30622 23588
rect 25372 23480 29132 23508
rect 25372 23468 25378 23480
rect 29362 23468 29368 23520
rect 29420 23508 29426 23520
rect 30282 23508 30288 23520
rect 29420 23480 30288 23508
rect 29420 23468 29426 23480
rect 30282 23468 30288 23480
rect 30340 23468 30346 23520
rect 1104 23418 31832 23440
rect 1104 23366 4791 23418
rect 4843 23366 4855 23418
rect 4907 23366 4919 23418
rect 4971 23366 4983 23418
rect 5035 23366 5047 23418
rect 5099 23366 12473 23418
rect 12525 23366 12537 23418
rect 12589 23366 12601 23418
rect 12653 23366 12665 23418
rect 12717 23366 12729 23418
rect 12781 23366 20155 23418
rect 20207 23366 20219 23418
rect 20271 23366 20283 23418
rect 20335 23366 20347 23418
rect 20399 23366 20411 23418
rect 20463 23366 27837 23418
rect 27889 23366 27901 23418
rect 27953 23366 27965 23418
rect 28017 23366 28029 23418
rect 28081 23366 28093 23418
rect 28145 23366 31832 23418
rect 1104 23344 31832 23366
rect 4157 23307 4215 23313
rect 4157 23273 4169 23307
rect 4203 23304 4215 23307
rect 4246 23304 4252 23316
rect 4203 23276 4252 23304
rect 4203 23273 4215 23276
rect 4157 23267 4215 23273
rect 4246 23264 4252 23276
rect 4304 23264 4310 23316
rect 5810 23304 5816 23316
rect 5771 23276 5816 23304
rect 5810 23264 5816 23276
rect 5868 23264 5874 23316
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 8478 23304 8484 23316
rect 5960 23276 8484 23304
rect 5960 23264 5966 23276
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 9217 23307 9275 23313
rect 9217 23273 9229 23307
rect 9263 23304 9275 23307
rect 9582 23304 9588 23316
rect 9263 23276 9588 23304
rect 9263 23273 9275 23276
rect 9217 23267 9275 23273
rect 9582 23264 9588 23276
rect 9640 23304 9646 23316
rect 9677 23307 9735 23313
rect 9677 23304 9689 23307
rect 9640 23276 9689 23304
rect 9640 23264 9646 23276
rect 9677 23273 9689 23276
rect 9723 23273 9735 23307
rect 9677 23267 9735 23273
rect 10321 23307 10379 23313
rect 10321 23273 10333 23307
rect 10367 23304 10379 23307
rect 10594 23304 10600 23316
rect 10367 23276 10600 23304
rect 10367 23273 10379 23276
rect 10321 23267 10379 23273
rect 10594 23264 10600 23276
rect 10652 23264 10658 23316
rect 12434 23304 12440 23316
rect 12176 23276 12440 23304
rect 4709 23239 4767 23245
rect 4709 23205 4721 23239
rect 4755 23236 4767 23239
rect 10134 23236 10140 23248
rect 4755 23208 10140 23236
rect 4755 23205 4767 23208
rect 4709 23199 4767 23205
rect 10134 23196 10140 23208
rect 10192 23196 10198 23248
rect 11054 23196 11060 23248
rect 11112 23236 11118 23248
rect 11333 23239 11391 23245
rect 11333 23236 11345 23239
rect 11112 23208 11345 23236
rect 11112 23196 11118 23208
rect 11333 23205 11345 23208
rect 11379 23205 11391 23239
rect 11333 23199 11391 23205
rect 11422 23196 11428 23248
rect 11480 23236 11486 23248
rect 12176 23236 12204 23276
rect 12434 23264 12440 23276
rect 12492 23304 12498 23316
rect 13630 23304 13636 23316
rect 12492 23276 13636 23304
rect 12492 23264 12498 23276
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 14366 23264 14372 23316
rect 14424 23304 14430 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14424 23276 14657 23304
rect 14424 23264 14430 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 14826 23304 14832 23316
rect 14787 23276 14832 23304
rect 14645 23267 14703 23273
rect 11480 23208 12204 23236
rect 12621 23239 12679 23245
rect 11480 23196 11486 23208
rect 12621 23205 12633 23239
rect 12667 23205 12679 23239
rect 12621 23199 12679 23205
rect 5442 23128 5448 23180
rect 5500 23168 5506 23180
rect 9582 23168 9588 23180
rect 5500 23140 9588 23168
rect 5500 23128 5506 23140
rect 9582 23128 9588 23140
rect 9640 23128 9646 23180
rect 12636 23168 12664 23199
rect 13722 23196 13728 23248
rect 13780 23236 13786 23248
rect 14182 23236 14188 23248
rect 13780 23208 14188 23236
rect 13780 23196 13786 23208
rect 14182 23196 14188 23208
rect 14240 23196 14246 23248
rect 14660 23236 14688 23267
rect 14826 23264 14832 23276
rect 14884 23264 14890 23316
rect 14918 23264 14924 23316
rect 14976 23304 14982 23316
rect 15286 23304 15292 23316
rect 14976 23276 15292 23304
rect 14976 23264 14982 23276
rect 15286 23264 15292 23276
rect 15344 23264 15350 23316
rect 15838 23264 15844 23316
rect 15896 23304 15902 23316
rect 16574 23304 16580 23316
rect 15896 23276 16580 23304
rect 15896 23264 15902 23276
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 16666 23264 16672 23316
rect 16724 23304 16730 23316
rect 16724 23276 18644 23304
rect 16724 23264 16730 23276
rect 14660 23208 14872 23236
rect 14844 23180 14872 23208
rect 15378 23196 15384 23248
rect 15436 23236 15442 23248
rect 15473 23239 15531 23245
rect 15473 23236 15485 23239
rect 15436 23208 15485 23236
rect 15436 23196 15442 23208
rect 15473 23205 15485 23208
rect 15519 23205 15531 23239
rect 15473 23199 15531 23205
rect 15580 23208 18276 23236
rect 11164 23140 12664 23168
rect 1578 23100 1584 23112
rect 1539 23072 1584 23100
rect 1578 23060 1584 23072
rect 1636 23060 1642 23112
rect 5074 23060 5080 23112
rect 5132 23100 5138 23112
rect 5261 23103 5319 23109
rect 5261 23100 5273 23103
rect 5132 23072 5273 23100
rect 5132 23060 5138 23072
rect 5261 23069 5273 23072
rect 5307 23100 5319 23103
rect 8018 23100 8024 23112
rect 5307 23072 8024 23100
rect 5307 23069 5319 23072
rect 5261 23063 5319 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 9398 23060 9404 23112
rect 9456 23100 9462 23112
rect 10502 23100 10508 23112
rect 9456 23072 10508 23100
rect 9456 23060 9462 23072
rect 10502 23060 10508 23072
rect 10560 23060 10566 23112
rect 6365 23035 6423 23041
rect 6365 23001 6377 23035
rect 6411 23032 6423 23035
rect 6546 23032 6552 23044
rect 6411 23004 6552 23032
rect 6411 23001 6423 23004
rect 6365 22995 6423 23001
rect 6546 22992 6552 23004
rect 6604 22992 6610 23044
rect 6638 22992 6644 23044
rect 6696 23032 6702 23044
rect 11164 23032 11192 23140
rect 12986 23128 12992 23180
rect 13044 23168 13050 23180
rect 13044 23140 14780 23168
rect 13044 23128 13050 23140
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 11333 23103 11391 23109
rect 11333 23100 11345 23103
rect 11296 23072 11345 23100
rect 11296 23060 11302 23072
rect 11333 23069 11345 23072
rect 11379 23069 11391 23103
rect 11333 23063 11391 23069
rect 6696 23004 11192 23032
rect 11348 23032 11376 23063
rect 11422 23060 11428 23112
rect 11480 23100 11486 23112
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 11480 23072 11529 23100
rect 11480 23060 11486 23072
rect 11517 23069 11529 23072
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 11606 23060 11612 23112
rect 11664 23100 11670 23112
rect 11977 23103 12035 23109
rect 11977 23100 11989 23103
rect 11664 23072 11989 23100
rect 11664 23060 11670 23072
rect 11977 23069 11989 23072
rect 12023 23069 12035 23103
rect 11977 23063 12035 23069
rect 12158 23060 12164 23112
rect 12216 23100 12222 23112
rect 12621 23103 12679 23109
rect 12621 23100 12633 23103
rect 12216 23072 12633 23100
rect 12216 23060 12222 23072
rect 12621 23069 12633 23072
rect 12667 23069 12679 23103
rect 12802 23100 12808 23112
rect 12763 23072 12808 23100
rect 12621 23063 12679 23069
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 12897 23103 12955 23109
rect 12897 23069 12909 23103
rect 12943 23100 12955 23103
rect 13446 23100 13452 23112
rect 12943 23072 13452 23100
rect 12943 23069 12955 23072
rect 12897 23063 12955 23069
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 13538 23060 13544 23112
rect 13596 23100 13602 23112
rect 13596 23072 13641 23100
rect 13596 23060 13602 23072
rect 13906 23060 13912 23112
rect 13964 23100 13970 23112
rect 14366 23100 14372 23112
rect 13964 23072 14372 23100
rect 13964 23060 13970 23072
rect 14366 23060 14372 23072
rect 14424 23100 14430 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 14424 23072 14473 23100
rect 14424 23060 14430 23072
rect 14461 23069 14473 23072
rect 14507 23069 14519 23103
rect 14642 23100 14648 23112
rect 14603 23072 14648 23100
rect 14461 23063 14519 23069
rect 14642 23060 14648 23072
rect 14700 23060 14706 23112
rect 14752 23100 14780 23140
rect 14826 23128 14832 23180
rect 14884 23128 14890 23180
rect 15580 23168 15608 23208
rect 14936 23140 15608 23168
rect 14936 23100 14964 23140
rect 16114 23128 16120 23180
rect 16172 23168 16178 23180
rect 17126 23168 17132 23180
rect 16172 23140 16344 23168
rect 16172 23128 16178 23140
rect 14752 23072 14964 23100
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23069 15439 23103
rect 15654 23100 15660 23112
rect 15615 23072 15660 23100
rect 15381 23063 15439 23069
rect 13357 23035 13415 23041
rect 13357 23032 13369 23035
rect 11348 23004 13369 23032
rect 6696 22992 6702 23004
rect 13357 23001 13369 23004
rect 13403 23001 13415 23035
rect 15286 23032 15292 23044
rect 15247 23004 15292 23032
rect 13357 22995 13415 23001
rect 15286 22992 15292 23004
rect 15344 22992 15350 23044
rect 15396 23032 15424 23063
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23100 15807 23103
rect 15838 23100 15844 23112
rect 15795 23072 15844 23100
rect 15795 23069 15807 23072
rect 15749 23063 15807 23069
rect 15838 23060 15844 23072
rect 15896 23060 15902 23112
rect 16206 23100 16212 23112
rect 16167 23072 16212 23100
rect 16206 23060 16212 23072
rect 16264 23060 16270 23112
rect 16316 23109 16344 23140
rect 16592 23140 17132 23168
rect 16301 23103 16359 23109
rect 16301 23069 16313 23103
rect 16347 23069 16359 23103
rect 16301 23063 16359 23069
rect 16390 23060 16396 23112
rect 16448 23100 16454 23112
rect 16592 23109 16620 23140
rect 17126 23128 17132 23140
rect 17184 23128 17190 23180
rect 17773 23171 17831 23177
rect 17773 23137 17785 23171
rect 17819 23168 17831 23171
rect 17862 23168 17868 23180
rect 17819 23140 17868 23168
rect 17819 23137 17831 23140
rect 17773 23131 17831 23137
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 18248 23177 18276 23208
rect 18414 23196 18420 23248
rect 18472 23196 18478 23248
rect 18616 23236 18644 23276
rect 19978 23264 19984 23316
rect 20036 23304 20042 23316
rect 20036 23276 21220 23304
rect 20036 23264 20042 23276
rect 18616 23208 19472 23236
rect 18233 23171 18291 23177
rect 18233 23137 18245 23171
rect 18279 23137 18291 23171
rect 18432 23168 18460 23196
rect 19334 23168 19340 23180
rect 18432 23140 18552 23168
rect 18233 23131 18291 23137
rect 16485 23103 16543 23109
rect 16485 23100 16497 23103
rect 16448 23072 16497 23100
rect 16448 23060 16454 23072
rect 16485 23069 16497 23072
rect 16531 23069 16543 23103
rect 16485 23063 16543 23069
rect 16577 23103 16635 23109
rect 16577 23069 16589 23103
rect 16623 23069 16635 23103
rect 16577 23063 16635 23069
rect 16761 23103 16819 23109
rect 16761 23069 16773 23103
rect 16807 23100 16819 23103
rect 16850 23100 16856 23112
rect 16807 23072 16856 23100
rect 16807 23069 16819 23072
rect 16761 23063 16819 23069
rect 15930 23032 15936 23044
rect 15396 23004 15936 23032
rect 15930 22992 15936 23004
rect 15988 22992 15994 23044
rect 16114 22992 16120 23044
rect 16172 23032 16178 23044
rect 16592 23032 16620 23063
rect 16850 23060 16856 23072
rect 16908 23060 16914 23112
rect 16942 23060 16948 23112
rect 17000 23100 17006 23112
rect 17221 23103 17279 23109
rect 17221 23100 17233 23103
rect 17000 23072 17233 23100
rect 17000 23060 17006 23072
rect 17221 23069 17233 23072
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 17310 23060 17316 23112
rect 17368 23100 17374 23112
rect 17494 23100 17500 23112
rect 17368 23072 17413 23100
rect 17455 23072 17500 23100
rect 17368 23060 17374 23072
rect 17494 23060 17500 23072
rect 17552 23060 17558 23112
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23100 17647 23103
rect 17678 23100 17684 23112
rect 17635 23072 17684 23100
rect 17635 23069 17647 23072
rect 17589 23063 17647 23069
rect 17678 23060 17684 23072
rect 17736 23060 17742 23112
rect 18524 23109 18552 23140
rect 18754 23140 19340 23168
rect 18754 23109 18782 23140
rect 19334 23128 19340 23140
rect 19392 23128 19398 23180
rect 19444 23168 19472 23208
rect 19518 23196 19524 23248
rect 19576 23236 19582 23248
rect 20806 23236 20812 23248
rect 19576 23208 20812 23236
rect 19576 23196 19582 23208
rect 20806 23196 20812 23208
rect 20864 23196 20870 23248
rect 21192 23236 21220 23276
rect 21266 23264 21272 23316
rect 21324 23304 21330 23316
rect 24854 23304 24860 23316
rect 21324 23276 24860 23304
rect 21324 23264 21330 23276
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 26786 23304 26792 23316
rect 24964 23276 26792 23304
rect 22554 23236 22560 23248
rect 21192 23208 22560 23236
rect 22554 23196 22560 23208
rect 22612 23196 22618 23248
rect 24026 23196 24032 23248
rect 24084 23236 24090 23248
rect 24964 23236 24992 23276
rect 26786 23264 26792 23276
rect 26844 23264 26850 23316
rect 27706 23264 27712 23316
rect 27764 23304 27770 23316
rect 28353 23307 28411 23313
rect 28353 23304 28365 23307
rect 27764 23276 28365 23304
rect 27764 23264 27770 23276
rect 28353 23273 28365 23276
rect 28399 23273 28411 23307
rect 28353 23267 28411 23273
rect 28534 23264 28540 23316
rect 28592 23304 28598 23316
rect 28629 23307 28687 23313
rect 28629 23304 28641 23307
rect 28592 23276 28641 23304
rect 28592 23264 28598 23276
rect 28629 23273 28641 23276
rect 28675 23273 28687 23307
rect 28810 23304 28816 23316
rect 28771 23276 28816 23304
rect 28629 23267 28687 23273
rect 28810 23264 28816 23276
rect 28868 23264 28874 23316
rect 29730 23264 29736 23316
rect 29788 23264 29794 23316
rect 30098 23264 30104 23316
rect 30156 23264 30162 23316
rect 30190 23264 30196 23316
rect 30248 23264 30254 23316
rect 24084 23208 24992 23236
rect 24084 23196 24090 23208
rect 26970 23196 26976 23248
rect 27028 23236 27034 23248
rect 27028 23208 27073 23236
rect 27028 23196 27034 23208
rect 27798 23196 27804 23248
rect 27856 23236 27862 23248
rect 29748 23236 29776 23264
rect 27856 23208 29776 23236
rect 27856 23196 27862 23208
rect 19444 23140 20116 23168
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23069 18475 23103
rect 18417 23063 18475 23069
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23069 18659 23103
rect 18601 23063 18659 23069
rect 18739 23103 18797 23109
rect 18739 23069 18751 23103
rect 18785 23069 18797 23103
rect 18739 23063 18797 23069
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23100 18935 23103
rect 19518 23100 19524 23112
rect 18923 23072 19524 23100
rect 18923 23069 18935 23072
rect 18877 23063 18935 23069
rect 16172 23004 16620 23032
rect 16172 22992 16178 23004
rect 17126 22992 17132 23044
rect 17184 23032 17190 23044
rect 17862 23032 17868 23044
rect 17184 23004 17868 23032
rect 17184 22992 17190 23004
rect 17862 22992 17868 23004
rect 17920 23032 17926 23044
rect 18432 23032 18460 23063
rect 17920 23004 18460 23032
rect 18616 23032 18644 23063
rect 19518 23060 19524 23072
rect 19576 23060 19582 23112
rect 19794 23060 19800 23112
rect 19852 23100 19858 23112
rect 20088 23109 20116 23140
rect 20346 23128 20352 23180
rect 20404 23168 20410 23180
rect 21450 23168 21456 23180
rect 20404 23140 21456 23168
rect 20404 23128 20410 23140
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 22094 23128 22100 23180
rect 22152 23168 22158 23180
rect 22281 23171 22339 23177
rect 22281 23168 22293 23171
rect 22152 23140 22293 23168
rect 22152 23128 22158 23140
rect 22281 23137 22293 23140
rect 22327 23137 22339 23171
rect 23106 23168 23112 23180
rect 22281 23131 22339 23137
rect 22579 23140 23112 23168
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 19852 23072 19901 23100
rect 19852 23060 19858 23072
rect 19889 23069 19901 23072
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23069 20131 23103
rect 20073 23063 20131 23069
rect 20165 23103 20223 23109
rect 20165 23069 20177 23103
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 20257 23103 20315 23109
rect 20257 23069 20269 23103
rect 20303 23069 20315 23103
rect 20257 23063 20315 23069
rect 19058 23032 19064 23044
rect 18616 23004 19064 23032
rect 17920 22992 17926 23004
rect 19058 22992 19064 23004
rect 19116 22992 19122 23044
rect 19150 22992 19156 23044
rect 19208 23032 19214 23044
rect 20180 23032 20208 23063
rect 19208 23004 20208 23032
rect 19208 22992 19214 23004
rect 6086 22924 6092 22976
rect 6144 22964 6150 22976
rect 6825 22967 6883 22973
rect 6825 22964 6837 22967
rect 6144 22936 6837 22964
rect 6144 22924 6150 22936
rect 6825 22933 6837 22936
rect 6871 22964 6883 22967
rect 7377 22967 7435 22973
rect 7377 22964 7389 22967
rect 6871 22936 7389 22964
rect 6871 22933 6883 22936
rect 6825 22927 6883 22933
rect 7377 22933 7389 22936
rect 7423 22933 7435 22967
rect 7377 22927 7435 22933
rect 7466 22924 7472 22976
rect 7524 22964 7530 22976
rect 7650 22964 7656 22976
rect 7524 22936 7656 22964
rect 7524 22924 7530 22936
rect 7650 22924 7656 22936
rect 7708 22964 7714 22976
rect 7929 22967 7987 22973
rect 7929 22964 7941 22967
rect 7708 22936 7941 22964
rect 7708 22924 7714 22936
rect 7929 22933 7941 22936
rect 7975 22933 7987 22967
rect 7929 22927 7987 22933
rect 8573 22967 8631 22973
rect 8573 22933 8585 22967
rect 8619 22964 8631 22967
rect 9030 22964 9036 22976
rect 8619 22936 9036 22964
rect 8619 22933 8631 22936
rect 8573 22927 8631 22933
rect 9030 22924 9036 22936
rect 9088 22924 9094 22976
rect 10870 22964 10876 22976
rect 10783 22936 10876 22964
rect 10870 22924 10876 22936
rect 10928 22964 10934 22976
rect 11698 22964 11704 22976
rect 10928 22936 11704 22964
rect 10928 22924 10934 22936
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 12066 22964 12072 22976
rect 12027 22936 12072 22964
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 12158 22924 12164 22976
rect 12216 22964 12222 22976
rect 13262 22964 13268 22976
rect 12216 22936 13268 22964
rect 12216 22924 12222 22936
rect 13262 22924 13268 22936
rect 13320 22964 13326 22976
rect 13725 22967 13783 22973
rect 13725 22964 13737 22967
rect 13320 22936 13737 22964
rect 13320 22924 13326 22936
rect 13725 22933 13737 22936
rect 13771 22933 13783 22967
rect 13725 22927 13783 22933
rect 14090 22924 14096 22976
rect 14148 22964 14154 22976
rect 16666 22964 16672 22976
rect 14148 22936 16672 22964
rect 14148 22924 14154 22936
rect 16666 22924 16672 22936
rect 16724 22924 16730 22976
rect 16758 22924 16764 22976
rect 16816 22964 16822 22976
rect 20272 22964 20300 23063
rect 20438 23060 20444 23112
rect 20496 23100 20502 23112
rect 21085 23103 21143 23109
rect 21085 23100 21097 23103
rect 20496 23072 21097 23100
rect 20496 23060 20502 23072
rect 21085 23069 21097 23072
rect 21131 23069 21143 23103
rect 21266 23100 21272 23112
rect 21227 23072 21272 23100
rect 21085 23063 21143 23069
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 21358 23060 21364 23112
rect 21416 23100 21422 23112
rect 21545 23103 21603 23109
rect 21545 23100 21557 23103
rect 21416 23072 21557 23100
rect 21416 23060 21422 23072
rect 21545 23069 21557 23072
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21634 23060 21640 23112
rect 21692 23100 21698 23112
rect 21818 23100 21824 23112
rect 21692 23072 21824 23100
rect 21692 23060 21698 23072
rect 21818 23060 21824 23072
rect 21876 23060 21882 23112
rect 22186 23060 22192 23112
rect 22244 23100 22250 23112
rect 22579 23100 22607 23140
rect 23106 23128 23112 23140
rect 23164 23128 23170 23180
rect 23658 23128 23664 23180
rect 23716 23168 23722 23180
rect 23716 23140 24992 23168
rect 23716 23128 23722 23140
rect 22244 23072 22607 23100
rect 24029 23103 24087 23109
rect 22244 23060 22250 23072
rect 24029 23069 24041 23103
rect 24075 23100 24087 23103
rect 24118 23100 24124 23112
rect 24075 23072 24124 23100
rect 24075 23069 24087 23072
rect 24029 23063 24087 23069
rect 24118 23060 24124 23072
rect 24176 23060 24182 23112
rect 24964 23086 24992 23140
rect 25038 23128 25044 23180
rect 25096 23168 25102 23180
rect 28721 23171 28779 23177
rect 28721 23168 28733 23171
rect 25096 23140 28733 23168
rect 25096 23128 25102 23140
rect 28721 23137 28733 23140
rect 28767 23137 28779 23171
rect 29270 23168 29276 23180
rect 28721 23131 28779 23137
rect 28920 23140 29276 23168
rect 26326 23060 26332 23112
rect 26384 23100 26390 23112
rect 26384 23072 26429 23100
rect 26384 23060 26390 23072
rect 26694 23060 26700 23112
rect 26752 23100 26758 23112
rect 26881 23103 26939 23109
rect 26881 23100 26893 23103
rect 26752 23072 26893 23100
rect 26752 23060 26758 23072
rect 26881 23069 26893 23072
rect 26927 23069 26939 23103
rect 27062 23100 27068 23112
rect 27023 23072 27068 23100
rect 26881 23063 26939 23069
rect 27062 23060 27068 23072
rect 27120 23060 27126 23112
rect 27614 23100 27620 23112
rect 27575 23072 27620 23100
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 27706 23060 27712 23112
rect 27764 23100 27770 23112
rect 28810 23100 28816 23112
rect 27764 23072 28816 23100
rect 27764 23060 27770 23072
rect 28810 23060 28816 23072
rect 28868 23060 28874 23112
rect 28920 23109 28948 23140
rect 29270 23128 29276 23140
rect 29328 23128 29334 23180
rect 29730 23168 29736 23180
rect 29691 23140 29736 23168
rect 29730 23128 29736 23140
rect 29788 23128 29794 23180
rect 28905 23103 28963 23109
rect 28905 23069 28917 23103
rect 28951 23069 28963 23103
rect 28905 23063 28963 23069
rect 29089 23103 29147 23109
rect 29089 23069 29101 23103
rect 29135 23100 29147 23103
rect 29546 23100 29552 23112
rect 29135 23072 29552 23100
rect 29135 23069 29147 23072
rect 29089 23063 29147 23069
rect 29546 23060 29552 23072
rect 29604 23060 29610 23112
rect 29638 23060 29644 23112
rect 29696 23100 29702 23112
rect 30116 23109 30144 23264
rect 30208 23236 30236 23264
rect 31110 23236 31116 23248
rect 30208 23208 31116 23236
rect 30208 23109 30236 23208
rect 31110 23196 31116 23208
rect 31168 23196 31174 23248
rect 30282 23128 30288 23180
rect 30340 23168 30346 23180
rect 30340 23140 30420 23168
rect 30340 23128 30346 23140
rect 30392 23109 30420 23140
rect 31018 23128 31024 23180
rect 31076 23168 31082 23180
rect 31297 23171 31355 23177
rect 31297 23168 31309 23171
rect 31076 23140 31309 23168
rect 31076 23128 31082 23140
rect 31297 23137 31309 23140
rect 31343 23137 31355 23171
rect 31297 23131 31355 23137
rect 30009 23103 30067 23109
rect 30009 23100 30021 23103
rect 29696 23072 30021 23100
rect 29696 23060 29702 23072
rect 30009 23069 30021 23072
rect 30055 23069 30067 23103
rect 30009 23063 30067 23069
rect 30098 23103 30156 23109
rect 30098 23069 30110 23103
rect 30144 23069 30156 23103
rect 30098 23063 30156 23069
rect 30193 23103 30251 23109
rect 30193 23069 30205 23103
rect 30239 23069 30251 23103
rect 30193 23063 30251 23069
rect 30377 23103 30435 23109
rect 30377 23069 30389 23103
rect 30423 23069 30435 23103
rect 30377 23063 30435 23069
rect 30837 23103 30895 23109
rect 30837 23069 30849 23103
rect 30883 23100 30895 23103
rect 30926 23100 30932 23112
rect 30883 23072 30932 23100
rect 30883 23069 30895 23072
rect 30837 23063 30895 23069
rect 20993 23035 21051 23041
rect 20993 23001 21005 23035
rect 21039 23032 21051 23035
rect 21450 23032 21456 23044
rect 21039 23004 21456 23032
rect 21039 23001 21051 23004
rect 20993 22995 21051 23001
rect 21450 22992 21456 23004
rect 21508 22992 21514 23044
rect 22094 22992 22100 23044
rect 22152 23032 22158 23044
rect 23753 23035 23811 23041
rect 22152 23004 22586 23032
rect 22152 22992 22158 23004
rect 23753 23001 23765 23035
rect 23799 23032 23811 23035
rect 24670 23032 24676 23044
rect 23799 23004 24676 23032
rect 23799 23001 23811 23004
rect 23753 22995 23811 23001
rect 24670 22992 24676 23004
rect 24728 22992 24734 23044
rect 26050 23032 26056 23044
rect 26011 23004 26056 23032
rect 26050 22992 26056 23004
rect 26108 22992 26114 23044
rect 30282 23032 30288 23044
rect 26159 23004 30288 23032
rect 16816 22936 20300 22964
rect 20533 22967 20591 22973
rect 16816 22924 16822 22936
rect 20533 22933 20545 22967
rect 20579 22964 20591 22967
rect 20622 22964 20628 22976
rect 20579 22936 20628 22964
rect 20579 22933 20591 22936
rect 20533 22927 20591 22933
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 21082 22924 21088 22976
rect 21140 22964 21146 22976
rect 24026 22964 24032 22976
rect 21140 22936 24032 22964
rect 21140 22924 21146 22936
rect 24026 22924 24032 22936
rect 24084 22924 24090 22976
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22964 24639 22967
rect 25406 22964 25412 22976
rect 24627 22936 25412 22964
rect 24627 22933 24639 22936
rect 24581 22927 24639 22933
rect 25406 22924 25412 22936
rect 25464 22924 25470 22976
rect 25682 22924 25688 22976
rect 25740 22964 25746 22976
rect 26159 22964 26187 23004
rect 30282 22992 30288 23004
rect 30340 22992 30346 23044
rect 30392 23032 30420 23063
rect 30926 23060 30932 23072
rect 30984 23060 30990 23112
rect 31113 23103 31171 23109
rect 31113 23069 31125 23103
rect 31159 23100 31171 23103
rect 32766 23100 32772 23112
rect 31159 23072 32772 23100
rect 31159 23069 31171 23072
rect 31113 23063 31171 23069
rect 32766 23060 32772 23072
rect 32824 23060 32830 23112
rect 31018 23032 31024 23044
rect 30392 23004 31024 23032
rect 31018 22992 31024 23004
rect 31076 22992 31082 23044
rect 25740 22936 26187 22964
rect 25740 22924 25746 22936
rect 26418 22924 26424 22976
rect 26476 22964 26482 22976
rect 27062 22964 27068 22976
rect 26476 22936 27068 22964
rect 26476 22924 26482 22936
rect 27062 22924 27068 22936
rect 27120 22924 27126 22976
rect 27246 22924 27252 22976
rect 27304 22964 27310 22976
rect 30742 22964 30748 22976
rect 27304 22936 30748 22964
rect 27304 22924 27310 22936
rect 30742 22924 30748 22936
rect 30800 22924 30806 22976
rect 30929 22967 30987 22973
rect 30929 22933 30941 22967
rect 30975 22964 30987 22967
rect 31478 22964 31484 22976
rect 30975 22936 31484 22964
rect 30975 22933 30987 22936
rect 30929 22927 30987 22933
rect 31478 22924 31484 22936
rect 31536 22924 31542 22976
rect 1104 22874 31992 22896
rect 1104 22822 8632 22874
rect 8684 22822 8696 22874
rect 8748 22822 8760 22874
rect 8812 22822 8824 22874
rect 8876 22822 8888 22874
rect 8940 22822 16314 22874
rect 16366 22822 16378 22874
rect 16430 22822 16442 22874
rect 16494 22822 16506 22874
rect 16558 22822 16570 22874
rect 16622 22822 23996 22874
rect 24048 22822 24060 22874
rect 24112 22822 24124 22874
rect 24176 22822 24188 22874
rect 24240 22822 24252 22874
rect 24304 22822 31678 22874
rect 31730 22822 31742 22874
rect 31794 22822 31806 22874
rect 31858 22822 31870 22874
rect 31922 22822 31934 22874
rect 31986 22822 31992 22874
rect 1104 22800 31992 22822
rect 4341 22763 4399 22769
rect 4341 22729 4353 22763
rect 4387 22760 4399 22763
rect 5626 22760 5632 22772
rect 4387 22732 5632 22760
rect 4387 22729 4399 22732
rect 4341 22723 4399 22729
rect 5626 22720 5632 22732
rect 5684 22720 5690 22772
rect 7098 22760 7104 22772
rect 7059 22732 7104 22760
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 8202 22760 8208 22772
rect 8163 22732 8208 22760
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 11149 22763 11207 22769
rect 11149 22729 11161 22763
rect 11195 22760 11207 22763
rect 11974 22760 11980 22772
rect 11195 22732 11980 22760
rect 11195 22729 11207 22732
rect 11149 22723 11207 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12342 22720 12348 22772
rect 12400 22760 12406 22772
rect 12437 22763 12495 22769
rect 12437 22760 12449 22763
rect 12400 22732 12449 22760
rect 12400 22720 12406 22732
rect 12437 22729 12449 22732
rect 12483 22729 12495 22763
rect 12437 22723 12495 22729
rect 12524 22763 12582 22769
rect 12524 22729 12536 22763
rect 12570 22760 12582 22763
rect 12710 22760 12716 22772
rect 12570 22732 12716 22760
rect 12570 22729 12582 22732
rect 12524 22723 12582 22729
rect 12710 22720 12716 22732
rect 12768 22720 12774 22772
rect 12894 22720 12900 22772
rect 12952 22760 12958 22772
rect 13265 22763 13323 22769
rect 13265 22760 13277 22763
rect 12952 22732 13277 22760
rect 12952 22720 12958 22732
rect 13265 22729 13277 22732
rect 13311 22729 13323 22763
rect 13265 22723 13323 22729
rect 13538 22720 13544 22772
rect 13596 22760 13602 22772
rect 13596 22732 14044 22760
rect 13596 22720 13602 22732
rect 4430 22652 4436 22704
rect 4488 22692 4494 22704
rect 5166 22692 5172 22704
rect 4488 22664 5172 22692
rect 4488 22652 4494 22664
rect 5166 22652 5172 22664
rect 5224 22692 5230 22704
rect 5353 22695 5411 22701
rect 5353 22692 5365 22695
rect 5224 22664 5365 22692
rect 5224 22652 5230 22664
rect 5353 22661 5365 22664
rect 5399 22661 5411 22695
rect 5353 22655 5411 22661
rect 7653 22695 7711 22701
rect 7653 22661 7665 22695
rect 7699 22692 7711 22695
rect 8110 22692 8116 22704
rect 7699 22664 8116 22692
rect 7699 22661 7711 22664
rect 7653 22655 7711 22661
rect 8110 22652 8116 22664
rect 8168 22652 8174 22704
rect 10410 22692 10416 22704
rect 10371 22664 10416 22692
rect 10410 22652 10416 22664
rect 10468 22652 10474 22704
rect 11422 22652 11428 22704
rect 11480 22692 11486 22704
rect 14016 22701 14044 22732
rect 14090 22720 14096 22772
rect 14148 22760 14154 22772
rect 14369 22763 14427 22769
rect 14369 22760 14381 22763
rect 14148 22732 14381 22760
rect 14148 22720 14154 22732
rect 14369 22729 14381 22732
rect 14415 22729 14427 22763
rect 16022 22760 16028 22772
rect 14369 22723 14427 22729
rect 15028 22732 16028 22760
rect 15028 22704 15056 22732
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 16114 22720 16120 22772
rect 16172 22760 16178 22772
rect 16301 22763 16359 22769
rect 16301 22760 16313 22763
rect 16172 22732 16313 22760
rect 16172 22720 16178 22732
rect 16301 22729 16313 22732
rect 16347 22729 16359 22763
rect 16301 22723 16359 22729
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 19702 22760 19708 22772
rect 16632 22732 19708 22760
rect 16632 22720 16638 22732
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 19794 22720 19800 22772
rect 19852 22760 19858 22772
rect 19889 22763 19947 22769
rect 19889 22760 19901 22763
rect 19852 22732 19901 22760
rect 19852 22720 19858 22732
rect 19889 22729 19901 22732
rect 19935 22760 19947 22763
rect 21174 22760 21180 22772
rect 19935 22732 21180 22760
rect 19935 22729 19947 22732
rect 19889 22723 19947 22729
rect 21174 22720 21180 22732
rect 21232 22720 21238 22772
rect 21266 22720 21272 22772
rect 21324 22760 21330 22772
rect 22002 22760 22008 22772
rect 21324 22732 22008 22760
rect 21324 22720 21330 22732
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 22738 22720 22744 22772
rect 22796 22760 22802 22772
rect 22796 22732 29868 22760
rect 22796 22720 22802 22732
rect 12621 22695 12679 22701
rect 12621 22692 12633 22695
rect 11480 22664 12633 22692
rect 11480 22652 11486 22664
rect 12621 22661 12633 22664
rect 12667 22661 12679 22695
rect 14001 22695 14059 22701
rect 12621 22655 12679 22661
rect 12912 22664 13952 22692
rect 12912 22636 12940 22664
rect 10318 22624 10324 22636
rect 10279 22596 10324 22624
rect 10318 22584 10324 22596
rect 10376 22584 10382 22636
rect 10502 22624 10508 22636
rect 10463 22596 10508 22624
rect 10502 22584 10508 22596
rect 10560 22584 10566 22636
rect 10965 22627 11023 22633
rect 10965 22593 10977 22627
rect 11011 22593 11023 22627
rect 10965 22587 11023 22593
rect 11149 22627 11207 22633
rect 11149 22593 11161 22627
rect 11195 22593 11207 22627
rect 11149 22587 11207 22593
rect 5902 22516 5908 22568
rect 5960 22556 5966 22568
rect 5960 22528 9674 22556
rect 5960 22516 5966 22528
rect 4893 22491 4951 22497
rect 4893 22457 4905 22491
rect 4939 22488 4951 22491
rect 5810 22488 5816 22500
rect 4939 22460 5816 22488
rect 4939 22457 4951 22460
rect 4893 22451 4951 22457
rect 5810 22448 5816 22460
rect 5868 22448 5874 22500
rect 6362 22448 6368 22500
rect 6420 22488 6426 22500
rect 9217 22491 9275 22497
rect 9217 22488 9229 22491
rect 6420 22460 9229 22488
rect 6420 22448 6426 22460
rect 9217 22457 9229 22460
rect 9263 22488 9275 22491
rect 9306 22488 9312 22500
rect 9263 22460 9312 22488
rect 9263 22457 9275 22460
rect 9217 22451 9275 22457
rect 9306 22448 9312 22460
rect 9364 22448 9370 22500
rect 5997 22423 6055 22429
rect 5997 22389 6009 22423
rect 6043 22420 6055 22423
rect 6086 22420 6092 22432
rect 6043 22392 6092 22420
rect 6043 22389 6055 22392
rect 5997 22383 6055 22389
rect 6086 22380 6092 22392
rect 6144 22380 6150 22432
rect 8754 22420 8760 22432
rect 8715 22392 8760 22420
rect 8754 22380 8760 22392
rect 8812 22380 8818 22432
rect 9646 22420 9674 22528
rect 9858 22488 9864 22500
rect 9819 22460 9864 22488
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 10980 22488 11008 22587
rect 11164 22556 11192 22587
rect 11606 22584 11612 22636
rect 11664 22624 11670 22636
rect 11701 22627 11759 22633
rect 11701 22624 11713 22627
rect 11664 22596 11713 22624
rect 11664 22584 11670 22596
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 12713 22627 12771 22633
rect 11701 22587 11759 22593
rect 12268 22596 12674 22624
rect 12268 22556 12296 22596
rect 11164 22528 12296 22556
rect 12345 22559 12403 22565
rect 12345 22525 12357 22559
rect 12391 22556 12403 22559
rect 12434 22556 12440 22568
rect 12391 22528 12440 22556
rect 12391 22525 12403 22528
rect 12345 22519 12403 22525
rect 12434 22516 12440 22528
rect 12492 22516 12498 22568
rect 12646 22556 12674 22596
rect 12713 22593 12725 22627
rect 12759 22624 12771 22627
rect 12802 22624 12808 22636
rect 12759 22596 12808 22624
rect 12759 22593 12771 22596
rect 12713 22587 12771 22593
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 12894 22584 12900 22636
rect 12952 22584 12958 22636
rect 13078 22584 13084 22636
rect 13136 22624 13142 22636
rect 13173 22627 13231 22633
rect 13173 22624 13185 22627
rect 13136 22596 13185 22624
rect 13136 22584 13142 22596
rect 13173 22593 13185 22596
rect 13219 22593 13231 22627
rect 13173 22587 13231 22593
rect 13354 22584 13360 22636
rect 13412 22633 13418 22636
rect 13412 22627 13457 22633
rect 13445 22593 13457 22627
rect 13412 22587 13457 22593
rect 13541 22627 13599 22633
rect 13541 22593 13553 22627
rect 13587 22624 13599 22627
rect 13814 22624 13820 22636
rect 13587 22596 13820 22624
rect 13587 22593 13599 22596
rect 13541 22587 13599 22593
rect 13412 22584 13418 22587
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 13924 22624 13952 22664
rect 14001 22661 14013 22695
rect 14047 22692 14059 22695
rect 14642 22692 14648 22704
rect 14047 22664 14648 22692
rect 14047 22661 14059 22664
rect 14001 22655 14059 22661
rect 14642 22652 14648 22664
rect 14700 22692 14706 22704
rect 14921 22695 14979 22701
rect 14700 22664 14872 22692
rect 14700 22652 14706 22664
rect 14844 22633 14872 22664
rect 14921 22661 14933 22695
rect 14967 22692 14979 22695
rect 15010 22692 15016 22704
rect 14967 22664 15016 22692
rect 14967 22661 14979 22664
rect 14921 22655 14979 22661
rect 15010 22652 15016 22664
rect 15068 22652 15074 22704
rect 15289 22695 15347 22701
rect 15289 22661 15301 22695
rect 15335 22692 15347 22695
rect 15470 22692 15476 22704
rect 15335 22664 15476 22692
rect 15335 22661 15347 22664
rect 15289 22655 15347 22661
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 15838 22652 15844 22704
rect 15896 22692 15902 22704
rect 16850 22692 16856 22704
rect 15896 22664 16856 22692
rect 15896 22652 15902 22664
rect 16850 22652 16856 22664
rect 16908 22652 16914 22704
rect 17402 22652 17408 22704
rect 17460 22692 17466 22704
rect 17862 22692 17868 22704
rect 17460 22664 17868 22692
rect 17460 22652 17466 22664
rect 17862 22652 17868 22664
rect 17920 22652 17926 22704
rect 18138 22652 18144 22704
rect 18196 22692 18202 22704
rect 18509 22695 18567 22701
rect 18509 22692 18521 22695
rect 18196 22664 18521 22692
rect 18196 22652 18202 22664
rect 18509 22661 18521 22664
rect 18555 22692 18567 22695
rect 20346 22692 20352 22704
rect 18555 22664 20352 22692
rect 18555 22661 18567 22664
rect 18509 22655 18567 22661
rect 20346 22652 20352 22664
rect 20404 22652 20410 22704
rect 21542 22652 21548 22704
rect 21600 22692 21606 22704
rect 21600 22664 23060 22692
rect 21600 22652 21606 22664
rect 20720 22636 20772 22642
rect 14185 22627 14243 22633
rect 14185 22624 14197 22627
rect 13924 22596 14197 22624
rect 14185 22593 14197 22596
rect 14231 22593 14243 22627
rect 14185 22587 14243 22593
rect 14829 22627 14887 22633
rect 14829 22593 14841 22627
rect 14875 22593 14887 22627
rect 15102 22624 15108 22636
rect 15063 22596 15108 22624
rect 14829 22587 14887 22593
rect 15102 22584 15108 22596
rect 15160 22584 15166 22636
rect 15933 22627 15991 22633
rect 15933 22624 15945 22627
rect 15488 22596 15945 22624
rect 13906 22556 13912 22568
rect 12646 22528 13912 22556
rect 13906 22516 13912 22528
rect 13964 22556 13970 22568
rect 13964 22528 14044 22556
rect 13964 22516 13970 22528
rect 11793 22491 11851 22497
rect 10980 22460 11744 22488
rect 10778 22420 10784 22432
rect 9646 22392 10784 22420
rect 10778 22380 10784 22392
rect 10836 22420 10842 22432
rect 11054 22420 11060 22432
rect 10836 22392 11060 22420
rect 10836 22380 10842 22392
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 11716 22420 11744 22460
rect 11793 22457 11805 22491
rect 11839 22488 11851 22491
rect 13262 22488 13268 22500
rect 11839 22460 13268 22488
rect 11839 22457 11851 22460
rect 11793 22451 11851 22457
rect 13262 22448 13268 22460
rect 13320 22448 13326 22500
rect 14016 22488 14044 22528
rect 14090 22516 14096 22568
rect 14148 22556 14154 22568
rect 15488 22556 15516 22596
rect 15933 22593 15945 22596
rect 15979 22593 15991 22627
rect 15933 22587 15991 22593
rect 16298 22584 16304 22636
rect 16356 22624 16362 22636
rect 16758 22624 16764 22636
rect 16356 22596 16764 22624
rect 16356 22584 16362 22596
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 17313 22627 17371 22633
rect 17313 22593 17325 22627
rect 17359 22624 17371 22627
rect 17586 22624 17592 22636
rect 17359 22596 17592 22624
rect 17359 22593 17371 22596
rect 17313 22587 17371 22593
rect 17586 22584 17592 22596
rect 17644 22584 17650 22636
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 18325 22627 18383 22633
rect 18325 22624 18337 22627
rect 18288 22596 18337 22624
rect 18288 22584 18294 22596
rect 18325 22593 18337 22596
rect 18371 22593 18383 22627
rect 18325 22587 18383 22593
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18690 22624 18696 22636
rect 18651 22596 18696 22624
rect 18417 22587 18475 22593
rect 14148 22528 15516 22556
rect 14148 22516 14154 22528
rect 15562 22516 15568 22568
rect 15620 22556 15626 22568
rect 15841 22559 15899 22565
rect 15841 22556 15853 22559
rect 15620 22528 15853 22556
rect 15620 22516 15626 22528
rect 15841 22525 15853 22528
rect 15887 22525 15899 22559
rect 15841 22519 15899 22525
rect 16022 22516 16028 22568
rect 16080 22556 16086 22568
rect 17221 22559 17279 22565
rect 17221 22556 17233 22559
rect 16080 22528 17233 22556
rect 16080 22516 16086 22528
rect 17221 22525 17233 22528
rect 17267 22556 17279 22559
rect 17267 22528 17632 22556
rect 17267 22525 17279 22528
rect 17221 22519 17279 22525
rect 15010 22488 15016 22500
rect 14016 22460 15016 22488
rect 15010 22448 15016 22460
rect 15068 22448 15074 22500
rect 16206 22448 16212 22500
rect 16264 22488 16270 22500
rect 16482 22488 16488 22500
rect 16264 22460 16488 22488
rect 16264 22448 16270 22460
rect 16482 22448 16488 22460
rect 16540 22448 16546 22500
rect 16758 22448 16764 22500
rect 16816 22488 16822 22500
rect 16942 22488 16948 22500
rect 16816 22460 16948 22488
rect 16816 22448 16822 22460
rect 16942 22448 16948 22460
rect 17000 22448 17006 22500
rect 17034 22448 17040 22500
rect 17092 22488 17098 22500
rect 17310 22488 17316 22500
rect 17092 22460 17316 22488
rect 17092 22448 17098 22460
rect 17310 22448 17316 22460
rect 17368 22448 17374 22500
rect 12342 22420 12348 22432
rect 11716 22392 12348 22420
rect 12342 22380 12348 22392
rect 12400 22420 12406 22432
rect 12710 22420 12716 22432
rect 12400 22392 12716 22420
rect 12400 22380 12406 22392
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 13541 22423 13599 22429
rect 13541 22389 13553 22423
rect 13587 22420 13599 22423
rect 17402 22420 17408 22432
rect 13587 22392 17408 22420
rect 13587 22389 13599 22392
rect 13541 22383 13599 22389
rect 17402 22380 17408 22392
rect 17460 22380 17466 22432
rect 17604 22420 17632 22528
rect 17770 22516 17776 22568
rect 17828 22556 17834 22568
rect 18432 22556 18460 22587
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 18782 22584 18788 22636
rect 18840 22624 18846 22636
rect 18840 22596 18885 22624
rect 18840 22584 18846 22596
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19024 22596 19625 22624
rect 19024 22584 19030 22596
rect 19613 22593 19625 22596
rect 19659 22593 19671 22627
rect 19613 22587 19671 22593
rect 19730 22627 19788 22633
rect 19730 22593 19742 22627
rect 19776 22624 19788 22627
rect 19978 22624 19984 22636
rect 19776 22596 19984 22624
rect 19776 22593 19788 22596
rect 19730 22587 19788 22593
rect 19242 22556 19248 22568
rect 17828 22528 18460 22556
rect 19203 22528 19248 22556
rect 17828 22516 17834 22528
rect 19242 22516 19248 22528
rect 19300 22516 19306 22568
rect 19518 22556 19524 22568
rect 19479 22528 19524 22556
rect 19518 22516 19524 22528
rect 19576 22516 19582 22568
rect 19628 22556 19656 22587
rect 19978 22584 19984 22596
rect 20036 22584 20042 22636
rect 21361 22627 21419 22633
rect 20772 22586 20852 22614
rect 21361 22593 21373 22627
rect 21407 22624 21419 22627
rect 21910 22624 21916 22636
rect 21407 22596 21916 22624
rect 21407 22593 21419 22596
rect 21361 22587 21419 22593
rect 20720 22578 20772 22584
rect 20824 22556 20852 22586
rect 21910 22584 21916 22596
rect 21968 22584 21974 22636
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22624 22247 22627
rect 22646 22624 22652 22636
rect 22235 22596 22652 22624
rect 22235 22593 22247 22596
rect 22189 22587 22247 22593
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 21542 22556 21548 22568
rect 19628 22528 20668 22556
rect 20824 22528 21548 22556
rect 17681 22491 17739 22497
rect 17681 22457 17693 22491
rect 17727 22488 17739 22491
rect 17954 22488 17960 22500
rect 17727 22460 17960 22488
rect 17727 22457 17739 22460
rect 17681 22451 17739 22457
rect 17954 22448 17960 22460
rect 18012 22448 18018 22500
rect 18141 22491 18199 22497
rect 18141 22457 18153 22491
rect 18187 22488 18199 22491
rect 18506 22488 18512 22500
rect 18187 22460 18512 22488
rect 18187 22457 18199 22460
rect 18141 22451 18199 22457
rect 18506 22448 18512 22460
rect 18564 22448 18570 22500
rect 19334 22448 19340 22500
rect 19392 22488 19398 22500
rect 19978 22488 19984 22500
rect 19392 22460 19984 22488
rect 19392 22448 19398 22460
rect 19978 22448 19984 22460
rect 20036 22448 20042 22500
rect 19518 22420 19524 22432
rect 17604 22392 19524 22420
rect 19518 22380 19524 22392
rect 19576 22420 19582 22432
rect 20070 22420 20076 22432
rect 19576 22392 20076 22420
rect 19576 22380 19582 22392
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 20640 22420 20668 22528
rect 21542 22516 21548 22528
rect 21600 22516 21606 22568
rect 21634 22516 21640 22568
rect 21692 22556 21698 22568
rect 22370 22556 22376 22568
rect 21692 22528 22376 22556
rect 21692 22516 21698 22528
rect 22370 22516 22376 22528
rect 22428 22516 22434 22568
rect 22465 22559 22523 22565
rect 22465 22525 22477 22559
rect 22511 22556 22523 22559
rect 22738 22556 22744 22568
rect 22511 22528 22744 22556
rect 22511 22525 22523 22528
rect 22465 22519 22523 22525
rect 22738 22516 22744 22528
rect 22796 22516 22802 22568
rect 22922 22556 22928 22568
rect 22883 22528 22928 22556
rect 22922 22516 22928 22528
rect 22980 22516 22986 22568
rect 23032 22556 23060 22664
rect 25314 22652 25320 22704
rect 25372 22652 25378 22704
rect 25958 22652 25964 22704
rect 26016 22692 26022 22704
rect 29638 22692 29644 22704
rect 26016 22664 29644 22692
rect 26016 22652 26022 22664
rect 29638 22652 29644 22664
rect 29696 22652 29702 22704
rect 23750 22624 23756 22636
rect 23711 22596 23756 22624
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22624 23995 22627
rect 24578 22624 24584 22636
rect 23983 22596 24584 22624
rect 23983 22593 23995 22596
rect 23937 22587 23995 22593
rect 24578 22584 24584 22596
rect 24636 22584 24642 22636
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 26384 22596 26429 22624
rect 26384 22584 26390 22596
rect 26510 22584 26516 22636
rect 26568 22624 26574 22636
rect 26970 22624 26976 22636
rect 26568 22596 26976 22624
rect 26568 22584 26574 22596
rect 26970 22584 26976 22596
rect 27028 22624 27034 22636
rect 27246 22633 27252 22636
rect 27225 22627 27252 22633
rect 27028 22596 27187 22624
rect 27028 22584 27034 22596
rect 25958 22556 25964 22568
rect 23032 22528 25964 22556
rect 25958 22516 25964 22528
rect 26016 22516 26022 22568
rect 26053 22559 26111 22565
rect 26053 22525 26065 22559
rect 26099 22556 26111 22559
rect 26099 22528 26390 22556
rect 26099 22525 26111 22528
rect 26053 22519 26111 22525
rect 21082 22448 21088 22500
rect 21140 22488 21146 22500
rect 21140 22460 21588 22488
rect 21140 22448 21146 22460
rect 21174 22420 21180 22432
rect 20640 22392 21180 22420
rect 21174 22380 21180 22392
rect 21232 22380 21238 22432
rect 21560 22420 21588 22460
rect 21818 22448 21824 22500
rect 21876 22488 21882 22500
rect 23658 22488 23664 22500
rect 21876 22460 23664 22488
rect 21876 22448 21882 22460
rect 23658 22448 23664 22460
rect 23716 22448 23722 22500
rect 24581 22491 24639 22497
rect 24581 22457 24593 22491
rect 24627 22488 24639 22491
rect 24854 22488 24860 22500
rect 24627 22460 24860 22488
rect 24627 22457 24639 22460
rect 24581 22451 24639 22457
rect 24854 22448 24860 22460
rect 24912 22448 24918 22500
rect 26362 22488 26390 22528
rect 26418 22516 26424 22568
rect 26476 22556 26482 22568
rect 27159 22556 27187 22596
rect 27225 22593 27237 22627
rect 27225 22587 27252 22593
rect 27246 22584 27252 22587
rect 27304 22584 27310 22636
rect 27614 22624 27620 22636
rect 27575 22596 27620 22624
rect 27614 22584 27620 22596
rect 27672 22624 27678 22636
rect 28258 22624 28264 22636
rect 27672 22596 28264 22624
rect 27672 22584 27678 22596
rect 28258 22584 28264 22596
rect 28316 22584 28322 22636
rect 28353 22627 28411 22633
rect 28353 22593 28365 22627
rect 28399 22593 28411 22627
rect 28353 22587 28411 22593
rect 27433 22559 27491 22565
rect 27433 22556 27445 22559
rect 26476 22528 26648 22556
rect 27159 22528 27445 22556
rect 26476 22516 26482 22528
rect 26620 22488 26648 22528
rect 27433 22525 27445 22528
rect 27479 22525 27491 22559
rect 27433 22519 27491 22525
rect 28074 22516 28080 22568
rect 28132 22556 28138 22568
rect 28368 22556 28396 22587
rect 28442 22584 28448 22636
rect 28500 22624 28506 22636
rect 28629 22627 28687 22633
rect 28629 22624 28641 22627
rect 28500 22596 28641 22624
rect 28500 22584 28506 22596
rect 28629 22593 28641 22596
rect 28675 22593 28687 22627
rect 29089 22627 29147 22633
rect 28748 22622 28994 22626
rect 28629 22587 28687 22593
rect 28736 22598 28994 22622
rect 28736 22594 28776 22598
rect 28736 22556 28764 22594
rect 28132 22528 28396 22556
rect 28460 22528 28764 22556
rect 28966 22556 28994 22598
rect 29089 22593 29101 22627
rect 29135 22624 29147 22627
rect 29178 22624 29184 22636
rect 29135 22596 29184 22624
rect 29135 22593 29147 22596
rect 29089 22587 29147 22593
rect 29178 22584 29184 22596
rect 29236 22584 29242 22636
rect 29546 22624 29552 22636
rect 29507 22596 29552 22624
rect 29546 22584 29552 22596
rect 29604 22584 29610 22636
rect 29733 22627 29791 22633
rect 29733 22593 29745 22627
rect 29779 22593 29791 22627
rect 29840 22624 29868 22732
rect 30282 22720 30288 22772
rect 30340 22760 30346 22772
rect 30929 22763 30987 22769
rect 30929 22760 30941 22763
rect 30340 22732 30941 22760
rect 30340 22720 30346 22732
rect 30929 22729 30941 22732
rect 30975 22729 30987 22763
rect 30929 22723 30987 22729
rect 31018 22720 31024 22772
rect 31076 22760 31082 22772
rect 31076 22732 31121 22760
rect 31076 22720 31082 22732
rect 31110 22692 31116 22704
rect 31071 22664 31116 22692
rect 31110 22652 31116 22664
rect 31168 22652 31174 22704
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 29840 22596 29929 22624
rect 29733 22587 29791 22593
rect 29917 22593 29929 22596
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 30101 22627 30159 22633
rect 30101 22593 30113 22627
rect 30147 22624 30159 22627
rect 30374 22624 30380 22636
rect 30147 22596 30380 22624
rect 30147 22593 30159 22596
rect 30101 22587 30159 22593
rect 29748 22556 29776 22587
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 30926 22584 30932 22636
rect 30984 22624 30990 22636
rect 32858 22624 32864 22636
rect 30984 22596 32864 22624
rect 30984 22584 30990 22596
rect 32858 22584 32864 22596
rect 32916 22584 32922 22636
rect 28966 22528 29776 22556
rect 28132 22516 28138 22528
rect 28460 22488 28488 22528
rect 29822 22516 29828 22568
rect 29880 22556 29886 22568
rect 30742 22556 30748 22568
rect 29880 22528 29925 22556
rect 30703 22528 30748 22556
rect 29880 22516 29886 22528
rect 30742 22516 30748 22528
rect 30800 22516 30806 22568
rect 30834 22516 30840 22568
rect 30892 22556 30898 22568
rect 32674 22556 32680 22568
rect 30892 22528 32680 22556
rect 30892 22516 30898 22528
rect 32674 22516 32680 22528
rect 32732 22516 32738 22568
rect 28718 22488 28724 22500
rect 26362 22460 26556 22488
rect 26620 22460 28488 22488
rect 28679 22460 28724 22488
rect 22005 22423 22063 22429
rect 22005 22420 22017 22423
rect 21560 22392 22017 22420
rect 22005 22389 22017 22392
rect 22051 22389 22063 22423
rect 22005 22383 22063 22389
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 22373 22423 22431 22429
rect 22373 22420 22385 22423
rect 22244 22392 22385 22420
rect 22244 22380 22250 22392
rect 22373 22389 22385 22392
rect 22419 22389 22431 22423
rect 22373 22383 22431 22389
rect 22462 22380 22468 22432
rect 22520 22420 22526 22432
rect 23106 22420 23112 22432
rect 22520 22392 23112 22420
rect 22520 22380 22526 22392
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 23934 22380 23940 22432
rect 23992 22420 23998 22432
rect 26418 22420 26424 22432
rect 23992 22392 26424 22420
rect 23992 22380 23998 22392
rect 26418 22380 26424 22392
rect 26476 22380 26482 22432
rect 26528 22420 26556 22460
rect 28718 22448 28724 22460
rect 28776 22448 28782 22500
rect 28813 22491 28871 22497
rect 28813 22457 28825 22491
rect 28859 22488 28871 22491
rect 29270 22488 29276 22500
rect 28859 22460 29276 22488
rect 28859 22457 28871 22460
rect 28813 22451 28871 22457
rect 29270 22448 29276 22460
rect 29328 22448 29334 22500
rect 29638 22448 29644 22500
rect 29696 22488 29702 22500
rect 31297 22491 31355 22497
rect 31297 22488 31309 22491
rect 29696 22460 31309 22488
rect 29696 22448 29702 22460
rect 31297 22457 31309 22460
rect 31343 22457 31355 22491
rect 31297 22451 31355 22457
rect 26694 22420 26700 22432
rect 26528 22392 26700 22420
rect 26694 22380 26700 22392
rect 26752 22380 26758 22432
rect 27246 22380 27252 22432
rect 27304 22420 27310 22432
rect 27341 22423 27399 22429
rect 27341 22420 27353 22423
rect 27304 22392 27353 22420
rect 27304 22380 27310 22392
rect 27341 22389 27353 22392
rect 27387 22389 27399 22423
rect 27522 22420 27528 22432
rect 27483 22392 27528 22420
rect 27341 22383 27399 22389
rect 27522 22380 27528 22392
rect 27580 22380 27586 22432
rect 27893 22423 27951 22429
rect 27893 22389 27905 22423
rect 27939 22420 27951 22423
rect 28626 22420 28632 22432
rect 27939 22392 28632 22420
rect 27939 22389 27951 22392
rect 27893 22383 27951 22389
rect 28626 22380 28632 22392
rect 28684 22380 28690 22432
rect 28905 22423 28963 22429
rect 28905 22389 28917 22423
rect 28951 22420 28963 22423
rect 28994 22420 29000 22432
rect 28951 22392 29000 22420
rect 28951 22389 28963 22392
rect 28905 22383 28963 22389
rect 28994 22380 29000 22392
rect 29052 22420 29058 22432
rect 30098 22420 30104 22432
rect 29052 22392 30104 22420
rect 29052 22380 29058 22392
rect 30098 22380 30104 22392
rect 30156 22380 30162 22432
rect 30282 22420 30288 22432
rect 30243 22392 30288 22420
rect 30282 22380 30288 22392
rect 30340 22380 30346 22432
rect 30742 22380 30748 22432
rect 30800 22420 30806 22432
rect 32122 22420 32128 22432
rect 30800 22392 32128 22420
rect 30800 22380 30806 22392
rect 32122 22380 32128 22392
rect 32180 22380 32186 22432
rect 1104 22330 31832 22352
rect 1104 22278 4791 22330
rect 4843 22278 4855 22330
rect 4907 22278 4919 22330
rect 4971 22278 4983 22330
rect 5035 22278 5047 22330
rect 5099 22278 12473 22330
rect 12525 22278 12537 22330
rect 12589 22278 12601 22330
rect 12653 22278 12665 22330
rect 12717 22278 12729 22330
rect 12781 22278 20155 22330
rect 20207 22278 20219 22330
rect 20271 22278 20283 22330
rect 20335 22278 20347 22330
rect 20399 22278 20411 22330
rect 20463 22278 27837 22330
rect 27889 22278 27901 22330
rect 27953 22278 27965 22330
rect 28017 22278 28029 22330
rect 28081 22278 28093 22330
rect 28145 22278 31832 22330
rect 1104 22256 31832 22278
rect 5534 22176 5540 22228
rect 5592 22216 5598 22228
rect 5813 22219 5871 22225
rect 5813 22216 5825 22219
rect 5592 22188 5825 22216
rect 5592 22176 5598 22188
rect 5813 22185 5825 22188
rect 5859 22216 5871 22219
rect 5902 22216 5908 22228
rect 5859 22188 5908 22216
rect 5859 22185 5871 22188
rect 5813 22179 5871 22185
rect 5902 22176 5908 22188
rect 5960 22176 5966 22228
rect 6362 22216 6368 22228
rect 6323 22188 6368 22216
rect 6362 22176 6368 22188
rect 6420 22176 6426 22228
rect 6546 22176 6552 22228
rect 6604 22216 6610 22228
rect 9582 22216 9588 22228
rect 6604 22188 9588 22216
rect 6604 22176 6610 22188
rect 9582 22176 9588 22188
rect 9640 22216 9646 22228
rect 9766 22216 9772 22228
rect 9640 22188 9772 22216
rect 9640 22176 9646 22188
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 11146 22216 11152 22228
rect 10888 22188 11152 22216
rect 9677 22151 9735 22157
rect 9677 22117 9689 22151
rect 9723 22148 9735 22151
rect 10888 22148 10916 22188
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 11974 22216 11980 22228
rect 11935 22188 11980 22216
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 14090 22216 14096 22228
rect 12176 22188 14096 22216
rect 11054 22148 11060 22160
rect 9723 22120 10916 22148
rect 11015 22120 11060 22148
rect 9723 22117 9735 22120
rect 9677 22111 9735 22117
rect 5261 22083 5319 22089
rect 5261 22049 5273 22083
rect 5307 22080 5319 22083
rect 5350 22080 5356 22092
rect 5307 22052 5356 22080
rect 5307 22049 5319 22052
rect 5261 22043 5319 22049
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 10778 22080 10784 22092
rect 9364 22052 10784 22080
rect 9364 22040 9370 22052
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 10888 22089 10916 22120
rect 11054 22108 11060 22120
rect 11112 22148 11118 22160
rect 12176 22148 12204 22188
rect 14090 22176 14096 22188
rect 14148 22176 14154 22228
rect 14274 22216 14280 22228
rect 14235 22188 14280 22216
rect 14274 22176 14280 22188
rect 14332 22176 14338 22228
rect 14458 22216 14464 22228
rect 14419 22188 14464 22216
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 17126 22216 17132 22228
rect 15166 22188 17132 22216
rect 13078 22148 13084 22160
rect 11112 22120 12204 22148
rect 12268 22120 13084 22148
rect 11112 22108 11118 22120
rect 10873 22083 10931 22089
rect 10873 22049 10885 22083
rect 10919 22049 10931 22083
rect 12268 22080 12296 22120
rect 13078 22108 13084 22120
rect 13136 22108 13142 22160
rect 15166 22148 15194 22188
rect 17126 22176 17132 22188
rect 17184 22176 17190 22228
rect 19150 22216 19156 22228
rect 17328 22188 19156 22216
rect 16574 22148 16580 22160
rect 13740 22120 15194 22148
rect 15228 22120 16580 22148
rect 10873 22043 10931 22049
rect 10980 22052 12296 22080
rect 4706 22012 4712 22024
rect 4667 21984 4712 22012
rect 4706 21972 4712 21984
rect 4764 21972 4770 22024
rect 9582 22012 9588 22024
rect 6932 21984 9444 22012
rect 9543 21984 9588 22012
rect 4246 21904 4252 21956
rect 4304 21944 4310 21956
rect 6932 21953 6960 21984
rect 6917 21947 6975 21953
rect 6917 21944 6929 21947
rect 4304 21916 6929 21944
rect 4304 21904 4310 21916
rect 6917 21913 6929 21916
rect 6963 21913 6975 21947
rect 6917 21907 6975 21913
rect 8021 21947 8079 21953
rect 8021 21913 8033 21947
rect 8067 21944 8079 21947
rect 9122 21944 9128 21956
rect 8067 21916 9128 21944
rect 8067 21913 8079 21916
rect 8021 21907 8079 21913
rect 9122 21904 9128 21916
rect 9180 21904 9186 21956
rect 4157 21879 4215 21885
rect 4157 21845 4169 21879
rect 4203 21876 4215 21879
rect 6546 21876 6552 21888
rect 4203 21848 6552 21876
rect 4203 21845 4215 21848
rect 4157 21839 4215 21845
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 7469 21879 7527 21885
rect 7469 21845 7481 21879
rect 7515 21876 7527 21879
rect 7558 21876 7564 21888
rect 7515 21848 7564 21876
rect 7515 21845 7527 21848
rect 7469 21839 7527 21845
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 8478 21876 8484 21888
rect 8439 21848 8484 21876
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 9416 21876 9444 21984
rect 9582 21972 9588 21984
rect 9640 21972 9646 22024
rect 10226 22012 10232 22024
rect 10187 21984 10232 22012
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10318 21972 10324 22024
rect 10376 22012 10382 22024
rect 10376 21984 10421 22012
rect 10376 21972 10382 21984
rect 9950 21904 9956 21956
rect 10008 21944 10014 21956
rect 10980 21944 11008 22052
rect 11146 22012 11152 22024
rect 11107 21984 11152 22012
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 11808 22021 11836 22052
rect 12342 22040 12348 22092
rect 12400 22080 12406 22092
rect 12805 22083 12863 22089
rect 12400 22052 12756 22080
rect 12400 22040 12406 22052
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11348 21984 11621 22012
rect 11348 21956 11376 21984
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 21981 11851 22015
rect 12437 22015 12495 22021
rect 12437 22012 12449 22015
rect 11793 21975 11851 21981
rect 12176 21984 12449 22012
rect 11330 21944 11336 21956
rect 10008 21916 11008 21944
rect 11072 21916 11336 21944
rect 10008 21904 10014 21916
rect 11072 21876 11100 21916
rect 11330 21904 11336 21916
rect 11388 21904 11394 21956
rect 11422 21904 11428 21956
rect 11480 21944 11486 21956
rect 12176 21944 12204 21984
rect 12437 21981 12449 21984
rect 12483 21981 12495 22015
rect 12618 22012 12624 22024
rect 12579 21984 12624 22012
rect 12437 21975 12495 21981
rect 12618 21972 12624 21984
rect 12676 21972 12682 22024
rect 12728 22012 12756 22052
rect 12805 22049 12817 22083
rect 12851 22080 12863 22083
rect 13630 22080 13636 22092
rect 12851 22052 13636 22080
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 13630 22040 13636 22052
rect 13688 22040 13694 22092
rect 13078 22012 13084 22024
rect 12728 21984 13084 22012
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 13446 22012 13452 22024
rect 13407 21984 13452 22012
rect 13446 21972 13452 21984
rect 13504 21972 13510 22024
rect 13740 22021 13768 22120
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 15228 21956 15256 22120
rect 16574 22108 16580 22120
rect 16632 22108 16638 22160
rect 16669 22151 16727 22157
rect 16669 22117 16681 22151
rect 16715 22148 16727 22151
rect 17328 22148 17356 22188
rect 19150 22176 19156 22188
rect 19208 22176 19214 22228
rect 20714 22216 20720 22228
rect 19260 22188 20720 22216
rect 16715 22120 17356 22148
rect 16715 22117 16727 22120
rect 16669 22111 16727 22117
rect 17402 22108 17408 22160
rect 17460 22148 17466 22160
rect 18046 22148 18052 22160
rect 17460 22120 18052 22148
rect 17460 22108 17466 22120
rect 18046 22108 18052 22120
rect 18104 22108 18110 22160
rect 18322 22108 18328 22160
rect 18380 22108 18386 22160
rect 18414 22108 18420 22160
rect 18472 22148 18478 22160
rect 19260 22148 19288 22188
rect 20714 22176 20720 22188
rect 20772 22176 20778 22228
rect 20990 22176 20996 22228
rect 21048 22216 21054 22228
rect 23397 22219 23455 22225
rect 23397 22216 23409 22219
rect 21048 22188 23409 22216
rect 21048 22176 21054 22188
rect 23397 22185 23409 22188
rect 23443 22185 23455 22219
rect 23397 22179 23455 22185
rect 23658 22176 23664 22228
rect 23716 22216 23722 22228
rect 24670 22216 24676 22228
rect 23716 22188 24676 22216
rect 23716 22176 23722 22188
rect 24670 22176 24676 22188
rect 24728 22176 24734 22228
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 25774 22216 25780 22228
rect 25188 22188 25780 22216
rect 25188 22176 25194 22188
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 26142 22176 26148 22228
rect 26200 22216 26206 22228
rect 26694 22216 26700 22228
rect 26200 22188 26700 22216
rect 26200 22176 26206 22188
rect 26694 22176 26700 22188
rect 26752 22176 26758 22228
rect 26970 22176 26976 22228
rect 27028 22216 27034 22228
rect 28442 22216 28448 22228
rect 27028 22188 28448 22216
rect 27028 22176 27034 22188
rect 28442 22176 28448 22188
rect 28500 22176 28506 22228
rect 28626 22176 28632 22228
rect 28684 22216 28690 22228
rect 29086 22216 29092 22228
rect 28684 22188 28994 22216
rect 29047 22188 29092 22216
rect 28684 22176 28690 22188
rect 18472 22120 19288 22148
rect 18472 22108 18478 22120
rect 15381 22083 15439 22089
rect 15381 22049 15393 22083
rect 15427 22080 15439 22083
rect 15654 22080 15660 22092
rect 15427 22052 15516 22080
rect 15615 22052 15660 22080
rect 15427 22049 15439 22052
rect 15381 22043 15439 22049
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 22012 15347 22015
rect 15488 22012 15516 22052
rect 15654 22040 15660 22052
rect 15712 22040 15718 22092
rect 16114 22040 16120 22092
rect 16172 22080 16178 22092
rect 16209 22083 16267 22089
rect 16209 22080 16221 22083
rect 16172 22052 16221 22080
rect 16172 22040 16178 22052
rect 16209 22049 16221 22052
rect 16255 22049 16267 22083
rect 16209 22043 16267 22049
rect 16942 22040 16948 22092
rect 17000 22080 17006 22092
rect 17000 22052 17264 22080
rect 17000 22040 17006 22052
rect 15930 22012 15936 22024
rect 15335 21984 15424 22012
rect 15488 21984 15936 22012
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 15396 21956 15424 21984
rect 15930 21972 15936 21984
rect 15988 21972 15994 22024
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 11480 21916 12204 21944
rect 11480 21904 11486 21916
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 14445 21947 14503 21953
rect 12308 21916 13676 21944
rect 12308 21904 12314 21916
rect 13648 21888 13676 21916
rect 14445 21913 14457 21947
rect 14491 21944 14503 21947
rect 14550 21944 14556 21956
rect 14491 21916 14556 21944
rect 14491 21913 14503 21916
rect 14445 21907 14503 21913
rect 14550 21904 14556 21916
rect 14608 21904 14614 21956
rect 14645 21947 14703 21953
rect 14645 21913 14657 21947
rect 14691 21944 14703 21947
rect 15194 21944 15200 21956
rect 14691 21916 15200 21944
rect 14691 21913 14703 21916
rect 14645 21907 14703 21913
rect 15194 21904 15200 21916
rect 15252 21944 15258 21956
rect 15252 21916 15345 21944
rect 15252 21904 15258 21916
rect 15378 21904 15384 21956
rect 15436 21904 15442 21956
rect 16022 21904 16028 21956
rect 16080 21944 16086 21956
rect 16316 21944 16344 21975
rect 16080 21916 16344 21944
rect 16080 21904 16086 21916
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 17129 21947 17187 21953
rect 17129 21944 17141 21947
rect 16540 21916 17141 21944
rect 16540 21904 16546 21916
rect 17129 21913 17141 21916
rect 17175 21913 17187 21947
rect 17236 21944 17264 22052
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 18340 22080 18368 22108
rect 17368 22052 17632 22080
rect 18340 22052 18552 22080
rect 17368 22040 17374 22052
rect 17402 22012 17408 22024
rect 17363 21984 17408 22012
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 17604 22021 17632 22052
rect 17497 22015 17555 22021
rect 17497 21981 17509 22015
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 21981 17647 22015
rect 17770 22012 17776 22024
rect 17731 21984 17776 22012
rect 17589 21975 17647 21981
rect 17512 21944 17540 21975
rect 17770 21972 17776 21984
rect 17828 21972 17834 22024
rect 18046 22012 18052 22024
rect 17880 21984 18052 22012
rect 17880 21944 17908 21984
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18138 21972 18144 22024
rect 18196 22012 18202 22024
rect 18233 22015 18291 22021
rect 18233 22012 18245 22015
rect 18196 21984 18245 22012
rect 18196 21972 18202 21984
rect 18233 21981 18245 21984
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 18524 22021 18552 22052
rect 18616 22021 18644 22120
rect 19518 22108 19524 22160
rect 19576 22148 19582 22160
rect 21910 22148 21916 22160
rect 19576 22120 19747 22148
rect 21871 22120 21916 22148
rect 19576 22108 19582 22120
rect 18874 22040 18880 22092
rect 18932 22080 18938 22092
rect 18932 22052 18977 22080
rect 18932 22040 18938 22052
rect 19242 22040 19248 22092
rect 19300 22080 19306 22092
rect 19613 22083 19671 22089
rect 19613 22080 19625 22083
rect 19300 22052 19625 22080
rect 19300 22040 19306 22052
rect 19613 22049 19625 22052
rect 19659 22049 19671 22083
rect 19719 22080 19747 22120
rect 21910 22108 21916 22120
rect 21968 22108 21974 22160
rect 26418 22108 26424 22160
rect 26476 22148 26482 22160
rect 26602 22148 26608 22160
rect 26476 22120 26608 22148
rect 26476 22108 26482 22120
rect 20990 22080 20996 22092
rect 19719 22052 20996 22080
rect 19613 22043 19671 22049
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 21450 22040 21456 22092
rect 21508 22080 21514 22092
rect 25590 22080 25596 22092
rect 21508 22052 25596 22080
rect 21508 22040 21514 22052
rect 25590 22040 25596 22052
rect 25648 22040 25654 22092
rect 26142 22080 26148 22092
rect 26103 22052 26148 22080
rect 26142 22040 26148 22052
rect 26200 22040 26206 22092
rect 18417 22015 18475 22021
rect 18417 22012 18429 22015
rect 18380 21984 18429 22012
rect 18380 21972 18386 21984
rect 18417 21981 18429 21984
rect 18463 21981 18475 22015
rect 18417 21975 18475 21981
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 21981 18659 22015
rect 19702 22012 19708 22024
rect 18601 21975 18659 21981
rect 18892 21984 19708 22012
rect 18892 21956 18920 21984
rect 19702 21972 19708 21984
rect 19760 21972 19766 22024
rect 21358 21972 21364 22024
rect 21416 22012 21422 22024
rect 23658 22021 23664 22024
rect 21416 21984 21461 22012
rect 21416 21972 21422 21984
rect 23654 21975 23664 22021
rect 23716 22012 23722 22024
rect 26421 22015 26479 22021
rect 23716 21984 23754 22012
rect 23658 21972 23664 21975
rect 23716 21972 23722 21984
rect 26421 21981 26433 22015
rect 26467 22012 26479 22015
rect 26528 22012 26556 22120
rect 26602 22108 26608 22120
rect 26660 22108 26666 22160
rect 28966 22148 28994 22188
rect 29086 22176 29092 22188
rect 29144 22176 29150 22228
rect 29270 22176 29276 22228
rect 29328 22216 29334 22228
rect 29328 22188 31340 22216
rect 29328 22176 29334 22188
rect 30282 22148 30288 22160
rect 26977 22120 28764 22148
rect 28966 22120 30288 22148
rect 26694 22040 26700 22092
rect 26752 22080 26758 22092
rect 26881 22083 26939 22089
rect 26881 22080 26893 22083
rect 26752 22052 26893 22080
rect 26752 22040 26758 22052
rect 26881 22049 26893 22052
rect 26927 22049 26939 22083
rect 26881 22043 26939 22049
rect 26467 21984 26556 22012
rect 26467 21981 26479 21984
rect 26421 21975 26479 21981
rect 17236 21916 17467 21944
rect 17512 21916 17908 21944
rect 17129 21907 17187 21913
rect 9416 21848 11100 21876
rect 11149 21879 11207 21885
rect 11149 21845 11161 21879
rect 11195 21876 11207 21879
rect 12894 21876 12900 21888
rect 11195 21848 12900 21876
rect 11195 21845 11207 21848
rect 11149 21839 11207 21845
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 13262 21876 13268 21888
rect 13223 21848 13268 21876
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 13630 21876 13636 21888
rect 13591 21848 13636 21876
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 14182 21836 14188 21888
rect 14240 21876 14246 21888
rect 17310 21876 17316 21888
rect 14240 21848 17316 21876
rect 14240 21836 14246 21848
rect 17310 21836 17316 21848
rect 17368 21836 17374 21888
rect 17439 21876 17467 21916
rect 17954 21904 17960 21956
rect 18012 21944 18018 21956
rect 18782 21944 18788 21956
rect 18012 21916 18788 21944
rect 18012 21904 18018 21916
rect 18782 21904 18788 21916
rect 18840 21904 18846 21956
rect 18874 21904 18880 21956
rect 18932 21904 18938 21956
rect 19518 21904 19524 21956
rect 19576 21944 19582 21956
rect 21085 21947 21143 21953
rect 19576 21916 19918 21944
rect 19576 21904 19582 21916
rect 21085 21913 21097 21947
rect 21131 21944 21143 21947
rect 21174 21944 21180 21956
rect 21131 21916 21180 21944
rect 21131 21913 21143 21916
rect 21085 21907 21143 21913
rect 21174 21904 21180 21916
rect 21232 21904 21238 21956
rect 22370 21904 22376 21956
rect 22428 21904 22434 21956
rect 23290 21904 23296 21956
rect 23348 21944 23354 21956
rect 24486 21944 24492 21956
rect 23348 21916 24492 21944
rect 23348 21904 23354 21916
rect 24486 21904 24492 21916
rect 24544 21904 24550 21956
rect 24762 21904 24768 21956
rect 24820 21944 24826 21956
rect 24820 21916 24978 21944
rect 24820 21904 24826 21916
rect 25866 21904 25872 21956
rect 25924 21944 25930 21956
rect 26977 21944 27005 22120
rect 27522 22080 27528 22092
rect 25924 21916 27005 21944
rect 27034 22052 27528 22080
rect 25924 21904 25930 21916
rect 22094 21876 22100 21888
rect 17439 21848 22100 21876
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 23014 21836 23020 21888
rect 23072 21876 23078 21888
rect 24578 21876 24584 21888
rect 23072 21848 24584 21876
rect 23072 21836 23078 21848
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 24673 21879 24731 21885
rect 24673 21845 24685 21879
rect 24719 21876 24731 21879
rect 27034 21876 27062 22052
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 28534 22080 28540 22092
rect 28198 22052 28540 22080
rect 28534 22040 28540 22052
rect 28592 22040 28598 22092
rect 28626 22040 28632 22092
rect 28684 22040 28690 22092
rect 27246 22012 27252 22024
rect 27207 21984 27252 22012
rect 27246 21972 27252 21984
rect 27304 21972 27310 22024
rect 27985 22018 28043 22021
rect 27982 21966 27988 22018
rect 28040 22012 28046 22018
rect 28644 22012 28672 22040
rect 28736 22021 28764 22120
rect 30282 22108 30288 22120
rect 30340 22108 30346 22160
rect 29089 22083 29147 22089
rect 29089 22049 29101 22083
rect 29135 22080 29147 22083
rect 30558 22080 30564 22092
rect 29135 22052 29224 22080
rect 29135 22049 29147 22052
rect 29089 22043 29147 22049
rect 28040 21984 28079 22012
rect 28184 21984 28672 22012
rect 28721 22015 28779 22021
rect 28040 21966 28046 21984
rect 28184 21956 28212 21984
rect 28721 21981 28733 22015
rect 28767 21981 28779 22015
rect 28721 21975 28779 21981
rect 28813 22015 28871 22021
rect 28813 21981 28825 22015
rect 28859 21981 28871 22015
rect 28813 21975 28871 21981
rect 27338 21904 27344 21956
rect 27396 21944 27402 21956
rect 27396 21916 27844 21944
rect 27396 21904 27402 21916
rect 24719 21848 27062 21876
rect 24719 21845 24731 21848
rect 24673 21839 24731 21845
rect 27154 21836 27160 21888
rect 27212 21876 27218 21888
rect 27430 21876 27436 21888
rect 27212 21848 27436 21876
rect 27212 21836 27218 21848
rect 27430 21836 27436 21848
rect 27488 21876 27494 21888
rect 27642 21879 27700 21885
rect 27642 21876 27654 21879
rect 27488 21848 27654 21876
rect 27488 21836 27494 21848
rect 27642 21845 27654 21848
rect 27688 21845 27700 21879
rect 27816 21876 27844 21916
rect 28166 21904 28172 21956
rect 28224 21904 28230 21956
rect 28828 21876 28856 21975
rect 28902 21972 28908 22024
rect 28960 21972 28966 22024
rect 28994 21972 29000 22024
rect 29052 22012 29058 22024
rect 29052 21984 29097 22012
rect 29052 21972 29058 21984
rect 28920 21944 28948 21972
rect 28920 21916 29040 21944
rect 27816 21848 28856 21876
rect 27642 21839 27700 21845
rect 28902 21836 28908 21888
rect 28960 21876 28966 21888
rect 29012 21876 29040 21916
rect 29086 21904 29092 21956
rect 29144 21944 29150 21956
rect 29196 21944 29224 22052
rect 30116 22052 30564 22080
rect 30116 22024 30144 22052
rect 30558 22040 30564 22052
rect 30616 22040 30622 22092
rect 29270 21972 29276 22024
rect 29328 22012 29334 22024
rect 29546 22012 29552 22024
rect 29328 21984 29552 22012
rect 29328 21972 29334 21984
rect 29546 21972 29552 21984
rect 29604 21972 29610 22024
rect 29638 21972 29644 22024
rect 29696 22012 29702 22024
rect 29733 22015 29791 22021
rect 29733 22012 29745 22015
rect 29696 21984 29745 22012
rect 29696 21972 29702 21984
rect 29733 21981 29745 21984
rect 29779 21981 29791 22015
rect 30098 22012 30104 22024
rect 30059 21984 30104 22012
rect 29733 21975 29791 21981
rect 30098 21972 30104 21984
rect 30156 21972 30162 22024
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 29822 21944 29828 21956
rect 29144 21916 29224 21944
rect 29783 21916 29828 21944
rect 29144 21904 29150 21916
rect 29822 21904 29828 21916
rect 29880 21904 29886 21956
rect 28960 21848 29040 21876
rect 28960 21836 28966 21848
rect 30098 21836 30104 21888
rect 30156 21876 30162 21888
rect 30208 21876 30236 21975
rect 30374 21972 30380 22024
rect 30432 22012 30438 22024
rect 30837 22015 30895 22021
rect 30837 22012 30849 22015
rect 30432 21984 30849 22012
rect 30432 21972 30438 21984
rect 30837 21981 30849 21984
rect 30883 21981 30895 22015
rect 31018 22012 31024 22024
rect 30979 21984 31024 22012
rect 30837 21975 30895 21981
rect 31018 21972 31024 21984
rect 31076 21972 31082 22024
rect 31312 22021 31340 22188
rect 31297 22015 31355 22021
rect 31297 21981 31309 22015
rect 31343 22012 31355 22015
rect 31478 22012 31484 22024
rect 31343 21984 31484 22012
rect 31343 21981 31355 21984
rect 31297 21975 31355 21981
rect 31478 21972 31484 21984
rect 31536 21972 31542 22024
rect 30156 21848 30236 21876
rect 30156 21836 30162 21848
rect 30282 21836 30288 21888
rect 30340 21876 30346 21888
rect 30377 21879 30435 21885
rect 30377 21876 30389 21879
rect 30340 21848 30389 21876
rect 30340 21836 30346 21848
rect 30377 21845 30389 21848
rect 30423 21845 30435 21879
rect 31110 21876 31116 21888
rect 31071 21848 31116 21876
rect 30377 21839 30435 21845
rect 31110 21836 31116 21848
rect 31168 21836 31174 21888
rect 1104 21786 31992 21808
rect 1104 21734 8632 21786
rect 8684 21734 8696 21786
rect 8748 21734 8760 21786
rect 8812 21734 8824 21786
rect 8876 21734 8888 21786
rect 8940 21734 16314 21786
rect 16366 21734 16378 21786
rect 16430 21734 16442 21786
rect 16494 21734 16506 21786
rect 16558 21734 16570 21786
rect 16622 21734 23996 21786
rect 24048 21734 24060 21786
rect 24112 21734 24124 21786
rect 24176 21734 24188 21786
rect 24240 21734 24252 21786
rect 24304 21734 31678 21786
rect 31730 21734 31742 21786
rect 31794 21734 31806 21786
rect 31858 21734 31870 21786
rect 31922 21734 31934 21786
rect 31986 21734 31992 21786
rect 1104 21712 31992 21734
rect 5442 21672 5448 21684
rect 5403 21644 5448 21672
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 5810 21632 5816 21684
rect 5868 21672 5874 21684
rect 5905 21675 5963 21681
rect 5905 21672 5917 21675
rect 5868 21644 5917 21672
rect 5868 21632 5874 21644
rect 5905 21641 5917 21644
rect 5951 21672 5963 21675
rect 7929 21675 7987 21681
rect 7929 21672 7941 21675
rect 5951 21644 7941 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 7929 21641 7941 21644
rect 7975 21672 7987 21675
rect 8481 21675 8539 21681
rect 8481 21672 8493 21675
rect 7975 21644 8493 21672
rect 7975 21641 7987 21644
rect 7929 21635 7987 21641
rect 8481 21641 8493 21644
rect 8527 21672 8539 21675
rect 9858 21672 9864 21684
rect 8527 21644 9864 21672
rect 8527 21641 8539 21644
rect 8481 21635 8539 21641
rect 9858 21632 9864 21644
rect 9916 21632 9922 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 11238 21672 11244 21684
rect 11195 21644 11244 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 11238 21632 11244 21644
rect 11296 21632 11302 21684
rect 11330 21632 11336 21684
rect 11388 21672 11394 21684
rect 11974 21672 11980 21684
rect 11388 21644 11980 21672
rect 11388 21632 11394 21644
rect 11974 21632 11980 21644
rect 12032 21632 12038 21684
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21672 12311 21675
rect 13262 21672 13268 21684
rect 12299 21644 13268 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 13262 21632 13268 21644
rect 13320 21632 13326 21684
rect 13446 21632 13452 21684
rect 13504 21672 13510 21684
rect 14277 21675 14335 21681
rect 13504 21644 14228 21672
rect 13504 21632 13510 21644
rect 4893 21607 4951 21613
rect 4893 21573 4905 21607
rect 4939 21604 4951 21607
rect 5534 21604 5540 21616
rect 4939 21576 5540 21604
rect 4939 21573 4951 21576
rect 4893 21567 4951 21573
rect 5534 21564 5540 21576
rect 5592 21564 5598 21616
rect 7558 21564 7564 21616
rect 7616 21604 7622 21616
rect 11422 21604 11428 21616
rect 7616 21576 11428 21604
rect 7616 21564 7622 21576
rect 11422 21564 11428 21576
rect 11480 21604 11486 21616
rect 11790 21604 11796 21616
rect 11480 21576 11796 21604
rect 11480 21564 11486 21576
rect 11790 21564 11796 21576
rect 11848 21564 11854 21616
rect 11992 21576 12940 21604
rect 9766 21536 9772 21548
rect 9727 21508 9772 21536
rect 9766 21496 9772 21508
rect 9824 21496 9830 21548
rect 10229 21539 10287 21545
rect 10229 21505 10241 21539
rect 10275 21536 10287 21539
rect 10594 21536 10600 21548
rect 10275 21508 10600 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 10870 21536 10876 21548
rect 10831 21508 10876 21536
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21536 11023 21539
rect 11992 21536 12020 21576
rect 12158 21536 12164 21548
rect 11011 21508 12020 21536
rect 12119 21508 12164 21536
rect 11011 21505 11023 21508
rect 10965 21499 11023 21505
rect 12158 21496 12164 21508
rect 12216 21496 12222 21548
rect 12529 21539 12587 21545
rect 12268 21508 12480 21536
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 9732 21440 9777 21468
rect 9732 21428 9738 21440
rect 9858 21428 9864 21480
rect 9916 21468 9922 21480
rect 11149 21471 11207 21477
rect 11149 21468 11161 21471
rect 9916 21440 11161 21468
rect 9916 21428 9922 21440
rect 11149 21437 11161 21440
rect 11195 21468 11207 21471
rect 12268 21468 12296 21508
rect 11195 21440 12296 21468
rect 12345 21471 12403 21477
rect 11195 21437 11207 21440
rect 11149 21431 11207 21437
rect 12345 21437 12357 21471
rect 12391 21437 12403 21471
rect 12452 21468 12480 21508
rect 12529 21505 12541 21539
rect 12575 21536 12587 21539
rect 12710 21536 12716 21548
rect 12575 21508 12716 21536
rect 12575 21505 12587 21508
rect 12529 21499 12587 21505
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 12912 21536 12940 21576
rect 12986 21564 12992 21616
rect 13044 21604 13050 21616
rect 13998 21604 14004 21616
rect 13044 21576 14004 21604
rect 13044 21564 13050 21576
rect 13998 21564 14004 21576
rect 14056 21564 14062 21616
rect 14200 21604 14228 21644
rect 14277 21641 14289 21675
rect 14323 21672 14335 21675
rect 14918 21672 14924 21684
rect 14323 21644 14924 21672
rect 14323 21641 14335 21644
rect 14277 21635 14335 21641
rect 14918 21632 14924 21644
rect 14976 21632 14982 21684
rect 16022 21672 16028 21684
rect 15580 21644 16028 21672
rect 15580 21604 15608 21644
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 16114 21632 16120 21684
rect 16172 21672 16178 21684
rect 16574 21672 16580 21684
rect 16172 21644 16580 21672
rect 16172 21632 16178 21644
rect 16574 21632 16580 21644
rect 16632 21672 16638 21684
rect 16838 21672 16844 21684
rect 16632 21644 16844 21672
rect 16632 21632 16638 21644
rect 16838 21632 16844 21644
rect 16896 21632 16902 21684
rect 17034 21632 17040 21684
rect 17092 21672 17098 21684
rect 17221 21675 17279 21681
rect 17221 21672 17233 21675
rect 17092 21644 17233 21672
rect 17092 21632 17098 21644
rect 17221 21641 17233 21644
rect 17267 21672 17279 21675
rect 17310 21672 17316 21684
rect 17267 21644 17316 21672
rect 17267 21641 17279 21644
rect 17221 21635 17279 21641
rect 17310 21632 17316 21644
rect 17368 21632 17374 21684
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 18138 21672 18144 21684
rect 17460 21644 18144 21672
rect 17460 21632 17466 21644
rect 18138 21632 18144 21644
rect 18196 21632 18202 21684
rect 18230 21632 18236 21684
rect 18288 21672 18294 21684
rect 18509 21675 18567 21681
rect 18509 21672 18521 21675
rect 18288 21644 18521 21672
rect 18288 21632 18294 21644
rect 18509 21641 18521 21644
rect 18555 21641 18567 21675
rect 18509 21635 18567 21641
rect 18601 21675 18659 21681
rect 18601 21641 18613 21675
rect 18647 21672 18659 21675
rect 19334 21672 19340 21684
rect 18647 21644 19340 21672
rect 18647 21641 18659 21644
rect 18601 21635 18659 21641
rect 16298 21604 16304 21616
rect 14200 21576 15608 21604
rect 15780 21576 16304 21604
rect 13173 21539 13231 21545
rect 13173 21536 13185 21539
rect 12912 21508 13185 21536
rect 13173 21505 13185 21508
rect 13219 21536 13231 21539
rect 14093 21539 14151 21545
rect 14093 21536 14105 21539
rect 13219 21508 14105 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 14093 21505 14105 21508
rect 14139 21505 14151 21539
rect 14093 21499 14151 21505
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21536 15163 21539
rect 15286 21536 15292 21548
rect 15151 21508 15292 21536
rect 15151 21505 15163 21508
rect 15105 21499 15163 21505
rect 13817 21471 13875 21477
rect 13817 21468 13829 21471
rect 12452 21440 13829 21468
rect 12345 21431 12403 21437
rect 13817 21437 13829 21440
rect 13863 21437 13875 21471
rect 13817 21431 13875 21437
rect 6917 21403 6975 21409
rect 6917 21369 6929 21403
rect 6963 21400 6975 21403
rect 9306 21400 9312 21412
rect 6963 21372 9312 21400
rect 6963 21369 6975 21372
rect 6917 21363 6975 21369
rect 9306 21360 9312 21372
rect 9364 21360 9370 21412
rect 10413 21403 10471 21409
rect 10413 21369 10425 21403
rect 10459 21400 10471 21403
rect 10962 21400 10968 21412
rect 10459 21372 10968 21400
rect 10459 21369 10471 21372
rect 10413 21363 10471 21369
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 12250 21360 12256 21412
rect 12308 21400 12314 21412
rect 12360 21400 12388 21431
rect 12526 21400 12532 21412
rect 12308 21372 12388 21400
rect 12487 21372 12532 21400
rect 12308 21360 12314 21372
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 7469 21335 7527 21341
rect 7469 21301 7481 21335
rect 7515 21332 7527 21335
rect 7926 21332 7932 21344
rect 7515 21304 7932 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 7926 21292 7932 21304
rect 7984 21292 7990 21344
rect 8938 21292 8944 21344
rect 8996 21332 9002 21344
rect 9033 21335 9091 21341
rect 9033 21332 9045 21335
rect 8996 21304 9045 21332
rect 8996 21292 9002 21304
rect 9033 21301 9045 21304
rect 9079 21332 9091 21335
rect 9214 21332 9220 21344
rect 9079 21304 9220 21332
rect 9079 21301 9091 21304
rect 9033 21295 9091 21301
rect 9214 21292 9220 21304
rect 9272 21292 9278 21344
rect 10502 21292 10508 21344
rect 10560 21332 10566 21344
rect 12986 21332 12992 21344
rect 10560 21304 12992 21332
rect 10560 21292 10566 21304
rect 12986 21292 12992 21304
rect 13044 21292 13050 21344
rect 13354 21332 13360 21344
rect 13315 21304 13360 21332
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 13832 21332 13860 21431
rect 13906 21428 13912 21480
rect 13964 21468 13970 21480
rect 13964 21440 14009 21468
rect 13964 21428 13970 21440
rect 14108 21400 14136 21499
rect 15286 21496 15292 21508
rect 15344 21496 15350 21548
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 14700 21440 14749 21468
rect 14700 21428 14706 21440
rect 14737 21437 14749 21440
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 15197 21471 15255 21477
rect 15197 21437 15209 21471
rect 15243 21468 15255 21471
rect 15780 21468 15808 21576
rect 16298 21564 16304 21576
rect 16356 21564 16362 21616
rect 16666 21564 16672 21616
rect 16724 21604 16730 21616
rect 17589 21607 17647 21613
rect 17589 21604 17601 21607
rect 16724 21576 17601 21604
rect 16724 21564 16730 21576
rect 17589 21573 17601 21576
rect 17635 21604 17647 21607
rect 18616 21604 18644 21635
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 19886 21632 19892 21684
rect 19944 21672 19950 21684
rect 21358 21672 21364 21684
rect 19944 21644 21364 21672
rect 19944 21632 19950 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 22554 21672 22560 21684
rect 22336 21644 22560 21672
rect 22336 21632 22342 21644
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 23382 21672 23388 21684
rect 22796 21644 23388 21672
rect 22796 21632 22802 21644
rect 23382 21632 23388 21644
rect 23440 21672 23446 21684
rect 23658 21672 23664 21684
rect 23440 21644 23664 21672
rect 23440 21632 23446 21644
rect 23658 21632 23664 21644
rect 23716 21672 23722 21684
rect 23716 21644 23796 21672
rect 23716 21632 23722 21644
rect 17635 21576 18644 21604
rect 17635 21573 17647 21576
rect 17589 21567 17647 21573
rect 18690 21564 18696 21616
rect 18748 21604 18754 21616
rect 19150 21604 19156 21616
rect 18748 21576 19156 21604
rect 18748 21564 18754 21576
rect 19150 21564 19156 21576
rect 19208 21564 19214 21616
rect 19904 21604 19932 21632
rect 19444 21576 19932 21604
rect 15930 21536 15936 21548
rect 15891 21508 15936 21536
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 16022 21496 16028 21548
rect 16080 21536 16086 21548
rect 17405 21539 17463 21545
rect 17405 21536 17417 21539
rect 16080 21508 17417 21536
rect 16080 21496 16086 21508
rect 17405 21505 17417 21508
rect 17451 21505 17463 21539
rect 17405 21499 17463 21505
rect 17497 21539 17555 21545
rect 17497 21505 17509 21539
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 15243 21440 15808 21468
rect 15841 21471 15899 21477
rect 15243 21437 15255 21440
rect 15197 21431 15255 21437
rect 15841 21437 15853 21471
rect 15887 21468 15899 21471
rect 17512 21468 17540 21499
rect 17678 21496 17684 21548
rect 17736 21536 17742 21548
rect 17773 21539 17831 21545
rect 17773 21536 17785 21539
rect 17736 21508 17785 21536
rect 17736 21496 17742 21508
rect 17773 21505 17785 21508
rect 17819 21536 17831 21539
rect 18966 21536 18972 21548
rect 17819 21508 18972 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18966 21496 18972 21508
rect 19024 21496 19030 21548
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 19444 21545 19472 21576
rect 19978 21564 19984 21616
rect 20036 21604 20042 21616
rect 20036 21576 20194 21604
rect 20036 21564 20042 21576
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 21453 21607 21511 21613
rect 21453 21604 21465 21607
rect 21048 21576 21465 21604
rect 21048 21564 21054 21576
rect 21453 21573 21465 21576
rect 21499 21573 21511 21607
rect 23768 21604 23796 21644
rect 23842 21632 23848 21684
rect 23900 21672 23906 21684
rect 29822 21672 29828 21684
rect 23900 21644 29828 21672
rect 23900 21632 23906 21644
rect 29822 21632 29828 21644
rect 29880 21632 29886 21684
rect 30742 21632 30748 21684
rect 30800 21632 30806 21684
rect 23768 21576 23888 21604
rect 21453 21567 21511 21573
rect 19429 21539 19487 21545
rect 19429 21536 19441 21539
rect 19392 21508 19441 21536
rect 19392 21496 19398 21508
rect 19429 21505 19441 21508
rect 19475 21505 19487 21539
rect 19429 21499 19487 21505
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 23860 21545 23888 21576
rect 26326 21564 26332 21616
rect 26384 21604 26390 21616
rect 26694 21604 26700 21616
rect 26384 21576 26700 21604
rect 26384 21564 26390 21576
rect 26694 21564 26700 21576
rect 26752 21564 26758 21616
rect 26786 21564 26792 21616
rect 26844 21604 26850 21616
rect 26970 21604 26976 21616
rect 26844 21576 26976 21604
rect 26844 21564 26850 21576
rect 26970 21564 26976 21576
rect 27028 21564 27034 21616
rect 27154 21564 27160 21616
rect 27212 21604 27218 21616
rect 27433 21607 27491 21613
rect 27433 21604 27445 21607
rect 27212 21576 27445 21604
rect 27212 21564 27218 21576
rect 27433 21573 27445 21576
rect 27479 21573 27491 21607
rect 27433 21567 27491 21573
rect 28166 21564 28172 21616
rect 28224 21564 28230 21616
rect 28810 21564 28816 21616
rect 28868 21604 28874 21616
rect 28868 21576 29500 21604
rect 28868 21564 28874 21576
rect 23845 21539 23903 21545
rect 22152 21508 22494 21536
rect 22152 21496 22158 21508
rect 23845 21505 23857 21539
rect 23891 21505 23903 21539
rect 23845 21499 23903 21505
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 24728 21508 25254 21536
rect 24728 21496 24734 21508
rect 26602 21496 26608 21548
rect 26660 21536 26666 21548
rect 26660 21508 27200 21536
rect 26660 21496 26666 21508
rect 17586 21468 17592 21480
rect 15887 21440 17592 21468
rect 15887 21437 15899 21440
rect 15841 21431 15899 21437
rect 15856 21400 15884 21431
rect 17586 21428 17592 21440
rect 17644 21468 17650 21480
rect 18230 21468 18236 21480
rect 17644 21440 18236 21468
rect 17644 21428 17650 21440
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 18414 21468 18420 21480
rect 18375 21440 18420 21468
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 18506 21428 18512 21480
rect 18564 21468 18570 21480
rect 18690 21468 18696 21480
rect 18564 21440 18696 21468
rect 18564 21428 18570 21440
rect 18690 21428 18696 21440
rect 18748 21428 18754 21480
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 19705 21471 19763 21477
rect 19705 21468 19717 21471
rect 18840 21440 19717 21468
rect 18840 21428 18846 21440
rect 19705 21437 19717 21440
rect 19751 21437 19763 21471
rect 19705 21431 19763 21437
rect 19794 21428 19800 21480
rect 19852 21468 19858 21480
rect 23569 21471 23627 21477
rect 23569 21468 23581 21471
rect 19852 21440 23581 21468
rect 19852 21428 19858 21440
rect 23569 21437 23581 21440
rect 23615 21437 23627 21471
rect 23569 21431 23627 21437
rect 26329 21471 26387 21477
rect 26329 21437 26341 21471
rect 26375 21468 26387 21471
rect 26970 21468 26976 21480
rect 26375 21440 26976 21468
rect 26375 21437 26387 21440
rect 26329 21431 26387 21437
rect 26970 21428 26976 21440
rect 27028 21428 27034 21480
rect 27172 21477 27200 21508
rect 28902 21496 28908 21548
rect 28960 21536 28966 21548
rect 29472 21545 29500 21576
rect 29546 21564 29552 21616
rect 29604 21604 29610 21616
rect 29641 21607 29699 21613
rect 29641 21604 29653 21607
rect 29604 21576 29653 21604
rect 29604 21564 29610 21576
rect 29641 21573 29653 21576
rect 29687 21573 29699 21607
rect 29641 21567 29699 21573
rect 29733 21607 29791 21613
rect 29733 21573 29745 21607
rect 29779 21604 29791 21607
rect 29914 21604 29920 21616
rect 29779 21576 29920 21604
rect 29779 21573 29791 21576
rect 29733 21567 29791 21573
rect 29914 21564 29920 21576
rect 29972 21564 29978 21616
rect 29365 21539 29423 21545
rect 29365 21536 29377 21539
rect 28960 21508 29377 21536
rect 28960 21496 28966 21508
rect 29365 21505 29377 21508
rect 29411 21505 29423 21539
rect 29365 21499 29423 21505
rect 29457 21539 29515 21545
rect 29457 21505 29469 21539
rect 29503 21505 29515 21539
rect 29457 21499 29515 21505
rect 29825 21539 29883 21545
rect 29825 21505 29837 21539
rect 29871 21536 29883 21539
rect 30282 21536 30288 21548
rect 29871 21508 30288 21536
rect 29871 21505 29883 21508
rect 29825 21499 29883 21505
rect 30282 21496 30288 21508
rect 30340 21496 30346 21548
rect 30469 21539 30527 21545
rect 30469 21505 30481 21539
rect 30515 21505 30527 21539
rect 30650 21536 30656 21548
rect 30611 21508 30656 21536
rect 30469 21499 30527 21505
rect 27157 21471 27215 21477
rect 27157 21437 27169 21471
rect 27203 21437 27215 21471
rect 30374 21468 30380 21480
rect 27157 21431 27215 21437
rect 27264 21440 30380 21468
rect 14108 21372 15884 21400
rect 15930 21360 15936 21412
rect 15988 21400 15994 21412
rect 17678 21400 17684 21412
rect 15988 21372 17684 21400
rect 15988 21360 15994 21372
rect 17678 21360 17684 21372
rect 17736 21360 17742 21412
rect 17770 21360 17776 21412
rect 17828 21400 17834 21412
rect 17828 21372 19012 21400
rect 17828 21360 17834 21372
rect 15948 21332 15976 21360
rect 13832 21304 15976 21332
rect 16301 21335 16359 21341
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 18414 21332 18420 21344
rect 16347 21304 18420 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 18984 21341 19012 21372
rect 19242 21360 19248 21412
rect 19300 21400 19306 21412
rect 19426 21400 19432 21412
rect 19300 21372 19432 21400
rect 19300 21360 19306 21372
rect 19426 21360 19432 21372
rect 19484 21360 19490 21412
rect 20714 21360 20720 21412
rect 20772 21400 20778 21412
rect 20772 21372 20944 21400
rect 20772 21360 20778 21372
rect 18969 21335 19027 21341
rect 18969 21301 18981 21335
rect 19015 21332 19027 21335
rect 20806 21332 20812 21344
rect 19015 21304 20812 21332
rect 19015 21301 19027 21304
rect 18969 21295 19027 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 20916 21332 20944 21372
rect 20990 21360 20996 21412
rect 21048 21400 21054 21412
rect 21818 21400 21824 21412
rect 21048 21372 21824 21400
rect 21048 21360 21054 21372
rect 21818 21360 21824 21372
rect 21876 21360 21882 21412
rect 22097 21403 22155 21409
rect 22097 21369 22109 21403
rect 22143 21400 22155 21403
rect 22462 21400 22468 21412
rect 22143 21372 22468 21400
rect 22143 21369 22155 21372
rect 22097 21363 22155 21369
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 24857 21403 24915 21409
rect 24857 21369 24869 21403
rect 24903 21400 24915 21403
rect 24946 21400 24952 21412
rect 24903 21372 24952 21400
rect 24903 21369 24915 21372
rect 24857 21363 24915 21369
rect 24946 21360 24952 21372
rect 25004 21360 25010 21412
rect 27264 21400 27292 21440
rect 30374 21428 30380 21440
rect 30432 21428 30438 21480
rect 26528 21372 27292 21400
rect 23014 21332 23020 21344
rect 20916 21304 23020 21332
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 23198 21292 23204 21344
rect 23256 21332 23262 21344
rect 26528 21332 26556 21372
rect 28442 21360 28448 21412
rect 28500 21400 28506 21412
rect 29362 21400 29368 21412
rect 28500 21372 29368 21400
rect 28500 21360 28506 21372
rect 29362 21360 29368 21372
rect 29420 21360 29426 21412
rect 30484 21400 30512 21499
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 30760 21545 30788 21632
rect 30745 21539 30803 21545
rect 30745 21505 30757 21539
rect 30791 21505 30803 21539
rect 30745 21499 30803 21505
rect 30834 21496 30840 21548
rect 30892 21536 30898 21548
rect 30892 21508 30937 21536
rect 30892 21496 30898 21508
rect 30650 21400 30656 21412
rect 30484 21372 30656 21400
rect 30650 21360 30656 21372
rect 30708 21360 30714 21412
rect 23256 21304 26556 21332
rect 23256 21292 23262 21304
rect 26970 21292 26976 21344
rect 27028 21332 27034 21344
rect 28810 21332 28816 21344
rect 27028 21304 28816 21332
rect 27028 21292 27034 21304
rect 28810 21292 28816 21304
rect 28868 21292 28874 21344
rect 28902 21292 28908 21344
rect 28960 21332 28966 21344
rect 28960 21304 29005 21332
rect 28960 21292 28966 21304
rect 29454 21292 29460 21344
rect 29512 21332 29518 21344
rect 30009 21335 30067 21341
rect 30009 21332 30021 21335
rect 29512 21304 30021 21332
rect 29512 21292 29518 21304
rect 30009 21301 30021 21304
rect 30055 21301 30067 21335
rect 31110 21332 31116 21344
rect 31071 21304 31116 21332
rect 30009 21295 30067 21301
rect 31110 21292 31116 21304
rect 31168 21292 31174 21344
rect 1104 21242 31832 21264
rect 1104 21190 4791 21242
rect 4843 21190 4855 21242
rect 4907 21190 4919 21242
rect 4971 21190 4983 21242
rect 5035 21190 5047 21242
rect 5099 21190 12473 21242
rect 12525 21190 12537 21242
rect 12589 21190 12601 21242
rect 12653 21190 12665 21242
rect 12717 21190 12729 21242
rect 12781 21190 20155 21242
rect 20207 21190 20219 21242
rect 20271 21190 20283 21242
rect 20335 21190 20347 21242
rect 20399 21190 20411 21242
rect 20463 21190 27837 21242
rect 27889 21190 27901 21242
rect 27953 21190 27965 21242
rect 28017 21190 28029 21242
rect 28081 21190 28093 21242
rect 28145 21190 31832 21242
rect 1104 21168 31832 21190
rect 5261 21131 5319 21137
rect 5261 21097 5273 21131
rect 5307 21128 5319 21131
rect 7466 21128 7472 21140
rect 5307 21100 7472 21128
rect 5307 21097 5319 21100
rect 5261 21091 5319 21097
rect 7466 21088 7472 21100
rect 7524 21088 7530 21140
rect 7650 21088 7656 21140
rect 7708 21128 7714 21140
rect 8294 21128 8300 21140
rect 7708 21100 8300 21128
rect 7708 21088 7714 21100
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 9122 21088 9128 21140
rect 9180 21128 9186 21140
rect 11790 21128 11796 21140
rect 9180 21100 11796 21128
rect 9180 21088 9186 21100
rect 11790 21088 11796 21100
rect 11848 21088 11854 21140
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 12529 21131 12587 21137
rect 12529 21128 12541 21131
rect 12492 21100 12541 21128
rect 12492 21088 12498 21100
rect 12529 21097 12541 21100
rect 12575 21097 12587 21131
rect 12529 21091 12587 21097
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 14461 21131 14519 21137
rect 14461 21128 14473 21131
rect 13412 21100 14473 21128
rect 13412 21088 13418 21100
rect 14461 21097 14473 21100
rect 14507 21097 14519 21131
rect 14461 21091 14519 21097
rect 15378 21088 15384 21140
rect 15436 21128 15442 21140
rect 16482 21128 16488 21140
rect 15436 21100 16488 21128
rect 15436 21088 15442 21100
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 16577 21131 16635 21137
rect 16577 21097 16589 21131
rect 16623 21128 16635 21131
rect 17862 21128 17868 21140
rect 16623 21100 17868 21128
rect 16623 21097 16635 21100
rect 16577 21091 16635 21097
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 18046 21088 18052 21140
rect 18104 21128 18110 21140
rect 18104 21100 18644 21128
rect 18104 21088 18110 21100
rect 10594 21020 10600 21072
rect 10652 21060 10658 21072
rect 14277 21063 14335 21069
rect 14277 21060 14289 21063
rect 10652 21032 14289 21060
rect 10652 21020 10658 21032
rect 14277 21029 14289 21032
rect 14323 21029 14335 21063
rect 15010 21060 15016 21072
rect 14277 21023 14335 21029
rect 14400 21032 15016 21060
rect 6917 20995 6975 21001
rect 6917 20961 6929 20995
rect 6963 20992 6975 20995
rect 8294 20992 8300 21004
rect 6963 20964 8300 20992
rect 6963 20961 6975 20964
rect 6917 20955 6975 20961
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 9306 20952 9312 21004
rect 9364 20992 9370 21004
rect 11241 21000 11299 21001
rect 11422 21000 11428 21004
rect 11241 20995 11428 21000
rect 9364 20964 11192 20992
rect 9364 20952 9370 20964
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20924 9735 20927
rect 9950 20924 9956 20936
rect 9723 20896 9956 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 9950 20884 9956 20896
rect 10008 20924 10014 20936
rect 10226 20924 10232 20936
rect 10008 20896 10232 20924
rect 10008 20884 10014 20896
rect 10226 20884 10232 20896
rect 10284 20884 10290 20936
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20893 10379 20927
rect 10502 20924 10508 20936
rect 10463 20896 10508 20924
rect 10321 20887 10379 20893
rect 8294 20816 8300 20868
rect 8352 20856 8358 20868
rect 8938 20856 8944 20868
rect 8352 20828 8944 20856
rect 8352 20816 8358 20828
rect 8938 20816 8944 20828
rect 8996 20856 9002 20868
rect 9125 20859 9183 20865
rect 9125 20856 9137 20859
rect 8996 20828 9137 20856
rect 8996 20816 9002 20828
rect 9125 20825 9137 20828
rect 9171 20825 9183 20859
rect 9125 20819 9183 20825
rect 5813 20791 5871 20797
rect 5813 20757 5825 20791
rect 5859 20788 5871 20791
rect 5994 20788 6000 20800
rect 5859 20760 6000 20788
rect 5859 20757 5871 20760
rect 5813 20751 5871 20757
rect 5994 20748 6000 20760
rect 6052 20748 6058 20800
rect 6365 20791 6423 20797
rect 6365 20757 6377 20791
rect 6411 20788 6423 20791
rect 7374 20788 7380 20800
rect 6411 20760 7380 20788
rect 6411 20757 6423 20760
rect 6365 20751 6423 20757
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 8018 20788 8024 20800
rect 7979 20760 8024 20788
rect 8018 20748 8024 20760
rect 8076 20748 8082 20800
rect 8110 20748 8116 20800
rect 8168 20788 8174 20800
rect 8386 20788 8392 20800
rect 8168 20760 8392 20788
rect 8168 20748 8174 20760
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 8573 20791 8631 20797
rect 8573 20757 8585 20791
rect 8619 20788 8631 20791
rect 9030 20788 9036 20800
rect 8619 20760 9036 20788
rect 8619 20757 8631 20760
rect 8573 20751 8631 20757
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 9140 20788 9168 20819
rect 9490 20816 9496 20868
rect 9548 20856 9554 20868
rect 10336 20856 10364 20887
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 10870 20884 10876 20936
rect 10928 20924 10934 20936
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 10928 20896 10977 20924
rect 10928 20884 10934 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11057 20927 11115 20933
rect 11057 20893 11069 20927
rect 11103 20893 11115 20927
rect 11164 20924 11192 20964
rect 11241 20961 11253 20995
rect 11287 20972 11428 20995
rect 11287 20961 11299 20972
rect 11241 20955 11299 20961
rect 11422 20952 11428 20972
rect 11480 20952 11486 21004
rect 11974 20952 11980 21004
rect 12032 20992 12038 21004
rect 12713 20995 12771 21001
rect 12032 20964 12664 20992
rect 12032 20952 12038 20964
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 11164 20896 11713 20924
rect 11057 20887 11115 20893
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 9548 20828 10364 20856
rect 9548 20816 9554 20828
rect 11072 20800 11100 20887
rect 11146 20816 11152 20868
rect 11204 20856 11210 20868
rect 11716 20856 11744 20887
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 11885 20927 11943 20933
rect 11885 20924 11897 20927
rect 11848 20896 11897 20924
rect 11848 20884 11854 20896
rect 11885 20893 11897 20896
rect 11931 20893 11943 20927
rect 12066 20924 12072 20936
rect 12027 20896 12072 20924
rect 11885 20887 11943 20893
rect 12066 20884 12072 20896
rect 12124 20884 12130 20936
rect 12526 20924 12532 20936
rect 12487 20896 12532 20924
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 12636 20924 12664 20964
rect 12713 20961 12725 20995
rect 12759 20992 12771 20995
rect 13170 20992 13176 21004
rect 12759 20964 13176 20992
rect 12759 20961 12771 20964
rect 12713 20955 12771 20961
rect 12897 20927 12955 20933
rect 12897 20924 12909 20927
rect 12636 20896 12909 20924
rect 12897 20893 12909 20896
rect 12943 20893 12955 20927
rect 12897 20887 12955 20893
rect 13004 20856 13032 20964
rect 13170 20952 13176 20964
rect 13228 20952 13234 21004
rect 13446 20952 13452 21004
rect 13504 20952 13510 21004
rect 13725 20995 13783 21001
rect 13725 20961 13737 20995
rect 13771 20992 13783 20995
rect 14400 20992 14428 21032
rect 15010 21020 15016 21032
rect 15068 21060 15074 21072
rect 15105 21063 15163 21069
rect 15105 21060 15117 21063
rect 15068 21032 15117 21060
rect 15068 21020 15074 21032
rect 15105 21029 15117 21032
rect 15151 21029 15163 21063
rect 16114 21060 16120 21072
rect 15105 21023 15163 21029
rect 15196 21032 16120 21060
rect 13771 20964 14428 20992
rect 13771 20961 13783 20964
rect 13725 20955 13783 20961
rect 14458 20952 14464 21004
rect 14516 20992 14522 21004
rect 15196 20992 15224 21032
rect 16114 21020 16120 21032
rect 16172 21020 16178 21072
rect 16298 21020 16304 21072
rect 16356 21060 16362 21072
rect 16850 21060 16856 21072
rect 16356 21032 16856 21060
rect 16356 21020 16362 21032
rect 16850 21020 16856 21032
rect 16908 21020 16914 21072
rect 17770 21060 17776 21072
rect 17052 21032 17776 21060
rect 16390 20992 16396 21004
rect 14516 20964 15224 20992
rect 15488 20964 16396 20992
rect 14516 20952 14522 20964
rect 13350 20927 13408 20933
rect 13350 20893 13362 20927
rect 13396 20924 13408 20927
rect 13464 20924 13492 20952
rect 15488 20933 15516 20964
rect 16390 20952 16396 20964
rect 16448 20952 16454 21004
rect 16482 20952 16488 21004
rect 16540 20992 16546 21004
rect 17052 20992 17080 21032
rect 17770 21020 17776 21032
rect 17828 21020 17834 21072
rect 18616 21060 18644 21100
rect 18690 21088 18696 21140
rect 18748 21128 18754 21140
rect 19978 21128 19984 21140
rect 18748 21100 19984 21128
rect 18748 21088 18754 21100
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 21450 21128 21456 21140
rect 20088 21100 21456 21128
rect 18782 21060 18788 21072
rect 18616 21032 18788 21060
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 18877 21063 18935 21069
rect 18877 21029 18889 21063
rect 18923 21060 18935 21063
rect 20088 21060 20116 21100
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 24765 21131 24823 21137
rect 24765 21097 24777 21131
rect 24811 21128 24823 21131
rect 25498 21128 25504 21140
rect 24811 21100 25504 21128
rect 24811 21097 24823 21100
rect 24765 21091 24823 21097
rect 25498 21088 25504 21100
rect 25556 21088 25562 21140
rect 25590 21088 25596 21140
rect 25648 21128 25654 21140
rect 28994 21128 29000 21140
rect 25648 21100 29000 21128
rect 25648 21088 25654 21100
rect 28994 21088 29000 21100
rect 29052 21088 29058 21140
rect 29362 21088 29368 21140
rect 29420 21128 29426 21140
rect 30837 21131 30895 21137
rect 30837 21128 30849 21131
rect 29420 21100 30849 21128
rect 29420 21088 29426 21100
rect 30837 21097 30849 21100
rect 30883 21097 30895 21131
rect 31294 21128 31300 21140
rect 31255 21100 31300 21128
rect 30837 21091 30895 21097
rect 31294 21088 31300 21100
rect 31352 21088 31358 21140
rect 29730 21060 29736 21072
rect 18923 21032 20116 21060
rect 21252 21032 23612 21060
rect 29691 21032 29736 21060
rect 18923 21029 18935 21032
rect 18877 21023 18935 21029
rect 17586 20992 17592 21004
rect 16540 20964 17080 20992
rect 17328 20964 17592 20992
rect 16540 20952 16546 20964
rect 15381 20927 15439 20933
rect 15381 20924 15393 20927
rect 13396 20896 13492 20924
rect 13648 20896 15393 20924
rect 13396 20893 13408 20896
rect 13350 20887 13408 20893
rect 11204 20828 11652 20856
rect 11716 20828 11928 20856
rect 11204 20816 11210 20828
rect 9582 20788 9588 20800
rect 9140 20760 9588 20788
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 9766 20788 9772 20800
rect 9727 20760 9772 20788
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 10410 20788 10416 20800
rect 10371 20760 10416 20788
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 11054 20748 11060 20800
rect 11112 20748 11118 20800
rect 11238 20788 11244 20800
rect 11199 20760 11244 20788
rect 11238 20748 11244 20760
rect 11296 20748 11302 20800
rect 11624 20788 11652 20828
rect 11790 20788 11796 20800
rect 11624 20760 11796 20788
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 11900 20788 11928 20828
rect 12544 20828 13032 20856
rect 13449 20859 13507 20865
rect 12544 20788 12572 20828
rect 13449 20825 13461 20859
rect 13495 20856 13507 20859
rect 13648 20856 13676 20896
rect 15381 20893 15393 20896
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20893 15531 20927
rect 15473 20887 15531 20893
rect 14645 20859 14703 20865
rect 14645 20856 14657 20859
rect 13495 20828 13676 20856
rect 13740 20828 14657 20856
rect 13495 20825 13507 20828
rect 13449 20819 13507 20825
rect 11900 20760 12572 20788
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 12805 20791 12863 20797
rect 12805 20788 12817 20791
rect 12676 20760 12817 20788
rect 12676 20748 12682 20760
rect 12805 20757 12817 20760
rect 12851 20757 12863 20791
rect 12805 20751 12863 20757
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 13541 20791 13599 20797
rect 13541 20788 13553 20791
rect 13136 20760 13553 20788
rect 13136 20748 13142 20760
rect 13541 20757 13553 20760
rect 13587 20788 13599 20791
rect 13630 20788 13636 20800
rect 13587 20760 13636 20788
rect 13587 20757 13599 20760
rect 13541 20751 13599 20757
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 13740 20797 13768 20828
rect 14645 20825 14657 20828
rect 14691 20856 14703 20859
rect 15194 20856 15200 20868
rect 14691 20828 15200 20856
rect 14691 20825 14703 20828
rect 14645 20819 14703 20825
rect 15194 20816 15200 20828
rect 15252 20816 15258 20868
rect 15396 20856 15424 20887
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 15804 20896 16313 20924
rect 15804 20884 15810 20896
rect 16301 20893 16313 20896
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 17328 20933 17356 20964
rect 17586 20952 17592 20964
rect 17644 20992 17650 21004
rect 20714 20992 20720 21004
rect 17644 20964 20720 20992
rect 17644 20952 17650 20964
rect 17117 20927 17175 20933
rect 17117 20924 17129 20927
rect 16632 20896 17129 20924
rect 16632 20884 16638 20896
rect 17117 20893 17129 20896
rect 17163 20893 17175 20927
rect 17117 20887 17175 20893
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 18230 20924 18236 20936
rect 17543 20921 17954 20924
rect 17543 20896 18092 20921
rect 18191 20896 18236 20924
rect 17543 20893 17555 20896
rect 17926 20893 18092 20896
rect 17497 20887 17555 20893
rect 15838 20856 15844 20868
rect 15396 20828 15844 20856
rect 15838 20816 15844 20828
rect 15896 20816 15902 20868
rect 16022 20816 16028 20868
rect 16080 20856 16086 20868
rect 16758 20856 16764 20868
rect 16080 20828 16764 20856
rect 16080 20816 16086 20828
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 17328 20856 17356 20887
rect 17144 20828 17356 20856
rect 14458 20797 14464 20800
rect 13725 20791 13783 20797
rect 13725 20757 13737 20791
rect 13771 20757 13783 20791
rect 13725 20751 13783 20757
rect 14445 20791 14464 20797
rect 14445 20757 14457 20791
rect 14445 20751 14464 20757
rect 14458 20748 14464 20751
rect 14516 20748 14522 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 15289 20791 15347 20797
rect 15289 20788 15301 20791
rect 14792 20760 15301 20788
rect 14792 20748 14798 20760
rect 15289 20757 15301 20760
rect 15335 20788 15347 20791
rect 15470 20788 15476 20800
rect 15335 20760 15476 20788
rect 15335 20757 15347 20760
rect 15289 20751 15347 20757
rect 15470 20748 15476 20760
rect 15528 20748 15534 20800
rect 15654 20788 15660 20800
rect 15615 20760 15660 20788
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 17144 20788 17172 20828
rect 15988 20760 17172 20788
rect 15988 20748 15994 20760
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 17420 20788 17448 20887
rect 17678 20816 17684 20868
rect 17736 20856 17742 20868
rect 17773 20859 17831 20865
rect 17773 20856 17785 20859
rect 17736 20828 17785 20856
rect 17736 20816 17742 20828
rect 17773 20825 17785 20828
rect 17819 20825 17831 20859
rect 18064 20856 18092 20893
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 18322 20884 18328 20936
rect 18380 20924 18386 20936
rect 18524 20933 18552 20964
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 21252 20992 21280 21032
rect 20864 20964 21280 20992
rect 20864 20952 20870 20964
rect 21542 20952 21548 21004
rect 21600 20992 21606 21004
rect 23584 21001 23612 21032
rect 29730 21020 29736 21032
rect 29788 21020 29794 21072
rect 30006 21020 30012 21072
rect 30064 21060 30070 21072
rect 30064 21032 30972 21060
rect 30064 21020 30070 21032
rect 22005 20995 22063 21001
rect 22005 20992 22017 20995
rect 21600 20964 22017 20992
rect 21600 20952 21606 20964
rect 22005 20961 22017 20964
rect 22051 20961 22063 20995
rect 22005 20955 22063 20961
rect 23569 20995 23627 21001
rect 23569 20961 23581 20995
rect 23615 20992 23627 20995
rect 27338 20992 27344 21004
rect 23615 20964 27344 20992
rect 23615 20961 23627 20964
rect 23569 20955 23627 20961
rect 27338 20952 27344 20964
rect 27396 20952 27402 21004
rect 27614 20952 27620 21004
rect 27672 20992 27678 21004
rect 27672 20964 28488 20992
rect 27672 20952 27678 20964
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18380 20896 18429 20924
rect 18380 20884 18386 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20893 18567 20927
rect 18509 20887 18567 20893
rect 18598 20884 18604 20936
rect 18656 20924 18662 20936
rect 18656 20896 18701 20924
rect 18656 20884 18662 20896
rect 18782 20884 18788 20936
rect 18840 20924 18846 20936
rect 19794 20924 19800 20936
rect 18840 20896 19800 20924
rect 18840 20884 18846 20896
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 19886 20884 19892 20936
rect 19944 20924 19950 20936
rect 19981 20927 20039 20933
rect 19981 20924 19993 20927
rect 19944 20896 19993 20924
rect 19944 20884 19950 20896
rect 19981 20893 19993 20896
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 22741 20927 22799 20933
rect 22741 20893 22753 20927
rect 22787 20893 22799 20927
rect 22741 20887 22799 20893
rect 23201 20927 23259 20933
rect 23201 20893 23213 20927
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 26513 20927 26571 20933
rect 26513 20893 26525 20927
rect 26559 20924 26571 20927
rect 26694 20924 26700 20936
rect 26559 20896 26700 20924
rect 26559 20893 26571 20896
rect 26513 20887 26571 20893
rect 18138 20856 18144 20868
rect 18064 20828 18144 20856
rect 17773 20819 17831 20825
rect 18138 20816 18144 20828
rect 18196 20816 18202 20868
rect 20264 20859 20322 20865
rect 18248 20828 20195 20856
rect 18248 20788 18276 20828
rect 17276 20760 18276 20788
rect 17276 20748 17282 20760
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 19521 20791 19579 20797
rect 19521 20788 19533 20791
rect 18380 20760 19533 20788
rect 18380 20748 18386 20760
rect 19521 20757 19533 20760
rect 19567 20788 19579 20791
rect 20070 20788 20076 20800
rect 19567 20760 20076 20788
rect 19567 20757 19579 20760
rect 19521 20751 19579 20757
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 20167 20788 20195 20828
rect 20264 20825 20276 20859
rect 20310 20856 20322 20859
rect 20530 20856 20536 20868
rect 20310 20828 20536 20856
rect 20310 20825 20322 20828
rect 20264 20819 20322 20825
rect 20530 20816 20536 20828
rect 20588 20816 20594 20868
rect 20990 20816 20996 20868
rect 21048 20816 21054 20868
rect 20622 20788 20628 20800
rect 20167 20760 20628 20788
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 20898 20748 20904 20800
rect 20956 20788 20962 20800
rect 22756 20788 22784 20887
rect 23216 20856 23244 20887
rect 26694 20884 26700 20896
rect 26752 20884 26758 20936
rect 26962 20927 27020 20933
rect 26962 20924 26974 20927
rect 26896 20896 26974 20924
rect 23216 20828 24992 20856
rect 20956 20760 22784 20788
rect 24964 20788 24992 20828
rect 25222 20816 25228 20868
rect 25280 20816 25286 20868
rect 26234 20856 26240 20868
rect 26195 20828 26240 20856
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 26602 20816 26608 20868
rect 26660 20856 26666 20868
rect 26896 20856 26924 20896
rect 26962 20893 26974 20896
rect 27008 20893 27020 20927
rect 28460 20924 28488 20964
rect 28534 20952 28540 21004
rect 28592 20992 28598 21004
rect 29822 20992 29828 21004
rect 28592 20964 29828 20992
rect 28592 20952 28598 20964
rect 29822 20952 29828 20964
rect 29880 20952 29886 21004
rect 30101 20995 30159 21001
rect 30101 20961 30113 20995
rect 30147 20992 30159 20995
rect 30190 20992 30196 21004
rect 30147 20964 30196 20992
rect 30147 20961 30159 20964
rect 30101 20955 30159 20961
rect 30190 20952 30196 20964
rect 30248 20952 30254 21004
rect 30944 21001 30972 21032
rect 30929 20995 30987 21001
rect 30929 20961 30941 20995
rect 30975 20961 30987 20995
rect 30929 20955 30987 20961
rect 28460 20896 30141 20924
rect 26962 20887 27020 20893
rect 27246 20856 27252 20868
rect 26660 20828 26924 20856
rect 27207 20828 27252 20856
rect 26660 20816 26666 20828
rect 27246 20816 27252 20828
rect 27304 20816 27310 20868
rect 28534 20856 28540 20868
rect 28474 20828 28540 20856
rect 28534 20816 28540 20828
rect 28592 20816 28598 20868
rect 29638 20816 29644 20868
rect 29696 20856 29702 20868
rect 29892 20859 29950 20865
rect 29892 20856 29904 20859
rect 29696 20828 29904 20856
rect 29696 20816 29702 20828
rect 29892 20825 29904 20828
rect 29938 20825 29950 20859
rect 30113 20856 30141 20896
rect 30282 20884 30288 20936
rect 30340 20924 30346 20936
rect 30377 20927 30435 20933
rect 30377 20924 30389 20927
rect 30340 20896 30389 20924
rect 30340 20884 30346 20896
rect 30377 20893 30389 20896
rect 30423 20893 30435 20927
rect 31113 20927 31171 20933
rect 31113 20924 31125 20927
rect 30377 20887 30435 20893
rect 30484 20896 31125 20924
rect 30484 20856 30512 20896
rect 31113 20893 31125 20896
rect 31159 20924 31171 20927
rect 31294 20924 31300 20936
rect 31159 20896 31300 20924
rect 31159 20893 31171 20896
rect 31113 20887 31171 20893
rect 31294 20884 31300 20896
rect 31352 20884 31358 20936
rect 30834 20856 30840 20868
rect 30113 20828 30512 20856
rect 30795 20828 30840 20856
rect 29892 20819 29950 20825
rect 30834 20816 30840 20828
rect 30892 20816 30898 20868
rect 25958 20788 25964 20800
rect 24964 20760 25964 20788
rect 20956 20748 20962 20760
rect 25958 20748 25964 20760
rect 26016 20748 26022 20800
rect 26050 20748 26056 20800
rect 26108 20788 26114 20800
rect 28626 20788 28632 20800
rect 26108 20760 28632 20788
rect 26108 20748 26114 20760
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 28721 20791 28779 20797
rect 28721 20757 28733 20791
rect 28767 20788 28779 20791
rect 29362 20788 29368 20800
rect 28767 20760 29368 20788
rect 28767 20757 28779 20760
rect 28721 20751 28779 20757
rect 29362 20748 29368 20760
rect 29420 20748 29426 20800
rect 29730 20748 29736 20800
rect 29788 20788 29794 20800
rect 30009 20791 30067 20797
rect 30009 20788 30021 20791
rect 29788 20760 30021 20788
rect 29788 20748 29794 20760
rect 30009 20757 30021 20760
rect 30055 20788 30067 20791
rect 30190 20788 30196 20800
rect 30055 20760 30196 20788
rect 30055 20757 30067 20760
rect 30009 20751 30067 20757
rect 30190 20748 30196 20760
rect 30248 20748 30254 20800
rect 1104 20698 31992 20720
rect 1104 20646 8632 20698
rect 8684 20646 8696 20698
rect 8748 20646 8760 20698
rect 8812 20646 8824 20698
rect 8876 20646 8888 20698
rect 8940 20646 16314 20698
rect 16366 20646 16378 20698
rect 16430 20646 16442 20698
rect 16494 20646 16506 20698
rect 16558 20646 16570 20698
rect 16622 20646 23996 20698
rect 24048 20646 24060 20698
rect 24112 20646 24124 20698
rect 24176 20646 24188 20698
rect 24240 20646 24252 20698
rect 24304 20646 31678 20698
rect 31730 20646 31742 20698
rect 31794 20646 31806 20698
rect 31858 20646 31870 20698
rect 31922 20646 31934 20698
rect 31986 20646 31992 20698
rect 1104 20624 31992 20646
rect 6917 20587 6975 20593
rect 6917 20553 6929 20587
rect 6963 20584 6975 20587
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 6963 20556 7941 20584
rect 6963 20553 6975 20556
rect 6917 20547 6975 20553
rect 7929 20553 7941 20556
rect 7975 20584 7987 20587
rect 8294 20584 8300 20596
rect 7975 20556 8300 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 9858 20584 9864 20596
rect 8404 20556 9864 20584
rect 5905 20519 5963 20525
rect 5905 20485 5917 20519
rect 5951 20516 5963 20519
rect 8404 20516 8432 20556
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 10413 20587 10471 20593
rect 10413 20553 10425 20587
rect 10459 20584 10471 20587
rect 12437 20587 12495 20593
rect 12437 20584 12449 20587
rect 10459 20556 12449 20584
rect 10459 20553 10471 20556
rect 10413 20547 10471 20553
rect 12437 20553 12449 20556
rect 12483 20584 12495 20587
rect 12894 20584 12900 20596
rect 12483 20556 12900 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 12894 20544 12900 20556
rect 12952 20544 12958 20596
rect 13998 20584 14004 20596
rect 13004 20556 14004 20584
rect 5951 20488 8432 20516
rect 5951 20485 5963 20488
rect 5905 20479 5963 20485
rect 9674 20476 9680 20528
rect 9732 20516 9738 20528
rect 13004 20516 13032 20556
rect 13998 20544 14004 20556
rect 14056 20584 14062 20596
rect 14109 20587 14167 20593
rect 14109 20584 14121 20587
rect 14056 20556 14121 20584
rect 14056 20544 14062 20556
rect 14109 20553 14121 20556
rect 14155 20553 14167 20587
rect 14109 20547 14167 20553
rect 16301 20587 16359 20593
rect 16301 20553 16313 20587
rect 16347 20584 16359 20587
rect 16942 20584 16948 20596
rect 16347 20556 16948 20584
rect 16347 20553 16359 20556
rect 16301 20547 16359 20553
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 22370 20584 22376 20596
rect 18012 20556 22376 20584
rect 18012 20544 18018 20556
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 23753 20587 23811 20593
rect 23753 20584 23765 20587
rect 22480 20556 23765 20584
rect 9732 20488 13032 20516
rect 9732 20476 9738 20488
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 9585 20451 9643 20457
rect 9585 20448 9597 20451
rect 8619 20420 9597 20448
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 9585 20417 9597 20420
rect 9631 20448 9643 20451
rect 9950 20448 9956 20460
rect 9631 20420 9956 20448
rect 9631 20417 9643 20420
rect 9585 20411 9643 20417
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 10226 20448 10232 20460
rect 10187 20420 10232 20448
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10413 20451 10471 20457
rect 10413 20417 10425 20451
rect 10459 20448 10471 20451
rect 10594 20448 10600 20460
rect 10459 20420 10600 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 10870 20448 10876 20460
rect 10831 20420 10876 20448
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 11149 20451 11207 20457
rect 11149 20417 11161 20451
rect 11195 20448 11207 20451
rect 11330 20448 11336 20460
rect 11195 20420 11336 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 1578 20380 1584 20392
rect 1539 20352 1584 20380
rect 1578 20340 1584 20352
rect 1636 20340 1642 20392
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 10980 20380 11008 20411
rect 11330 20408 11336 20420
rect 11388 20408 11394 20460
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11716 20380 11744 20411
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 12360 20457 12388 20488
rect 13078 20476 13084 20528
rect 13136 20516 13142 20528
rect 13281 20519 13339 20525
rect 13136 20488 13181 20516
rect 13136 20476 13142 20488
rect 13281 20485 13293 20519
rect 13327 20516 13339 20519
rect 13446 20516 13452 20528
rect 13327 20488 13452 20516
rect 13327 20485 13339 20488
rect 13281 20479 13339 20485
rect 13446 20476 13452 20488
rect 13504 20476 13510 20528
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 13909 20519 13967 20525
rect 13909 20516 13921 20519
rect 13596 20488 13921 20516
rect 13596 20476 13602 20488
rect 13909 20485 13921 20488
rect 13955 20485 13967 20519
rect 13909 20479 13967 20485
rect 14936 20488 16988 20516
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11848 20420 11897 20448
rect 11848 20408 11854 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 12345 20451 12403 20457
rect 12345 20417 12357 20451
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20448 12679 20451
rect 14090 20448 14096 20460
rect 12667 20420 14096 20448
rect 12667 20417 12679 20420
rect 12621 20411 12679 20417
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 14936 20457 14964 20488
rect 14921 20451 14979 20457
rect 14921 20448 14933 20451
rect 14332 20420 14933 20448
rect 14332 20408 14338 20420
rect 14921 20417 14933 20420
rect 14967 20417 14979 20451
rect 14921 20411 14979 20417
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 15712 20420 15761 20448
rect 15712 20408 15718 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 15749 20411 15807 20417
rect 15856 20420 16865 20448
rect 12158 20380 12164 20392
rect 7432 20352 11284 20380
rect 11716 20352 12164 20380
rect 7432 20340 7438 20352
rect 5445 20315 5503 20321
rect 5445 20281 5457 20315
rect 5491 20312 5503 20315
rect 7466 20312 7472 20324
rect 5491 20284 7472 20312
rect 5491 20281 5503 20284
rect 5445 20275 5503 20281
rect 7466 20272 7472 20284
rect 7524 20272 7530 20324
rect 9674 20312 9680 20324
rect 9635 20284 9680 20312
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7650 20244 7656 20256
rect 7423 20216 7656 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 9030 20244 9036 20256
rect 7984 20216 9036 20244
rect 7984 20204 7990 20216
rect 9030 20204 9036 20216
rect 9088 20204 9094 20256
rect 11146 20244 11152 20256
rect 11107 20216 11152 20244
rect 11146 20204 11152 20216
rect 11204 20204 11210 20256
rect 11256 20244 11284 20352
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 13538 20380 13544 20392
rect 12544 20352 13544 20380
rect 11793 20315 11851 20321
rect 11793 20281 11805 20315
rect 11839 20312 11851 20315
rect 12544 20312 12572 20352
rect 13538 20340 13544 20352
rect 13596 20340 13602 20392
rect 13722 20340 13728 20392
rect 13780 20380 13786 20392
rect 14734 20380 14740 20392
rect 13780 20352 14740 20380
rect 13780 20340 13786 20352
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20349 15071 20383
rect 15286 20380 15292 20392
rect 15247 20352 15292 20380
rect 15013 20343 15071 20349
rect 11839 20284 12572 20312
rect 12621 20315 12679 20321
rect 11839 20281 11851 20284
rect 11793 20275 11851 20281
rect 12621 20281 12633 20315
rect 12667 20312 12679 20315
rect 12710 20312 12716 20324
rect 12667 20284 12716 20312
rect 12667 20281 12679 20284
rect 12621 20275 12679 20281
rect 12710 20272 12716 20284
rect 12768 20272 12774 20324
rect 12802 20272 12808 20324
rect 12860 20312 12866 20324
rect 14642 20312 14648 20324
rect 12860 20284 14648 20312
rect 12860 20272 12866 20284
rect 14642 20272 14648 20284
rect 14700 20272 14706 20324
rect 15028 20312 15056 20343
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 15470 20340 15476 20392
rect 15528 20380 15534 20392
rect 15856 20380 15884 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 15528 20352 15884 20380
rect 15528 20340 15534 20352
rect 15930 20340 15936 20392
rect 15988 20380 15994 20392
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 15988 20352 16037 20380
rect 15988 20340 15994 20352
rect 16025 20349 16037 20352
rect 16071 20380 16083 20383
rect 16758 20380 16764 20392
rect 16071 20352 16764 20380
rect 16071 20349 16083 20352
rect 16025 20343 16083 20349
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 16960 20380 16988 20488
rect 17218 20476 17224 20528
rect 17276 20516 17282 20528
rect 17497 20519 17555 20525
rect 17497 20516 17509 20519
rect 17276 20488 17509 20516
rect 17276 20476 17282 20488
rect 17497 20485 17509 20488
rect 17543 20485 17555 20519
rect 17497 20479 17555 20485
rect 17865 20519 17923 20525
rect 17865 20485 17877 20519
rect 17911 20516 17923 20519
rect 18322 20516 18328 20528
rect 17911 20488 18328 20516
rect 17911 20485 17923 20488
rect 17865 20479 17923 20485
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 19150 20516 19156 20528
rect 18708 20488 19156 20516
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 17402 20448 17408 20460
rect 17184 20420 17408 20448
rect 17184 20408 17190 20420
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 17681 20451 17739 20457
rect 17544 20446 17632 20448
rect 17681 20446 17693 20451
rect 17544 20420 17693 20446
rect 17544 20380 17572 20420
rect 17604 20418 17693 20420
rect 17681 20417 17693 20418
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 17773 20451 17831 20457
rect 17773 20417 17785 20451
rect 17819 20448 17831 20451
rect 17819 20420 17908 20448
rect 17819 20417 17831 20420
rect 17773 20411 17831 20417
rect 16960 20352 17572 20380
rect 16206 20312 16212 20324
rect 15028 20284 16212 20312
rect 16206 20272 16212 20284
rect 16264 20272 16270 20324
rect 16945 20315 17003 20321
rect 16945 20281 16957 20315
rect 16991 20312 17003 20315
rect 17402 20312 17408 20324
rect 16991 20284 17408 20312
rect 16991 20281 17003 20284
rect 16945 20275 17003 20281
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 17544 20312 17572 20352
rect 17544 20284 17632 20312
rect 12066 20244 12072 20256
rect 11256 20216 12072 20244
rect 12066 20204 12072 20216
rect 12124 20244 12130 20256
rect 12526 20244 12532 20256
rect 12124 20216 12532 20244
rect 12124 20204 12130 20216
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 12894 20204 12900 20256
rect 12952 20244 12958 20256
rect 13265 20247 13323 20253
rect 13265 20244 13277 20247
rect 12952 20216 13277 20244
rect 12952 20204 12958 20216
rect 13265 20213 13277 20216
rect 13311 20213 13323 20247
rect 13265 20207 13323 20213
rect 13449 20247 13507 20253
rect 13449 20213 13461 20247
rect 13495 20244 13507 20247
rect 13906 20244 13912 20256
rect 13495 20216 13912 20244
rect 13495 20213 13507 20216
rect 13449 20207 13507 20213
rect 13906 20204 13912 20216
rect 13964 20204 13970 20256
rect 14090 20244 14096 20256
rect 14051 20216 14096 20244
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 14277 20247 14335 20253
rect 14277 20213 14289 20247
rect 14323 20244 14335 20247
rect 14458 20244 14464 20256
rect 14323 20216 14464 20244
rect 14323 20213 14335 20216
rect 14277 20207 14335 20213
rect 14458 20204 14464 20216
rect 14516 20244 14522 20256
rect 14826 20244 14832 20256
rect 14516 20216 14832 20244
rect 14516 20204 14522 20216
rect 14826 20204 14832 20216
rect 14884 20204 14890 20256
rect 15010 20204 15016 20256
rect 15068 20244 15074 20256
rect 15841 20247 15899 20253
rect 15841 20244 15853 20247
rect 15068 20216 15853 20244
rect 15068 20204 15074 20216
rect 15841 20213 15853 20216
rect 15887 20244 15899 20247
rect 16022 20244 16028 20256
rect 15887 20216 16028 20244
rect 15887 20213 15899 20216
rect 15841 20207 15899 20213
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 16114 20204 16120 20256
rect 16172 20244 16178 20256
rect 17494 20244 17500 20256
rect 16172 20216 17500 20244
rect 16172 20204 16178 20216
rect 17494 20204 17500 20216
rect 17552 20204 17558 20256
rect 17604 20244 17632 20284
rect 17880 20256 17908 20420
rect 17954 20408 17960 20460
rect 18012 20408 18018 20460
rect 18230 20408 18236 20460
rect 18288 20448 18294 20460
rect 18288 20420 18368 20448
rect 18288 20408 18294 20420
rect 17972 20380 18000 20408
rect 18340 20380 18368 20420
rect 18414 20408 18420 20460
rect 18472 20448 18478 20460
rect 18708 20457 18736 20488
rect 19150 20476 19156 20488
rect 19208 20476 19214 20528
rect 19886 20516 19892 20528
rect 19444 20488 19892 20516
rect 18509 20451 18567 20457
rect 18509 20448 18521 20451
rect 18472 20420 18521 20448
rect 18472 20408 18478 20420
rect 18509 20417 18521 20420
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 19242 20448 19248 20460
rect 18923 20420 19248 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 18800 20380 18828 20411
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 19444 20380 19472 20488
rect 19886 20476 19892 20488
rect 19944 20476 19950 20528
rect 20714 20476 20720 20528
rect 20772 20476 20778 20528
rect 21266 20476 21272 20528
rect 21324 20516 21330 20528
rect 22480 20516 22508 20556
rect 23753 20553 23765 20556
rect 23799 20584 23811 20587
rect 25590 20584 25596 20596
rect 23799 20556 25596 20584
rect 23799 20553 23811 20556
rect 23753 20547 23811 20553
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 26418 20544 26424 20596
rect 26476 20584 26482 20596
rect 29730 20584 29736 20596
rect 26476 20556 29736 20584
rect 26476 20544 26482 20556
rect 29730 20544 29736 20556
rect 29788 20544 29794 20596
rect 21324 20488 22508 20516
rect 21324 20476 21330 20488
rect 25682 20476 25688 20528
rect 25740 20476 25746 20528
rect 26142 20476 26148 20528
rect 26200 20516 26206 20528
rect 27706 20516 27712 20528
rect 26200 20488 27712 20516
rect 26200 20476 26206 20488
rect 27706 20476 27712 20488
rect 27764 20476 27770 20528
rect 29086 20476 29092 20528
rect 29144 20516 29150 20528
rect 29914 20516 29920 20528
rect 29144 20488 29920 20516
rect 29144 20476 29150 20488
rect 29914 20476 29920 20488
rect 29972 20476 29978 20528
rect 30558 20476 30564 20528
rect 30616 20516 30622 20528
rect 32030 20516 32036 20528
rect 30616 20488 32036 20516
rect 30616 20476 30622 20488
rect 17972 20352 18276 20380
rect 18340 20352 18828 20380
rect 18248 20312 18276 20352
rect 18800 20324 18828 20352
rect 18892 20352 19472 20380
rect 19536 20420 19833 20448
rect 18892 20324 18920 20352
rect 18690 20312 18696 20324
rect 18248 20284 18696 20312
rect 18690 20272 18696 20284
rect 18748 20272 18754 20324
rect 18782 20272 18788 20324
rect 18840 20272 18846 20324
rect 18874 20272 18880 20324
rect 18932 20272 18938 20324
rect 19153 20315 19211 20321
rect 19153 20281 19165 20315
rect 19199 20312 19211 20315
rect 19536 20312 19564 20420
rect 19805 20380 19833 20420
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 21910 20448 21916 20460
rect 21692 20420 21916 20448
rect 21692 20408 21698 20420
rect 21910 20408 21916 20420
rect 21968 20408 21974 20460
rect 26513 20451 26571 20457
rect 20806 20380 20812 20392
rect 19805 20352 20812 20380
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 21177 20383 21235 20389
rect 21177 20349 21189 20383
rect 21223 20380 21235 20383
rect 21223 20352 21404 20380
rect 21223 20349 21235 20352
rect 21177 20343 21235 20349
rect 19199 20284 19564 20312
rect 19199 20281 19211 20284
rect 19153 20275 19211 20281
rect 19610 20272 19616 20324
rect 19668 20312 19674 20324
rect 19705 20315 19763 20321
rect 19705 20312 19717 20315
rect 19668 20284 19717 20312
rect 19668 20272 19674 20284
rect 19705 20281 19717 20284
rect 19751 20281 19763 20315
rect 19978 20312 19984 20324
rect 19705 20275 19763 20281
rect 19812 20284 19984 20312
rect 17678 20244 17684 20256
rect 17604 20216 17684 20244
rect 17678 20204 17684 20216
rect 17736 20204 17742 20256
rect 17862 20204 17868 20256
rect 17920 20204 17926 20256
rect 18046 20244 18052 20256
rect 18007 20216 18052 20244
rect 18046 20204 18052 20216
rect 18104 20204 18110 20256
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 19812 20244 19840 20284
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 21376 20312 21404 20352
rect 21450 20340 21456 20392
rect 21508 20380 21514 20392
rect 22005 20383 22063 20389
rect 22005 20380 22017 20383
rect 21508 20352 22017 20380
rect 21508 20340 21514 20352
rect 22005 20349 22017 20352
rect 22051 20380 22063 20383
rect 22278 20380 22284 20392
rect 22051 20349 22072 20380
rect 22239 20352 22284 20380
rect 22005 20343 22072 20349
rect 21634 20312 21640 20324
rect 21376 20284 21640 20312
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 18288 20216 19840 20244
rect 18288 20204 18294 20216
rect 19886 20204 19892 20256
rect 19944 20244 19950 20256
rect 21542 20244 21548 20256
rect 19944 20216 21548 20244
rect 19944 20204 19950 20216
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 22044 20244 22072 20343
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 22370 20340 22376 20392
rect 22428 20380 22434 20392
rect 23400 20380 23428 20434
rect 26513 20417 26525 20451
rect 26559 20448 26571 20451
rect 26694 20448 26700 20460
rect 26559 20420 26700 20448
rect 26559 20417 26571 20420
rect 26513 20411 26571 20417
rect 26694 20408 26700 20420
rect 26752 20448 26758 20460
rect 26970 20448 26976 20460
rect 26752 20420 26976 20448
rect 26752 20408 26758 20420
rect 26970 20408 26976 20420
rect 27028 20408 27034 20460
rect 27157 20451 27215 20457
rect 27157 20417 27169 20451
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 22428 20352 23428 20380
rect 22428 20340 22434 20352
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 25866 20380 25872 20392
rect 23532 20352 25872 20380
rect 23532 20340 23538 20352
rect 25866 20340 25872 20352
rect 25924 20340 25930 20392
rect 26237 20383 26295 20389
rect 26237 20349 26249 20383
rect 26283 20380 26295 20383
rect 26283 20352 26556 20380
rect 26283 20349 26295 20352
rect 26237 20343 26295 20349
rect 23750 20272 23756 20324
rect 23808 20312 23814 20324
rect 24765 20315 24823 20321
rect 24765 20312 24777 20315
rect 23808 20284 24777 20312
rect 23808 20272 23814 20284
rect 24765 20281 24777 20284
rect 24811 20281 24823 20315
rect 24765 20275 24823 20281
rect 22738 20244 22744 20256
rect 22044 20216 22744 20244
rect 22738 20204 22744 20216
rect 22796 20204 22802 20256
rect 24780 20244 24808 20275
rect 25774 20244 25780 20256
rect 24780 20216 25780 20244
rect 25774 20204 25780 20216
rect 25832 20204 25838 20256
rect 26528 20244 26556 20352
rect 26602 20340 26608 20392
rect 26660 20380 26666 20392
rect 27172 20380 27200 20411
rect 28534 20408 28540 20460
rect 28592 20408 28598 20460
rect 28810 20408 28816 20460
rect 28868 20448 28874 20460
rect 29454 20448 29460 20460
rect 28868 20420 29460 20448
rect 28868 20408 28874 20420
rect 29454 20408 29460 20420
rect 29512 20408 29518 20460
rect 30760 20457 30788 20488
rect 32030 20476 32036 20488
rect 32088 20476 32094 20528
rect 29825 20451 29883 20457
rect 29825 20417 29837 20451
rect 29871 20417 29883 20451
rect 29825 20411 29883 20417
rect 30653 20451 30711 20457
rect 30653 20417 30665 20451
rect 30699 20417 30711 20451
rect 30653 20411 30711 20417
rect 30745 20451 30803 20457
rect 30745 20417 30757 20451
rect 30791 20417 30803 20451
rect 30745 20411 30803 20417
rect 26660 20352 27200 20380
rect 27433 20383 27491 20389
rect 26660 20340 26666 20352
rect 27433 20349 27445 20383
rect 27479 20380 27491 20383
rect 27522 20380 27528 20392
rect 27479 20352 27528 20380
rect 27479 20349 27491 20352
rect 27433 20343 27491 20349
rect 27522 20340 27528 20352
rect 27580 20340 27586 20392
rect 27890 20340 27896 20392
rect 27948 20380 27954 20392
rect 27948 20352 28488 20380
rect 27948 20340 27954 20352
rect 28460 20312 28488 20352
rect 28718 20340 28724 20392
rect 28776 20380 28782 20392
rect 29638 20380 29644 20392
rect 28776 20352 29644 20380
rect 28776 20340 28782 20352
rect 29638 20340 29644 20352
rect 29696 20340 29702 20392
rect 29457 20315 29515 20321
rect 29457 20312 29469 20315
rect 28460 20284 29469 20312
rect 29457 20281 29469 20284
rect 29503 20281 29515 20315
rect 29840 20312 29868 20411
rect 29917 20383 29975 20389
rect 29917 20349 29929 20383
rect 29963 20380 29975 20383
rect 30558 20380 30564 20392
rect 29963 20352 30564 20380
rect 29963 20349 29975 20352
rect 29917 20343 29975 20349
rect 30558 20340 30564 20352
rect 30616 20340 30622 20392
rect 30006 20312 30012 20324
rect 29840 20284 30012 20312
rect 29457 20275 29515 20281
rect 30006 20272 30012 20284
rect 30064 20312 30070 20324
rect 30668 20312 30696 20411
rect 30834 20408 30840 20460
rect 30892 20448 30898 20460
rect 31021 20451 31079 20457
rect 31021 20448 31033 20451
rect 30892 20420 31033 20448
rect 30892 20408 30898 20420
rect 31021 20417 31033 20420
rect 31067 20448 31079 20451
rect 31570 20448 31576 20460
rect 31067 20420 31576 20448
rect 31067 20417 31079 20420
rect 31021 20411 31079 20417
rect 31570 20408 31576 20420
rect 31628 20408 31634 20460
rect 32858 20408 32864 20460
rect 32916 20448 32922 20460
rect 32916 20420 32996 20448
rect 32916 20408 32922 20420
rect 30926 20380 30932 20392
rect 30887 20352 30932 20380
rect 30926 20340 30932 20352
rect 30984 20340 30990 20392
rect 32858 20312 32864 20324
rect 30064 20284 30604 20312
rect 30668 20284 32864 20312
rect 30064 20272 30070 20284
rect 28718 20244 28724 20256
rect 26528 20216 28724 20244
rect 28718 20204 28724 20216
rect 28776 20204 28782 20256
rect 28905 20247 28963 20253
rect 28905 20213 28917 20247
rect 28951 20244 28963 20247
rect 30282 20244 30288 20256
rect 28951 20216 30288 20244
rect 28951 20213 28963 20216
rect 28905 20207 28963 20213
rect 30282 20204 30288 20216
rect 30340 20204 30346 20256
rect 30466 20244 30472 20256
rect 30427 20216 30472 20244
rect 30466 20204 30472 20216
rect 30524 20204 30530 20256
rect 30576 20244 30604 20284
rect 32858 20272 32864 20284
rect 32916 20272 32922 20324
rect 32582 20244 32588 20256
rect 30576 20216 32588 20244
rect 32582 20204 32588 20216
rect 32640 20204 32646 20256
rect 1104 20154 31832 20176
rect 1104 20102 4791 20154
rect 4843 20102 4855 20154
rect 4907 20102 4919 20154
rect 4971 20102 4983 20154
rect 5035 20102 5047 20154
rect 5099 20102 12473 20154
rect 12525 20102 12537 20154
rect 12589 20102 12601 20154
rect 12653 20102 12665 20154
rect 12717 20102 12729 20154
rect 12781 20102 20155 20154
rect 20207 20102 20219 20154
rect 20271 20102 20283 20154
rect 20335 20102 20347 20154
rect 20399 20102 20411 20154
rect 20463 20102 27837 20154
rect 27889 20102 27901 20154
rect 27953 20102 27965 20154
rect 28017 20102 28029 20154
rect 28081 20102 28093 20154
rect 28145 20102 31832 20154
rect 32858 20136 32864 20188
rect 32916 20176 32922 20188
rect 32968 20176 32996 20420
rect 32916 20148 32996 20176
rect 32916 20136 32922 20148
rect 1104 20080 31832 20102
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 7984 20012 8493 20040
rect 7984 20000 7990 20012
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 8481 20003 8539 20009
rect 10597 20043 10655 20049
rect 10597 20009 10609 20043
rect 10643 20040 10655 20043
rect 10643 20012 12112 20040
rect 10643 20009 10655 20012
rect 10597 20003 10655 20009
rect 11425 19975 11483 19981
rect 11425 19941 11437 19975
rect 11471 19972 11483 19975
rect 11514 19972 11520 19984
rect 11471 19944 11520 19972
rect 11471 19941 11483 19944
rect 11425 19935 11483 19941
rect 11514 19932 11520 19944
rect 11572 19932 11578 19984
rect 11885 19975 11943 19981
rect 11885 19941 11897 19975
rect 11931 19972 11943 19975
rect 11974 19972 11980 19984
rect 11931 19944 11980 19972
rect 11931 19941 11943 19944
rect 11885 19935 11943 19941
rect 11974 19932 11980 19944
rect 12032 19932 12038 19984
rect 12084 19972 12112 20012
rect 12158 20000 12164 20052
rect 12216 20040 12222 20052
rect 13722 20040 13728 20052
rect 12216 20012 13308 20040
rect 13683 20012 13728 20040
rect 12216 20000 12222 20012
rect 13170 19972 13176 19984
rect 12084 19944 13176 19972
rect 13170 19932 13176 19944
rect 13228 19932 13234 19984
rect 13280 19972 13308 20012
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 13964 20012 18184 20040
rect 13964 20000 13970 20012
rect 14274 19972 14280 19984
rect 13280 19944 14280 19972
rect 14274 19932 14280 19944
rect 14332 19932 14338 19984
rect 14461 19975 14519 19981
rect 14461 19941 14473 19975
rect 14507 19972 14519 19975
rect 17954 19972 17960 19984
rect 14507 19944 17960 19972
rect 14507 19941 14519 19944
rect 14461 19935 14519 19941
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 18156 19972 18184 20012
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 19702 20040 19708 20052
rect 18288 20012 19708 20040
rect 18288 20000 18294 20012
rect 19702 20000 19708 20012
rect 19760 20000 19766 20052
rect 19805 20012 21588 20040
rect 18156 19944 18644 19972
rect 10870 19904 10876 19916
rect 7944 19876 10876 19904
rect 7944 19848 7972 19876
rect 10870 19864 10876 19876
rect 10928 19904 10934 19916
rect 10928 19876 12204 19904
rect 10928 19864 10934 19876
rect 7466 19836 7472 19848
rect 7379 19808 7472 19836
rect 7466 19796 7472 19808
rect 7524 19836 7530 19848
rect 7926 19836 7932 19848
rect 7524 19808 7932 19836
rect 7524 19796 7530 19808
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 10226 19796 10232 19848
rect 10284 19836 10290 19848
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 10284 19808 10517 19836
rect 10284 19796 10290 19808
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 6365 19771 6423 19777
rect 6365 19737 6377 19771
rect 6411 19768 6423 19771
rect 8018 19768 8024 19780
rect 6411 19740 8024 19768
rect 6411 19737 6423 19740
rect 6365 19731 6423 19737
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 9493 19771 9551 19777
rect 9493 19737 9505 19771
rect 9539 19768 9551 19771
rect 9858 19768 9864 19780
rect 9539 19740 9864 19768
rect 9539 19737 9551 19740
rect 9493 19731 9551 19737
rect 9858 19728 9864 19740
rect 9916 19728 9922 19780
rect 10520 19768 10548 19799
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 11164 19845 11192 19876
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 10652 19808 10701 19836
rect 10652 19796 10658 19808
rect 10689 19805 10701 19808
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 11149 19839 11207 19845
rect 11149 19805 11161 19839
rect 11195 19805 11207 19839
rect 11149 19799 11207 19805
rect 11425 19839 11483 19845
rect 11425 19805 11437 19839
rect 11471 19805 11483 19839
rect 11425 19799 11483 19805
rect 11440 19768 11468 19799
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 11885 19839 11943 19845
rect 11885 19836 11897 19839
rect 11572 19808 11897 19836
rect 11572 19796 11578 19808
rect 11885 19805 11897 19808
rect 11931 19805 11943 19839
rect 12066 19836 12072 19848
rect 12027 19808 12072 19836
rect 11885 19799 11943 19805
rect 12066 19796 12072 19808
rect 12124 19796 12130 19848
rect 12176 19845 12204 19876
rect 12342 19864 12348 19916
rect 12400 19904 12406 19916
rect 13630 19904 13636 19916
rect 12400 19876 13636 19904
rect 12400 19864 12406 19876
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 16206 19904 16212 19916
rect 13872 19876 16068 19904
rect 16167 19876 16212 19904
rect 13872 19864 13878 19876
rect 12161 19839 12219 19845
rect 12161 19805 12173 19839
rect 12207 19836 12219 19839
rect 12250 19836 12256 19848
rect 12207 19808 12256 19836
rect 12207 19805 12219 19808
rect 12161 19799 12219 19805
rect 12250 19796 12256 19808
rect 12308 19796 12314 19848
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 13262 19836 13268 19848
rect 12676 19808 13268 19836
rect 12676 19796 12682 19808
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 13504 19808 13553 19836
rect 13504 19796 13510 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19836 13783 19839
rect 14274 19836 14280 19848
rect 13771 19808 14280 19836
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 14734 19836 14740 19848
rect 14476 19808 14740 19836
rect 12084 19768 12112 19796
rect 12710 19768 12716 19780
rect 10520 19740 11376 19768
rect 11440 19740 12112 19768
rect 12671 19740 12716 19768
rect 6914 19700 6920 19712
rect 6875 19672 6920 19700
rect 6914 19660 6920 19672
rect 6972 19700 6978 19712
rect 7374 19700 7380 19712
rect 6972 19672 7380 19700
rect 6972 19660 6978 19672
rect 7374 19660 7380 19672
rect 7432 19700 7438 19712
rect 7929 19703 7987 19709
rect 7929 19700 7941 19703
rect 7432 19672 7941 19700
rect 7432 19660 7438 19672
rect 7929 19669 7941 19672
rect 7975 19669 7987 19703
rect 9950 19700 9956 19712
rect 9911 19672 9956 19700
rect 7929 19663 7987 19669
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 11238 19700 11244 19712
rect 11199 19672 11244 19700
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 11348 19700 11376 19740
rect 12710 19728 12716 19740
rect 12768 19728 12774 19780
rect 12986 19728 12992 19780
rect 13044 19768 13050 19780
rect 14476 19768 14504 19808
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 14884 19808 14929 19836
rect 14884 19796 14890 19808
rect 15010 19796 15016 19848
rect 15068 19836 15074 19848
rect 15470 19836 15476 19848
rect 15068 19808 15476 19836
rect 15068 19796 15074 19808
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 15562 19796 15568 19848
rect 15620 19836 15626 19848
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 15620 19808 15761 19836
rect 15620 19796 15626 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 16040 19836 16068 19876
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19904 16727 19907
rect 17218 19904 17224 19916
rect 16715 19876 17224 19904
rect 16715 19873 16727 19876
rect 16669 19867 16727 19873
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 17328 19876 17509 19904
rect 16577 19839 16635 19845
rect 16577 19836 16589 19839
rect 16040 19808 16589 19836
rect 15749 19799 15807 19805
rect 16577 19805 16589 19808
rect 16623 19836 16635 19839
rect 17126 19836 17132 19848
rect 16623 19808 17132 19836
rect 16623 19805 16635 19808
rect 16577 19799 16635 19805
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 13044 19740 14504 19768
rect 13044 19728 13050 19740
rect 14642 19728 14648 19780
rect 14700 19768 14706 19780
rect 15102 19768 15108 19780
rect 14700 19740 15108 19768
rect 14700 19728 14706 19740
rect 15102 19728 15108 19740
rect 15160 19768 15166 19780
rect 15654 19768 15660 19780
rect 15160 19740 15660 19768
rect 15160 19728 15166 19740
rect 15654 19728 15660 19740
rect 15712 19768 15718 19780
rect 17328 19768 17356 19876
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 17773 19907 17831 19913
rect 17773 19904 17785 19907
rect 17497 19867 17555 19873
rect 17696 19876 17785 19904
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 15712 19740 17356 19768
rect 15712 19728 15718 19740
rect 17420 19712 17448 19799
rect 17512 19768 17540 19867
rect 17696 19848 17724 19876
rect 17773 19873 17785 19876
rect 17819 19904 17831 19907
rect 18616 19904 18644 19944
rect 18690 19932 18696 19984
rect 18748 19972 18754 19984
rect 19805 19972 19833 20012
rect 18748 19944 19833 19972
rect 21560 19972 21588 20012
rect 21634 20000 21640 20052
rect 21692 20040 21698 20052
rect 22557 20043 22615 20049
rect 22557 20040 22569 20043
rect 21692 20012 22569 20040
rect 21692 20000 21698 20012
rect 22557 20009 22569 20012
rect 22603 20009 22615 20043
rect 22557 20003 22615 20009
rect 23014 20000 23020 20052
rect 23072 20040 23078 20052
rect 25038 20040 25044 20052
rect 23072 20012 25044 20040
rect 23072 20000 23078 20012
rect 25038 20000 25044 20012
rect 25096 20000 25102 20052
rect 25314 20000 25320 20052
rect 25372 20040 25378 20052
rect 26510 20040 26516 20052
rect 25372 20012 26516 20040
rect 25372 20000 25378 20012
rect 26510 20000 26516 20012
rect 26568 20000 26574 20052
rect 26786 20000 26792 20052
rect 26844 20040 26850 20052
rect 26881 20043 26939 20049
rect 26881 20040 26893 20043
rect 26844 20012 26893 20040
rect 26844 20000 26850 20012
rect 26881 20009 26893 20012
rect 26927 20009 26939 20043
rect 27706 20040 27712 20052
rect 26881 20003 26939 20009
rect 26977 20012 27712 20040
rect 21910 19972 21916 19984
rect 21560 19944 21916 19972
rect 18748 19932 18754 19944
rect 21910 19932 21916 19944
rect 21968 19932 21974 19984
rect 22462 19932 22468 19984
rect 22520 19972 22526 19984
rect 23474 19972 23480 19984
rect 22520 19944 23480 19972
rect 22520 19932 22526 19944
rect 23474 19932 23480 19944
rect 23532 19932 23538 19984
rect 26142 19932 26148 19984
rect 26200 19972 26206 19984
rect 26977 19972 27005 20012
rect 27706 20000 27712 20012
rect 27764 20000 27770 20052
rect 28994 20040 29000 20052
rect 28173 20012 29000 20040
rect 26200 19944 27005 19972
rect 26200 19932 26206 19944
rect 27430 19932 27436 19984
rect 27488 19972 27494 19984
rect 28173 19972 28201 20012
rect 28994 20000 29000 20012
rect 29052 20000 29058 20052
rect 30834 20040 30840 20052
rect 29104 20012 30840 20040
rect 29104 19972 29132 20012
rect 30834 20000 30840 20012
rect 30892 20000 30898 20052
rect 31110 19972 31116 19984
rect 27488 19944 27533 19972
rect 27632 19944 28201 19972
rect 28736 19944 29132 19972
rect 29932 19944 31116 19972
rect 27488 19932 27494 19944
rect 23201 19907 23259 19913
rect 23201 19904 23213 19907
rect 17819 19876 18552 19904
rect 18616 19876 23213 19904
rect 17819 19873 17831 19876
rect 17773 19867 17831 19873
rect 17678 19796 17684 19848
rect 17736 19796 17742 19848
rect 18138 19796 18144 19848
rect 18196 19833 18202 19848
rect 18524 19845 18552 19876
rect 23201 19873 23213 19876
rect 23247 19873 23259 19907
rect 23750 19904 23756 19916
rect 23201 19867 23259 19873
rect 23308 19876 23756 19904
rect 18233 19839 18291 19845
rect 18233 19833 18245 19839
rect 18196 19805 18245 19833
rect 18279 19805 18291 19839
rect 18196 19796 18202 19805
rect 18233 19799 18291 19805
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 18966 19836 18972 19848
rect 18647 19808 18972 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 17512 19740 17815 19768
rect 12526 19700 12532 19712
rect 11348 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 12802 19700 12808 19712
rect 12763 19672 12808 19700
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 13357 19703 13415 19709
rect 13357 19669 13369 19703
rect 13403 19700 13415 19703
rect 13630 19700 13636 19712
rect 13403 19672 13636 19700
rect 13403 19669 13415 19672
rect 13357 19663 13415 19669
rect 13630 19660 13636 19672
rect 13688 19700 13694 19712
rect 14182 19700 14188 19712
rect 13688 19672 14188 19700
rect 13688 19660 13694 19672
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 14274 19660 14280 19712
rect 14332 19700 14338 19712
rect 15930 19700 15936 19712
rect 14332 19672 15936 19700
rect 14332 19660 14338 19672
rect 15930 19660 15936 19672
rect 15988 19660 15994 19712
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 17402 19700 17408 19712
rect 16080 19672 17408 19700
rect 16080 19660 16086 19672
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 17787 19700 17815 19740
rect 17954 19728 17960 19780
rect 18012 19768 18018 19780
rect 18432 19768 18460 19799
rect 18966 19796 18972 19808
rect 19024 19796 19030 19848
rect 19426 19836 19432 19848
rect 19387 19808 19432 19836
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 20073 19839 20131 19845
rect 20073 19836 20085 19839
rect 19812 19808 20085 19836
rect 18012 19740 18460 19768
rect 18012 19728 18018 19740
rect 18690 19728 18696 19780
rect 18748 19768 18754 19780
rect 19702 19768 19708 19780
rect 18748 19740 19708 19768
rect 18748 19728 18754 19740
rect 19702 19728 19708 19740
rect 19760 19768 19766 19780
rect 19812 19768 19840 19808
rect 20073 19805 20085 19808
rect 20119 19805 20131 19839
rect 22738 19836 22744 19848
rect 22699 19808 22744 19836
rect 20073 19799 20131 19805
rect 22738 19796 22744 19808
rect 22796 19796 22802 19848
rect 22830 19796 22836 19848
rect 22888 19836 22894 19848
rect 23308 19836 23336 19876
rect 23750 19864 23756 19876
rect 23808 19864 23814 19916
rect 24854 19864 24860 19916
rect 24912 19904 24918 19916
rect 26329 19907 26387 19913
rect 24912 19876 26280 19904
rect 24912 19864 24918 19876
rect 22888 19808 23336 19836
rect 22888 19796 22894 19808
rect 23382 19796 23388 19848
rect 23440 19836 23446 19848
rect 23477 19839 23535 19845
rect 23477 19836 23489 19839
rect 23440 19808 23489 19836
rect 23440 19796 23446 19808
rect 23477 19805 23489 19808
rect 23523 19805 23535 19839
rect 24578 19836 24584 19848
rect 24539 19808 24584 19836
rect 23477 19799 23535 19805
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 26252 19836 26280 19876
rect 26329 19873 26341 19907
rect 26375 19904 26387 19907
rect 26418 19904 26424 19916
rect 26375 19876 26424 19904
rect 26375 19873 26387 19876
rect 26329 19867 26387 19873
rect 26418 19864 26424 19876
rect 26476 19864 26482 19916
rect 26878 19864 26884 19916
rect 26936 19904 26942 19916
rect 27249 19907 27307 19913
rect 27249 19904 27261 19907
rect 26936 19876 27261 19904
rect 26936 19864 26942 19876
rect 27249 19873 27261 19876
rect 27295 19873 27307 19907
rect 27249 19867 27307 19873
rect 27341 19907 27399 19913
rect 27341 19873 27353 19907
rect 27387 19904 27399 19907
rect 27632 19904 27660 19944
rect 27387 19876 27660 19904
rect 27387 19873 27399 19876
rect 27341 19867 27399 19873
rect 27706 19864 27712 19916
rect 27764 19904 27770 19916
rect 28736 19913 28764 19944
rect 28629 19907 28687 19913
rect 28629 19904 28641 19907
rect 27764 19876 28641 19904
rect 27764 19864 27770 19876
rect 28629 19873 28641 19876
rect 28675 19873 28687 19907
rect 28629 19867 28687 19873
rect 28721 19907 28779 19913
rect 28721 19873 28733 19907
rect 28767 19873 28779 19907
rect 28721 19867 28779 19873
rect 26786 19836 26792 19848
rect 26252 19808 26792 19836
rect 26786 19796 26792 19808
rect 26844 19836 26850 19848
rect 27157 19839 27215 19845
rect 27157 19836 27169 19839
rect 26844 19808 27169 19836
rect 26844 19796 26850 19808
rect 27157 19805 27169 19808
rect 27203 19805 27215 19839
rect 27617 19839 27675 19845
rect 27157 19799 27215 19805
rect 27264 19808 27568 19836
rect 19760 19740 19840 19768
rect 19760 19728 19766 19740
rect 19886 19728 19892 19780
rect 19944 19728 19950 19780
rect 20254 19728 20260 19780
rect 20312 19768 20318 19780
rect 20349 19771 20407 19777
rect 20349 19768 20361 19771
rect 20312 19740 20361 19768
rect 20312 19728 20318 19740
rect 20349 19737 20361 19740
rect 20395 19737 20407 19771
rect 22094 19768 22100 19780
rect 21574 19740 21680 19768
rect 22055 19740 22100 19768
rect 20349 19731 20407 19737
rect 18506 19700 18512 19712
rect 17787 19672 18512 19700
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 18877 19703 18935 19709
rect 18877 19669 18889 19703
rect 18923 19700 18935 19703
rect 19334 19700 19340 19712
rect 18923 19672 19340 19700
rect 18923 19669 18935 19672
rect 18877 19663 18935 19669
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 19613 19703 19671 19709
rect 19613 19669 19625 19703
rect 19659 19700 19671 19703
rect 19794 19700 19800 19712
rect 19659 19672 19800 19700
rect 19659 19669 19671 19672
rect 19613 19663 19671 19669
rect 19794 19660 19800 19672
rect 19852 19660 19858 19712
rect 19904 19700 19932 19728
rect 21358 19700 21364 19712
rect 19904 19672 21364 19700
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 21652 19700 21680 19740
rect 22094 19728 22100 19740
rect 22152 19768 22158 19780
rect 22848 19768 22876 19796
rect 22152 19740 22876 19768
rect 22152 19728 22158 19740
rect 22922 19728 22928 19780
rect 22980 19768 22986 19780
rect 24854 19768 24860 19780
rect 22980 19740 24716 19768
rect 24815 19740 24860 19768
rect 22980 19728 22986 19740
rect 23290 19700 23296 19712
rect 21652 19672 23296 19700
rect 23290 19660 23296 19672
rect 23348 19660 23354 19712
rect 24688 19700 24716 19740
rect 24854 19728 24860 19740
rect 24912 19728 24918 19780
rect 25866 19728 25872 19780
rect 25924 19728 25930 19780
rect 26510 19728 26516 19780
rect 26568 19768 26574 19780
rect 27264 19768 27292 19808
rect 26568 19740 27292 19768
rect 27540 19768 27568 19808
rect 27617 19805 27629 19839
rect 27663 19836 27675 19839
rect 27890 19836 27896 19848
rect 27663 19808 27896 19836
rect 27663 19805 27675 19808
rect 27617 19799 27675 19805
rect 27890 19796 27896 19808
rect 27948 19796 27954 19848
rect 29932 19845 29960 19944
rect 31110 19932 31116 19944
rect 31168 19932 31174 19984
rect 30190 19904 30196 19916
rect 30151 19876 30196 19904
rect 30190 19864 30196 19876
rect 30248 19864 30254 19916
rect 30742 19904 30748 19916
rect 30703 19876 30748 19904
rect 30742 19864 30748 19876
rect 30800 19864 30806 19916
rect 31205 19907 31263 19913
rect 31205 19873 31217 19907
rect 31251 19904 31263 19907
rect 31570 19904 31576 19916
rect 31251 19876 31576 19904
rect 31251 19873 31263 19876
rect 31205 19867 31263 19873
rect 31570 19864 31576 19876
rect 31628 19864 31634 19916
rect 28258 19839 28316 19845
rect 28258 19805 28270 19839
rect 28304 19836 28316 19839
rect 29917 19839 29975 19845
rect 29917 19836 29929 19839
rect 28304 19808 29929 19836
rect 28304 19805 28316 19808
rect 28258 19799 28316 19805
rect 29917 19805 29929 19808
rect 29963 19805 29975 19839
rect 29917 19799 29975 19805
rect 30009 19839 30067 19845
rect 30009 19805 30021 19839
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 30285 19839 30343 19845
rect 30285 19805 30297 19839
rect 30331 19836 30343 19839
rect 30466 19836 30472 19848
rect 30331 19808 30472 19836
rect 30331 19805 30343 19808
rect 30285 19799 30343 19805
rect 27540 19740 28120 19768
rect 26568 19728 26574 19740
rect 27246 19700 27252 19712
rect 24688 19672 27252 19700
rect 27246 19660 27252 19672
rect 27304 19660 27310 19712
rect 28092 19709 28120 19740
rect 29730 19728 29736 19780
rect 29788 19768 29794 19780
rect 29788 19740 29833 19768
rect 29788 19728 29794 19740
rect 30024 19712 30052 19799
rect 30466 19796 30472 19808
rect 30524 19796 30530 19848
rect 31110 19836 31116 19848
rect 31071 19808 31116 19836
rect 31110 19796 31116 19808
rect 31168 19796 31174 19848
rect 28077 19703 28135 19709
rect 28077 19669 28089 19703
rect 28123 19669 28135 19703
rect 28258 19700 28264 19712
rect 28219 19672 28264 19700
rect 28077 19663 28135 19669
rect 28258 19660 28264 19672
rect 28316 19700 28322 19712
rect 30006 19700 30012 19712
rect 28316 19672 30012 19700
rect 28316 19660 28322 19672
rect 30006 19660 30012 19672
rect 30064 19660 30070 19712
rect 30282 19660 30288 19712
rect 30340 19700 30346 19712
rect 30466 19700 30472 19712
rect 30340 19672 30472 19700
rect 30340 19660 30346 19672
rect 30466 19660 30472 19672
rect 30524 19660 30530 19712
rect 1104 19610 31992 19632
rect 1104 19558 8632 19610
rect 8684 19558 8696 19610
rect 8748 19558 8760 19610
rect 8812 19558 8824 19610
rect 8876 19558 8888 19610
rect 8940 19558 16314 19610
rect 16366 19558 16378 19610
rect 16430 19558 16442 19610
rect 16494 19558 16506 19610
rect 16558 19558 16570 19610
rect 16622 19558 23996 19610
rect 24048 19558 24060 19610
rect 24112 19558 24124 19610
rect 24176 19558 24188 19610
rect 24240 19558 24252 19610
rect 24304 19558 31678 19610
rect 31730 19558 31742 19610
rect 31794 19558 31806 19610
rect 31858 19558 31870 19610
rect 31922 19558 31934 19610
rect 31986 19558 31992 19610
rect 1104 19536 31992 19558
rect 9030 19456 9036 19508
rect 9088 19496 9094 19508
rect 9953 19499 10011 19505
rect 9953 19496 9965 19499
rect 9088 19468 9965 19496
rect 9088 19456 9094 19468
rect 9953 19465 9965 19468
rect 9999 19496 10011 19499
rect 11422 19496 11428 19508
rect 9999 19468 11428 19496
rect 9999 19465 10011 19468
rect 9953 19459 10011 19465
rect 11422 19456 11428 19468
rect 11480 19496 11486 19508
rect 12158 19496 12164 19508
rect 11480 19468 12164 19496
rect 11480 19456 11486 19468
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 12798 19499 12856 19505
rect 12798 19465 12810 19499
rect 12844 19496 12856 19499
rect 13262 19496 13268 19508
rect 12844 19468 13268 19496
rect 12844 19465 12856 19468
rect 12798 19459 12856 19465
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 14090 19456 14096 19508
rect 14148 19496 14154 19508
rect 14461 19499 14519 19505
rect 14461 19496 14473 19499
rect 14148 19468 14473 19496
rect 14148 19456 14154 19468
rect 14461 19465 14473 19468
rect 14507 19496 14519 19499
rect 16758 19496 16764 19508
rect 14507 19468 16764 19496
rect 14507 19465 14519 19468
rect 14461 19459 14519 19465
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 16942 19456 16948 19508
rect 17000 19496 17006 19508
rect 17954 19496 17960 19508
rect 17000 19468 17960 19496
rect 17000 19456 17006 19468
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 18049 19499 18107 19505
rect 18049 19465 18061 19499
rect 18095 19496 18107 19499
rect 18874 19496 18880 19508
rect 18095 19468 18880 19496
rect 18095 19465 18107 19468
rect 18049 19459 18107 19465
rect 18874 19456 18880 19468
rect 18932 19456 18938 19508
rect 19150 19496 19156 19508
rect 19111 19468 19156 19496
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 19610 19496 19616 19508
rect 19536 19468 19616 19496
rect 8018 19388 8024 19440
rect 8076 19428 8082 19440
rect 9490 19428 9496 19440
rect 8076 19400 9496 19428
rect 8076 19388 8082 19400
rect 9490 19388 9496 19400
rect 9548 19428 9554 19440
rect 11330 19428 11336 19440
rect 9548 19400 11336 19428
rect 9548 19388 9554 19400
rect 11330 19388 11336 19400
rect 11388 19428 11394 19440
rect 11514 19428 11520 19440
rect 11388 19400 11520 19428
rect 11388 19388 11394 19400
rect 11514 19388 11520 19400
rect 11572 19388 11578 19440
rect 11698 19388 11704 19440
rect 11756 19388 11762 19440
rect 12066 19428 12072 19440
rect 12027 19400 12072 19428
rect 12066 19388 12072 19400
rect 12124 19388 12130 19440
rect 12526 19428 12532 19440
rect 12268 19400 12532 19428
rect 10870 19320 10876 19372
rect 10928 19360 10934 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10928 19332 10977 19360
rect 10928 19320 10934 19332
rect 10965 19329 10977 19332
rect 11011 19329 11023 19363
rect 10965 19323 11023 19329
rect 7193 19295 7251 19301
rect 7193 19261 7205 19295
rect 7239 19292 7251 19295
rect 9582 19292 9588 19304
rect 7239 19264 9588 19292
rect 7239 19261 7251 19264
rect 7193 19255 7251 19261
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 10042 19252 10048 19304
rect 10100 19292 10106 19304
rect 10980 19292 11008 19323
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11716 19360 11744 19388
rect 11977 19363 12035 19369
rect 11977 19360 11989 19363
rect 11112 19332 11157 19360
rect 11256 19332 11989 19360
rect 11112 19320 11118 19332
rect 11256 19292 11284 19332
rect 11977 19329 11989 19332
rect 12023 19360 12035 19363
rect 12268 19360 12296 19400
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 12894 19428 12900 19440
rect 12855 19400 12900 19428
rect 12894 19388 12900 19400
rect 12952 19388 12958 19440
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 13357 19431 13415 19437
rect 13357 19428 13369 19431
rect 13228 19400 13369 19428
rect 13228 19388 13234 19400
rect 13357 19397 13369 19400
rect 13403 19397 13415 19431
rect 13357 19391 13415 19397
rect 12023 19332 12296 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12618 19360 12624 19372
rect 12400 19332 12624 19360
rect 12400 19320 12406 19332
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 12802 19360 12808 19372
rect 12759 19332 12808 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 12802 19320 12808 19332
rect 12860 19360 12866 19372
rect 13078 19360 13084 19372
rect 12860 19332 13084 19360
rect 12860 19320 12866 19332
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 10100 19264 11284 19292
rect 10100 19252 10106 19264
rect 11330 19252 11336 19304
rect 11388 19292 11394 19304
rect 12894 19292 12900 19304
rect 11388 19264 12900 19292
rect 11388 19252 11394 19264
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 13170 19252 13176 19304
rect 13228 19292 13234 19304
rect 13372 19292 13400 19391
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 15749 19431 15807 19437
rect 15749 19428 15761 19431
rect 13780 19400 15761 19428
rect 13780 19388 13786 19400
rect 15749 19397 15761 19400
rect 15795 19428 15807 19431
rect 17310 19428 17316 19440
rect 15795 19400 17316 19428
rect 15795 19397 15807 19400
rect 15749 19391 15807 19397
rect 17310 19388 17316 19400
rect 17368 19388 17374 19440
rect 17402 19388 17408 19440
rect 17460 19428 17466 19440
rect 18414 19428 18420 19440
rect 17460 19400 18420 19428
rect 17460 19388 17466 19400
rect 13630 19360 13636 19372
rect 13591 19332 13636 19360
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 14274 19360 14280 19372
rect 14235 19332 14280 19360
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 14734 19320 14740 19372
rect 14792 19360 14798 19372
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14792 19332 14933 19360
rect 14792 19320 14798 19332
rect 14921 19329 14933 19332
rect 14967 19329 14979 19363
rect 15838 19360 15844 19372
rect 15799 19332 15844 19360
rect 14921 19323 14979 19329
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 15930 19320 15936 19372
rect 15988 19360 15994 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 15988 19332 16129 19360
rect 15988 19320 15994 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16298 19360 16304 19372
rect 16259 19332 16304 19360
rect 16117 19323 16175 19329
rect 16298 19320 16304 19332
rect 16356 19320 16362 19372
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 17034 19360 17040 19372
rect 16995 19332 17040 19360
rect 16853 19323 16911 19329
rect 13228 19264 13400 19292
rect 13464 19264 13860 19292
rect 13228 19252 13234 19264
rect 8849 19227 8907 19233
rect 8849 19193 8861 19227
rect 8895 19224 8907 19227
rect 9674 19224 9680 19236
rect 8895 19196 9680 19224
rect 8895 19193 8907 19196
rect 8849 19187 8907 19193
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 9766 19184 9772 19236
rect 9824 19224 9830 19236
rect 13464 19224 13492 19264
rect 9824 19196 13492 19224
rect 13541 19227 13599 19233
rect 9824 19184 9830 19196
rect 13541 19193 13553 19227
rect 13587 19224 13599 19227
rect 13722 19224 13728 19236
rect 13587 19196 13728 19224
rect 13587 19193 13599 19196
rect 13541 19187 13599 19193
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 13832 19224 13860 19264
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13964 19264 14105 19292
rect 13964 19252 13970 19264
rect 14093 19261 14105 19264
rect 14139 19292 14151 19295
rect 15013 19295 15071 19301
rect 15013 19292 15025 19295
rect 14139 19264 15025 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 15013 19261 15025 19264
rect 15059 19292 15071 19295
rect 15194 19292 15200 19304
rect 15059 19264 15200 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15470 19252 15476 19304
rect 15528 19292 15534 19304
rect 16758 19292 16764 19304
rect 15528 19264 16764 19292
rect 15528 19252 15534 19264
rect 16758 19252 16764 19264
rect 16816 19292 16822 19304
rect 16868 19292 16896 19323
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 17218 19320 17224 19372
rect 17276 19360 17282 19372
rect 17494 19360 17500 19372
rect 17276 19332 17500 19360
rect 17276 19320 17282 19332
rect 17494 19320 17500 19332
rect 17552 19360 17558 19372
rect 17696 19369 17724 19400
rect 18414 19388 18420 19400
rect 18472 19428 18478 19440
rect 18994 19431 19052 19437
rect 18994 19428 19006 19431
rect 18472 19400 19006 19428
rect 18472 19388 18478 19400
rect 18994 19397 19006 19400
rect 19040 19428 19052 19431
rect 19536 19428 19564 19468
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 20622 19496 20628 19508
rect 19910 19468 20628 19496
rect 19910 19428 19938 19468
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 20864 19468 21220 19496
rect 20864 19456 20870 19468
rect 19040 19400 19564 19428
rect 19628 19400 19938 19428
rect 19040 19397 19052 19400
rect 18994 19391 19052 19397
rect 17589 19363 17647 19369
rect 17589 19360 17601 19363
rect 17552 19332 17601 19360
rect 17552 19320 17558 19332
rect 17589 19329 17601 19332
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19329 17739 19363
rect 17681 19323 17739 19329
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19360 17923 19363
rect 17954 19360 17960 19372
rect 17911 19332 17960 19360
rect 17911 19329 17923 19332
rect 17865 19323 17923 19329
rect 17954 19320 17960 19332
rect 18012 19360 18018 19372
rect 18322 19360 18328 19372
rect 18012 19332 18328 19360
rect 18012 19320 18018 19332
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18782 19360 18788 19372
rect 18432 19332 18644 19360
rect 18743 19332 18788 19360
rect 16816 19264 16896 19292
rect 16945 19295 17003 19301
rect 16816 19252 16822 19264
rect 16945 19261 16957 19295
rect 16991 19292 17003 19295
rect 16991 19264 17572 19292
rect 16991 19261 17003 19264
rect 16945 19255 17003 19261
rect 15286 19224 15292 19236
rect 13832 19196 15194 19224
rect 15247 19196 15292 19224
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 6638 19156 6644 19168
rect 6052 19128 6644 19156
rect 6052 19116 6058 19128
rect 6638 19116 6644 19128
rect 6696 19116 6702 19168
rect 7650 19156 7656 19168
rect 7611 19128 7656 19156
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 9214 19156 9220 19168
rect 8343 19128 9220 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 9401 19159 9459 19165
rect 9401 19125 9413 19159
rect 9447 19156 9459 19159
rect 9858 19156 9864 19168
rect 9447 19128 9864 19156
rect 9447 19125 9459 19128
rect 9401 19119 9459 19125
rect 9858 19116 9864 19128
rect 9916 19156 9922 19168
rect 10505 19159 10563 19165
rect 10505 19156 10517 19159
rect 9916 19128 10517 19156
rect 9916 19116 9922 19128
rect 10505 19125 10517 19128
rect 10551 19156 10563 19159
rect 10778 19156 10784 19168
rect 10551 19128 10784 19156
rect 10551 19125 10563 19128
rect 10505 19119 10563 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11514 19116 11520 19168
rect 11572 19156 11578 19168
rect 13262 19156 13268 19168
rect 11572 19128 13268 19156
rect 11572 19116 11578 19128
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 13412 19128 13461 19156
rect 13412 19116 13418 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 14918 19156 14924 19168
rect 14879 19128 14924 19156
rect 13449 19119 13507 19125
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 15166 19156 15194 19196
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 15378 19184 15384 19236
rect 15436 19224 15442 19236
rect 16850 19224 16856 19236
rect 15436 19196 16856 19224
rect 15436 19184 15442 19196
rect 16850 19184 16856 19196
rect 16908 19184 16914 19236
rect 17544 19224 17572 19264
rect 17770 19252 17776 19304
rect 17828 19292 17834 19304
rect 18432 19292 18460 19332
rect 18616 19304 18644 19332
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 19628 19360 19656 19400
rect 19978 19388 19984 19440
rect 20036 19428 20042 19440
rect 21192 19428 21220 19468
rect 21266 19456 21272 19508
rect 21324 19496 21330 19508
rect 21361 19499 21419 19505
rect 21361 19496 21373 19499
rect 21324 19468 21373 19496
rect 21324 19456 21330 19468
rect 21361 19465 21373 19468
rect 21407 19496 21419 19499
rect 22646 19496 22652 19508
rect 21407 19468 22652 19496
rect 21407 19465 21419 19468
rect 21361 19459 21419 19465
rect 22646 19456 22652 19468
rect 22704 19496 22710 19508
rect 23198 19496 23204 19508
rect 22704 19468 23204 19496
rect 22704 19456 22710 19468
rect 23198 19456 23204 19468
rect 23256 19456 23262 19508
rect 23382 19456 23388 19508
rect 23440 19496 23446 19508
rect 25406 19496 25412 19508
rect 23440 19468 25412 19496
rect 23440 19456 23446 19468
rect 25406 19456 25412 19468
rect 25464 19456 25470 19508
rect 25590 19456 25596 19508
rect 25648 19496 25654 19508
rect 26602 19496 26608 19508
rect 25648 19468 26608 19496
rect 25648 19456 25654 19468
rect 26602 19456 26608 19468
rect 26660 19456 26666 19508
rect 26694 19456 26700 19508
rect 26752 19496 26758 19508
rect 27430 19496 27436 19508
rect 26752 19468 27436 19496
rect 26752 19456 26758 19468
rect 27430 19456 27436 19468
rect 27488 19456 27494 19508
rect 27522 19456 27528 19508
rect 27580 19496 27586 19508
rect 27798 19496 27804 19508
rect 27580 19468 27804 19496
rect 27580 19456 27586 19468
rect 27798 19456 27804 19468
rect 27856 19496 27862 19508
rect 28442 19496 28448 19508
rect 27856 19468 28448 19496
rect 27856 19456 27862 19468
rect 28442 19456 28448 19468
rect 28500 19456 28506 19508
rect 28626 19496 28632 19508
rect 28552 19468 28632 19496
rect 22186 19428 22192 19440
rect 20036 19400 20378 19428
rect 21192 19400 22192 19428
rect 20036 19388 20042 19400
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 23842 19428 23848 19440
rect 23782 19400 23848 19428
rect 23842 19388 23848 19400
rect 23900 19388 23906 19440
rect 25682 19388 25688 19440
rect 25740 19388 25746 19440
rect 26326 19388 26332 19440
rect 26384 19428 26390 19440
rect 28261 19431 28319 19437
rect 26384 19400 28212 19428
rect 26384 19388 26390 19400
rect 28184 19372 28212 19400
rect 28261 19397 28273 19431
rect 28307 19428 28319 19431
rect 28552 19428 28580 19468
rect 28626 19456 28632 19468
rect 28684 19456 28690 19508
rect 32306 19496 32312 19508
rect 29840 19468 32312 19496
rect 29840 19428 29868 19468
rect 32306 19456 32312 19468
rect 32364 19456 32370 19508
rect 28307 19400 28580 19428
rect 28644 19400 29868 19428
rect 28307 19397 28319 19400
rect 28261 19391 28319 19397
rect 19168 19332 19656 19360
rect 19168 19304 19196 19332
rect 22094 19320 22100 19372
rect 22152 19360 22158 19372
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 22152 19332 22293 19360
rect 22152 19320 22158 19332
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 22281 19323 22339 19329
rect 26605 19363 26663 19369
rect 26605 19329 26617 19363
rect 26651 19360 26663 19363
rect 26970 19360 26976 19372
rect 26651 19332 26976 19360
rect 26651 19329 26663 19332
rect 26605 19323 26663 19329
rect 26970 19320 26976 19332
rect 27028 19320 27034 19372
rect 27246 19320 27252 19372
rect 27304 19360 27310 19372
rect 27341 19363 27399 19369
rect 27341 19360 27353 19363
rect 27304 19332 27353 19360
rect 27304 19320 27310 19332
rect 27341 19329 27353 19332
rect 27387 19329 27399 19363
rect 27341 19323 27399 19329
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 27617 19363 27675 19369
rect 27617 19360 27629 19363
rect 27488 19332 27629 19360
rect 27488 19320 27494 19332
rect 27617 19329 27629 19332
rect 27663 19329 27675 19363
rect 27798 19360 27804 19372
rect 27759 19332 27804 19360
rect 27617 19323 27675 19329
rect 27798 19320 27804 19332
rect 27856 19320 27862 19372
rect 28166 19320 28172 19372
rect 28224 19320 28230 19372
rect 28644 19360 28672 19400
rect 29914 19388 29920 19440
rect 29972 19388 29978 19440
rect 30282 19388 30288 19440
rect 30340 19428 30346 19440
rect 32214 19428 32220 19440
rect 30340 19400 32220 19428
rect 30340 19388 30346 19400
rect 28369 19334 28672 19360
rect 28276 19332 28672 19334
rect 28721 19363 28779 19369
rect 28276 19306 28397 19332
rect 28721 19329 28733 19363
rect 28767 19360 28779 19363
rect 28994 19360 29000 19372
rect 28767 19332 29000 19360
rect 28767 19329 28779 19332
rect 28721 19323 28779 19329
rect 28994 19320 29000 19332
rect 29052 19360 29058 19372
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 29052 19332 29745 19360
rect 29052 19320 29058 19332
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29932 19360 29960 19388
rect 30377 19363 30435 19369
rect 30377 19360 30389 19363
rect 29932 19332 30389 19360
rect 29733 19323 29791 19329
rect 30377 19329 30389 19332
rect 30423 19329 30435 19363
rect 30377 19323 30435 19329
rect 30466 19320 30472 19372
rect 30524 19360 30530 19372
rect 30668 19369 30696 19400
rect 32214 19388 32220 19400
rect 32272 19388 32278 19440
rect 30653 19363 30711 19369
rect 30524 19332 30569 19360
rect 30524 19320 30530 19332
rect 30653 19329 30665 19363
rect 30699 19329 30711 19363
rect 30653 19323 30711 19329
rect 30745 19363 30803 19369
rect 30745 19329 30757 19363
rect 30791 19329 30803 19363
rect 30745 19323 30803 19329
rect 17828 19264 18460 19292
rect 18509 19295 18567 19301
rect 17828 19252 17834 19264
rect 18509 19261 18521 19295
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 18322 19224 18328 19236
rect 17544 19196 18328 19224
rect 18322 19184 18328 19196
rect 18380 19184 18386 19236
rect 18138 19156 18144 19168
rect 15166 19128 18144 19156
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 18414 19116 18420 19168
rect 18472 19156 18478 19168
rect 18527 19156 18555 19255
rect 18598 19252 18604 19304
rect 18656 19292 18662 19304
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18656 19264 18889 19292
rect 18656 19252 18662 19264
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 19150 19252 19156 19304
rect 19208 19252 19214 19304
rect 19892 19301 19898 19304
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19261 19671 19295
rect 19889 19292 19898 19301
rect 19853 19264 19898 19292
rect 19613 19255 19671 19261
rect 19889 19255 19898 19264
rect 19058 19184 19064 19236
rect 19116 19224 19122 19236
rect 19628 19224 19656 19255
rect 19892 19252 19898 19255
rect 19950 19252 19956 19304
rect 20346 19252 20352 19304
rect 20404 19292 20410 19304
rect 21450 19292 21456 19304
rect 20404 19264 21456 19292
rect 20404 19252 20410 19264
rect 21450 19252 21456 19264
rect 21508 19252 21514 19304
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 22066 19264 22569 19292
rect 19116 19196 19656 19224
rect 19116 19184 19122 19196
rect 21174 19184 21180 19236
rect 21232 19224 21238 19236
rect 22066 19224 22094 19264
rect 22557 19261 22569 19264
rect 22603 19261 22615 19295
rect 27525 19295 27583 19301
rect 27525 19292 27537 19295
rect 22557 19255 22615 19261
rect 23584 19264 27537 19292
rect 21232 19196 22094 19224
rect 21232 19184 21238 19196
rect 21266 19156 21272 19168
rect 18472 19128 21272 19156
rect 18472 19116 18478 19128
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 23584 19156 23612 19264
rect 27525 19261 27537 19264
rect 27571 19261 27583 19295
rect 27525 19255 27583 19261
rect 27890 19252 27896 19304
rect 27948 19292 27954 19304
rect 28276 19292 28304 19306
rect 27948 19264 28304 19292
rect 28629 19295 28687 19301
rect 27948 19252 27954 19264
rect 28629 19261 28641 19295
rect 28675 19292 28687 19295
rect 29178 19292 29184 19304
rect 28675 19264 29184 19292
rect 28675 19261 28687 19264
rect 28629 19255 28687 19261
rect 29178 19252 29184 19264
rect 29236 19252 29242 19304
rect 29365 19295 29423 19301
rect 29365 19261 29377 19295
rect 29411 19292 29423 19295
rect 29454 19292 29460 19304
rect 29411 19264 29460 19292
rect 29411 19261 29423 19264
rect 29365 19255 29423 19261
rect 29454 19252 29460 19264
rect 29512 19252 29518 19304
rect 29825 19295 29883 19301
rect 29825 19261 29837 19295
rect 29871 19292 29883 19295
rect 29914 19292 29920 19304
rect 29871 19264 29920 19292
rect 29871 19261 29883 19264
rect 29825 19255 29883 19261
rect 29914 19252 29920 19264
rect 29972 19252 29978 19304
rect 30282 19252 30288 19304
rect 30340 19292 30346 19304
rect 30760 19292 30788 19323
rect 30340 19264 30788 19292
rect 30340 19252 30346 19264
rect 24854 19224 24860 19236
rect 24815 19196 24860 19224
rect 24854 19184 24860 19196
rect 24912 19184 24918 19236
rect 26694 19184 26700 19236
rect 26752 19224 26758 19236
rect 27157 19227 27215 19233
rect 27157 19224 27169 19227
rect 26752 19196 27169 19224
rect 26752 19184 26758 19196
rect 27157 19193 27169 19196
rect 27203 19193 27215 19227
rect 27157 19187 27215 19193
rect 27246 19184 27252 19236
rect 27304 19224 27310 19236
rect 27433 19227 27491 19233
rect 27433 19224 27445 19227
rect 27304 19196 27445 19224
rect 27304 19184 27310 19196
rect 27433 19193 27445 19196
rect 27479 19193 27491 19227
rect 27433 19187 27491 19193
rect 27614 19184 27620 19236
rect 27672 19224 27678 19236
rect 28166 19224 28172 19236
rect 27672 19196 28172 19224
rect 27672 19184 27678 19196
rect 28166 19184 28172 19196
rect 28224 19184 28230 19236
rect 30742 19224 30748 19236
rect 28276 19196 30748 19224
rect 24026 19156 24032 19168
rect 21784 19128 23612 19156
rect 23987 19128 24032 19156
rect 21784 19116 21790 19128
rect 24026 19116 24032 19128
rect 24084 19116 24090 19168
rect 24210 19116 24216 19168
rect 24268 19156 24274 19168
rect 26234 19156 26240 19168
rect 24268 19128 26240 19156
rect 24268 19116 24274 19128
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 26347 19159 26405 19165
rect 26347 19125 26359 19159
rect 26393 19156 26405 19159
rect 28276 19156 28304 19196
rect 30742 19184 30748 19196
rect 30800 19184 30806 19236
rect 26393 19128 28304 19156
rect 26393 19125 26405 19128
rect 26347 19119 26405 19125
rect 28350 19116 28356 19168
rect 28408 19156 28414 19168
rect 28905 19159 28963 19165
rect 28408 19128 28453 19156
rect 28408 19116 28414 19128
rect 28905 19125 28917 19159
rect 28951 19156 28963 19159
rect 29178 19156 29184 19168
rect 28951 19128 29184 19156
rect 28951 19125 28963 19128
rect 28905 19119 28963 19125
rect 29178 19116 29184 19128
rect 29236 19156 29242 19168
rect 30650 19156 30656 19168
rect 29236 19128 30656 19156
rect 29236 19116 29242 19128
rect 30650 19116 30656 19128
rect 30708 19116 30714 19168
rect 30926 19156 30932 19168
rect 30887 19128 30932 19156
rect 30926 19116 30932 19128
rect 30984 19116 30990 19168
rect 1104 19066 31832 19088
rect 1104 19014 4791 19066
rect 4843 19014 4855 19066
rect 4907 19014 4919 19066
rect 4971 19014 4983 19066
rect 5035 19014 5047 19066
rect 5099 19014 12473 19066
rect 12525 19014 12537 19066
rect 12589 19014 12601 19066
rect 12653 19014 12665 19066
rect 12717 19014 12729 19066
rect 12781 19014 20155 19066
rect 20207 19014 20219 19066
rect 20271 19014 20283 19066
rect 20335 19014 20347 19066
rect 20399 19014 20411 19066
rect 20463 19014 27837 19066
rect 27889 19014 27901 19066
rect 27953 19014 27965 19066
rect 28017 19014 28029 19066
rect 28081 19014 28093 19066
rect 28145 19014 31832 19066
rect 1104 18992 31832 19014
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 13722 18952 13728 18964
rect 12308 18924 13728 18952
rect 12308 18912 12314 18924
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 14274 18912 14280 18964
rect 14332 18952 14338 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 14332 18924 14749 18952
rect 14332 18912 14338 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 14737 18915 14795 18921
rect 15010 18912 15016 18964
rect 15068 18952 15074 18964
rect 15470 18952 15476 18964
rect 15068 18924 15476 18952
rect 15068 18912 15074 18924
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 15988 18924 16681 18952
rect 15988 18912 15994 18924
rect 16669 18921 16681 18924
rect 16715 18921 16727 18955
rect 16669 18915 16727 18921
rect 16779 18924 17356 18952
rect 10505 18887 10563 18893
rect 10505 18853 10517 18887
rect 10551 18884 10563 18887
rect 12618 18884 12624 18896
rect 10551 18856 12624 18884
rect 10551 18853 10563 18856
rect 10505 18847 10563 18853
rect 12618 18844 12624 18856
rect 12676 18844 12682 18896
rect 13446 18884 13452 18896
rect 13407 18856 13452 18884
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 13538 18844 13544 18896
rect 13596 18884 13602 18896
rect 16779 18884 16807 18924
rect 13596 18856 16807 18884
rect 16853 18887 16911 18893
rect 13596 18844 13602 18856
rect 16853 18853 16865 18887
rect 16899 18884 16911 18887
rect 17126 18884 17132 18896
rect 16899 18856 17132 18884
rect 16899 18853 16911 18856
rect 16853 18847 16911 18853
rect 17126 18844 17132 18856
rect 17184 18844 17190 18896
rect 9950 18816 9956 18828
rect 9863 18788 9956 18816
rect 9950 18776 9956 18788
rect 10008 18816 10014 18828
rect 10962 18816 10968 18828
rect 10008 18788 10968 18816
rect 10008 18776 10014 18788
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11112 18788 13216 18816
rect 11112 18776 11118 18788
rect 1578 18748 1584 18760
rect 1539 18720 1584 18748
rect 1578 18708 1584 18720
rect 1636 18708 1642 18760
rect 11330 18748 11336 18760
rect 10888 18720 11336 18748
rect 7469 18683 7527 18689
rect 7469 18649 7481 18683
rect 7515 18680 7527 18683
rect 10042 18680 10048 18692
rect 7515 18652 10048 18680
rect 7515 18649 7527 18652
rect 7469 18643 7527 18649
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 7926 18612 7932 18624
rect 7887 18584 7932 18612
rect 7926 18572 7932 18584
rect 7984 18612 7990 18624
rect 8481 18615 8539 18621
rect 8481 18612 8493 18615
rect 7984 18584 8493 18612
rect 7984 18572 7990 18584
rect 8481 18581 8493 18584
rect 8527 18581 8539 18615
rect 8481 18575 8539 18581
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 9272 18584 9321 18612
rect 9272 18572 9278 18584
rect 9309 18581 9321 18584
rect 9355 18612 9367 18615
rect 10888 18612 10916 18720
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 11514 18748 11520 18760
rect 11475 18720 11520 18748
rect 11514 18708 11520 18720
rect 11572 18708 11578 18760
rect 12158 18748 12164 18760
rect 12119 18720 12164 18748
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 12345 18751 12403 18757
rect 12345 18748 12357 18751
rect 12308 18720 12357 18748
rect 12308 18708 12314 18720
rect 12345 18717 12357 18720
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 12805 18751 12863 18757
rect 12805 18717 12817 18751
rect 12851 18748 12863 18751
rect 12986 18748 12992 18760
rect 12851 18720 12992 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 13188 18748 13216 18788
rect 13262 18776 13268 18828
rect 13320 18816 13326 18828
rect 13320 18788 13676 18816
rect 13320 18776 13326 18788
rect 13648 18757 13676 18788
rect 13998 18776 14004 18828
rect 14056 18816 14062 18828
rect 15654 18816 15660 18828
rect 14056 18788 15660 18816
rect 14056 18776 14062 18788
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 15933 18819 15991 18825
rect 15933 18785 15945 18819
rect 15979 18816 15991 18819
rect 17328 18816 17356 18924
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17770 18952 17776 18964
rect 17552 18924 17776 18952
rect 17552 18912 17558 18924
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 17865 18955 17923 18961
rect 17865 18921 17877 18955
rect 17911 18952 17923 18955
rect 19334 18952 19340 18964
rect 17911 18924 19340 18952
rect 17911 18921 17923 18924
rect 17865 18915 17923 18921
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 19521 18955 19579 18961
rect 19521 18921 19533 18955
rect 19567 18952 19579 18955
rect 19610 18952 19616 18964
rect 19567 18924 19616 18952
rect 19567 18921 19579 18924
rect 19521 18915 19579 18921
rect 19610 18912 19616 18924
rect 19668 18952 19674 18964
rect 19978 18952 19984 18964
rect 19668 18924 19984 18952
rect 19668 18912 19674 18924
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20898 18952 20904 18964
rect 20088 18924 20904 18952
rect 17405 18887 17463 18893
rect 17405 18853 17417 18887
rect 17451 18884 17463 18887
rect 18138 18884 18144 18896
rect 17451 18856 18144 18884
rect 17451 18853 17463 18856
rect 17405 18847 17463 18853
rect 18138 18844 18144 18856
rect 18196 18844 18202 18896
rect 18322 18844 18328 18896
rect 18380 18884 18386 18896
rect 18877 18887 18935 18893
rect 18380 18856 18555 18884
rect 18380 18844 18386 18856
rect 17862 18816 17868 18828
rect 15979 18788 17264 18816
rect 15979 18785 15991 18788
rect 15933 18779 15991 18785
rect 13633 18751 13691 18757
rect 13188 18720 13584 18748
rect 11146 18640 11152 18692
rect 11204 18680 11210 18692
rect 13449 18683 13507 18689
rect 13449 18680 13461 18683
rect 11204 18652 13461 18680
rect 11204 18640 11210 18652
rect 13449 18649 13461 18652
rect 13495 18649 13507 18683
rect 13556 18680 13584 18720
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 13722 18708 13728 18760
rect 13780 18748 13786 18760
rect 16114 18748 16120 18760
rect 13780 18720 13825 18748
rect 14752 18720 16120 18748
rect 13780 18708 13786 18720
rect 14752 18680 14780 18720
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 16485 18751 16543 18757
rect 16485 18748 16497 18751
rect 16264 18720 16497 18748
rect 16264 18708 16270 18720
rect 16485 18717 16497 18720
rect 16531 18717 16543 18751
rect 16485 18711 16543 18717
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18748 16819 18751
rect 16850 18748 16856 18760
rect 16807 18720 16856 18748
rect 16807 18717 16819 18720
rect 16761 18711 16819 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 14918 18680 14924 18692
rect 13556 18652 14780 18680
rect 14879 18652 14924 18680
rect 13449 18643 13507 18649
rect 14918 18640 14924 18652
rect 14976 18640 14982 18692
rect 15102 18680 15108 18692
rect 15063 18652 15108 18680
rect 15102 18640 15108 18652
rect 15160 18640 15166 18692
rect 15562 18680 15568 18692
rect 15523 18652 15568 18680
rect 15562 18640 15568 18652
rect 15620 18640 15626 18692
rect 15749 18683 15807 18689
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 16022 18680 16028 18692
rect 15795 18652 16028 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 16393 18683 16451 18689
rect 16393 18649 16405 18683
rect 16439 18680 16451 18683
rect 17126 18680 17132 18692
rect 16439 18652 17132 18680
rect 16439 18649 16451 18652
rect 16393 18643 16451 18649
rect 9355 18584 10916 18612
rect 9355 18581 9367 18584
rect 9309 18575 9367 18581
rect 10962 18572 10968 18624
rect 11020 18612 11026 18624
rect 11422 18612 11428 18624
rect 11020 18584 11428 18612
rect 11020 18572 11026 18584
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 11609 18615 11667 18621
rect 11609 18581 11621 18615
rect 11655 18612 11667 18615
rect 12066 18612 12072 18624
rect 11655 18584 12072 18612
rect 11655 18581 11667 18584
rect 11609 18575 11667 18581
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12345 18615 12403 18621
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 12802 18612 12808 18624
rect 12391 18584 12808 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 12897 18615 12955 18621
rect 12897 18581 12909 18615
rect 12943 18612 12955 18615
rect 13538 18612 13544 18624
rect 12943 18584 13544 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 16408 18612 16436 18643
rect 17126 18640 17132 18652
rect 17184 18640 17190 18692
rect 17236 18680 17264 18788
rect 17328 18788 17868 18816
rect 17328 18757 17356 18788
rect 17862 18776 17868 18788
rect 17920 18776 17926 18828
rect 18414 18816 18420 18828
rect 17972 18788 18420 18816
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17529 18751 17587 18757
rect 17529 18748 17541 18751
rect 17460 18720 17541 18748
rect 17460 18708 17466 18720
rect 17529 18717 17541 18720
rect 17575 18717 17587 18751
rect 17678 18748 17684 18760
rect 17639 18720 17684 18748
rect 17529 18711 17587 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 17770 18708 17776 18760
rect 17828 18748 17834 18760
rect 17972 18748 18000 18788
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 18527 18816 18555 18856
rect 18877 18853 18889 18887
rect 18923 18884 18935 18887
rect 20088 18884 20116 18924
rect 20898 18912 20904 18924
rect 20956 18912 20962 18964
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 23845 18955 23903 18961
rect 23845 18952 23857 18955
rect 21876 18924 23857 18952
rect 21876 18912 21882 18924
rect 23845 18921 23857 18924
rect 23891 18921 23903 18955
rect 26326 18952 26332 18964
rect 23845 18915 23903 18921
rect 23952 18924 26332 18952
rect 22462 18884 22468 18896
rect 18923 18856 20116 18884
rect 22423 18856 22468 18884
rect 18923 18853 18935 18856
rect 18877 18847 18935 18853
rect 22462 18844 22468 18856
rect 22520 18844 22526 18896
rect 22738 18844 22744 18896
rect 22796 18884 22802 18896
rect 23661 18887 23719 18893
rect 23661 18884 23673 18887
rect 22796 18856 23673 18884
rect 22796 18844 22802 18856
rect 23661 18853 23673 18856
rect 23707 18853 23719 18887
rect 23661 18847 23719 18853
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 18527 18788 20269 18816
rect 20257 18785 20269 18788
rect 20303 18785 20315 18819
rect 20257 18779 20315 18785
rect 20346 18776 20352 18828
rect 20404 18816 20410 18828
rect 23017 18819 23075 18825
rect 23017 18816 23029 18819
rect 20404 18788 23029 18816
rect 20404 18776 20410 18788
rect 23017 18785 23029 18788
rect 23063 18785 23075 18819
rect 23017 18779 23075 18785
rect 23198 18776 23204 18828
rect 23256 18816 23262 18828
rect 23952 18816 23980 18924
rect 26326 18912 26332 18924
rect 26384 18912 26390 18964
rect 26970 18912 26976 18964
rect 27028 18952 27034 18964
rect 27028 18924 27568 18952
rect 27028 18912 27034 18924
rect 24946 18844 24952 18896
rect 25004 18844 25010 18896
rect 27430 18884 27436 18896
rect 26252 18856 27200 18884
rect 27391 18856 27436 18884
rect 23256 18788 23980 18816
rect 24964 18816 24992 18844
rect 26252 18816 26280 18856
rect 24964 18788 26280 18816
rect 23256 18776 23262 18788
rect 26326 18776 26332 18828
rect 26384 18816 26390 18828
rect 26602 18816 26608 18828
rect 26384 18788 26608 18816
rect 26384 18776 26390 18788
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 26786 18816 26792 18828
rect 26747 18788 26792 18816
rect 26786 18776 26792 18788
rect 26844 18776 26850 18828
rect 27172 18825 27200 18856
rect 27430 18844 27436 18856
rect 27488 18844 27494 18896
rect 27540 18884 27568 18924
rect 27706 18912 27712 18964
rect 27764 18952 27770 18964
rect 27893 18955 27951 18961
rect 27893 18952 27905 18955
rect 27764 18924 27905 18952
rect 27764 18912 27770 18924
rect 27893 18921 27905 18924
rect 27939 18921 27951 18955
rect 28074 18952 28080 18964
rect 27893 18915 27951 18921
rect 28000 18924 28080 18952
rect 28000 18884 28028 18924
rect 28074 18912 28080 18924
rect 28132 18912 28138 18964
rect 28350 18952 28356 18964
rect 28184 18924 28356 18952
rect 27540 18856 28028 18884
rect 27157 18819 27215 18825
rect 27157 18785 27169 18819
rect 27203 18816 27215 18819
rect 27890 18816 27896 18828
rect 27203 18788 27896 18816
rect 27203 18785 27215 18788
rect 27157 18779 27215 18785
rect 27890 18776 27896 18788
rect 27948 18776 27954 18828
rect 27982 18776 27988 18828
rect 28040 18816 28046 18828
rect 28184 18825 28212 18924
rect 28350 18912 28356 18924
rect 28408 18912 28414 18964
rect 28442 18912 28448 18964
rect 28500 18952 28506 18964
rect 29089 18955 29147 18961
rect 29089 18952 29101 18955
rect 28500 18924 29101 18952
rect 28500 18912 28506 18924
rect 29089 18921 29101 18924
rect 29135 18921 29147 18955
rect 29089 18915 29147 18921
rect 29546 18912 29552 18964
rect 29604 18952 29610 18964
rect 31205 18955 31263 18961
rect 31205 18952 31217 18955
rect 29604 18924 31217 18952
rect 29604 18912 29610 18924
rect 31205 18921 31217 18924
rect 31251 18921 31263 18955
rect 31205 18915 31263 18921
rect 29733 18887 29791 18893
rect 28460 18856 29040 18884
rect 28078 18819 28136 18825
rect 28078 18816 28090 18819
rect 28040 18788 28090 18816
rect 28040 18776 28046 18788
rect 28078 18785 28090 18788
rect 28124 18785 28136 18819
rect 28078 18779 28136 18785
rect 28169 18819 28227 18825
rect 28169 18785 28181 18819
rect 28215 18785 28227 18819
rect 28169 18779 28227 18785
rect 28261 18819 28319 18825
rect 28261 18785 28273 18819
rect 28307 18816 28319 18819
rect 28460 18816 28488 18856
rect 28307 18788 28488 18816
rect 28307 18785 28319 18788
rect 28261 18779 28319 18785
rect 28534 18776 28540 18828
rect 28592 18816 28598 18828
rect 28905 18819 28963 18825
rect 28905 18816 28917 18819
rect 28592 18788 28917 18816
rect 28592 18776 28598 18788
rect 28905 18785 28917 18788
rect 28951 18785 28963 18819
rect 29012 18816 29040 18856
rect 29733 18853 29745 18887
rect 29779 18884 29791 18887
rect 31110 18884 31116 18896
rect 29779 18856 31116 18884
rect 29779 18853 29791 18856
rect 29733 18847 29791 18853
rect 31110 18844 31116 18856
rect 31168 18844 31174 18896
rect 30006 18816 30012 18828
rect 29012 18788 30012 18816
rect 28905 18779 28963 18785
rect 30006 18776 30012 18788
rect 30064 18776 30070 18828
rect 30193 18819 30251 18825
rect 30193 18785 30205 18819
rect 30239 18816 30251 18819
rect 30926 18816 30932 18828
rect 30239 18788 30932 18816
rect 30239 18785 30251 18788
rect 30193 18779 30251 18785
rect 30926 18776 30932 18788
rect 30984 18776 30990 18828
rect 17828 18720 18000 18748
rect 17828 18708 17834 18720
rect 18046 18708 18052 18760
rect 18104 18748 18110 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18104 18720 18521 18748
rect 18104 18708 18110 18720
rect 18509 18717 18521 18720
rect 18555 18748 18567 18751
rect 18782 18748 18788 18760
rect 18555 18720 18788 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 18932 18720 19196 18748
rect 18932 18708 18938 18720
rect 19168 18680 19196 18720
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 19981 18751 20039 18757
rect 19981 18748 19993 18751
rect 19668 18720 19993 18748
rect 19668 18708 19674 18720
rect 19981 18717 19993 18720
rect 20027 18717 20039 18751
rect 19981 18711 20039 18717
rect 21634 18708 21640 18760
rect 21692 18748 21698 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 21692 18720 22937 18748
rect 21692 18708 21698 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 24210 18748 24216 18760
rect 22925 18711 22983 18717
rect 23446 18720 24216 18748
rect 20530 18680 20536 18692
rect 17236 18652 19104 18680
rect 19168 18652 20536 18680
rect 13780 18584 16436 18612
rect 13780 18572 13786 18584
rect 16482 18572 16488 18624
rect 16540 18612 16546 18624
rect 18874 18612 18880 18624
rect 16540 18584 18880 18612
rect 16540 18572 16546 18584
rect 18874 18572 18880 18584
rect 18932 18572 18938 18624
rect 19076 18612 19104 18652
rect 20530 18640 20536 18652
rect 20588 18640 20594 18692
rect 21266 18640 21272 18692
rect 21324 18640 21330 18692
rect 22002 18680 22008 18692
rect 21963 18652 22008 18680
rect 22002 18640 22008 18652
rect 22060 18680 22066 18692
rect 22833 18683 22891 18689
rect 22833 18680 22845 18683
rect 22060 18652 22845 18680
rect 22060 18640 22066 18652
rect 22833 18649 22845 18652
rect 22879 18680 22891 18683
rect 23446 18680 23474 18720
rect 24210 18708 24216 18720
rect 24268 18708 24274 18760
rect 24946 18708 24952 18760
rect 25004 18708 25010 18760
rect 27430 18708 27436 18760
rect 27488 18748 27494 18760
rect 28353 18751 28411 18757
rect 28353 18748 28365 18751
rect 27488 18720 28365 18748
rect 27488 18708 27494 18720
rect 28353 18717 28365 18720
rect 28399 18717 28411 18751
rect 28353 18711 28411 18717
rect 29181 18751 29239 18757
rect 29181 18717 29193 18751
rect 29227 18748 29239 18751
rect 30098 18748 30104 18760
rect 29227 18720 29408 18748
rect 30059 18720 30104 18748
rect 29227 18717 29239 18720
rect 29181 18711 29239 18717
rect 23813 18683 23871 18689
rect 23813 18680 23825 18683
rect 22879 18652 23474 18680
rect 23584 18652 23825 18680
rect 22879 18649 22891 18652
rect 22833 18643 22891 18649
rect 21818 18612 21824 18624
rect 19076 18584 21824 18612
rect 21818 18572 21824 18584
rect 21876 18572 21882 18624
rect 22278 18572 22284 18624
rect 22336 18612 22342 18624
rect 23584 18612 23612 18652
rect 23813 18649 23825 18652
rect 23859 18649 23871 18683
rect 23813 18643 23871 18649
rect 24029 18683 24087 18689
rect 24029 18649 24041 18683
rect 24075 18649 24087 18683
rect 24029 18643 24087 18649
rect 26053 18683 26111 18689
rect 26053 18649 26065 18683
rect 26099 18680 26111 18683
rect 26142 18680 26148 18692
rect 26099 18652 26148 18680
rect 26099 18649 26111 18652
rect 26053 18643 26111 18649
rect 22336 18584 23612 18612
rect 22336 18572 22342 18584
rect 23658 18572 23664 18624
rect 23716 18612 23722 18624
rect 24044 18612 24072 18643
rect 26142 18640 26148 18652
rect 26200 18640 26206 18692
rect 26970 18680 26976 18692
rect 26712 18652 26976 18680
rect 23716 18584 24072 18612
rect 24581 18615 24639 18621
rect 23716 18572 23722 18584
rect 24581 18581 24593 18615
rect 24627 18612 24639 18615
rect 25222 18612 25228 18624
rect 24627 18584 25228 18612
rect 24627 18581 24639 18584
rect 24581 18575 24639 18581
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 25958 18572 25964 18624
rect 26016 18612 26022 18624
rect 26712 18612 26740 18652
rect 26970 18640 26976 18652
rect 27028 18640 27034 18692
rect 27274 18683 27332 18689
rect 27274 18649 27286 18683
rect 27320 18649 27332 18683
rect 27274 18643 27332 18649
rect 26016 18584 26740 18612
rect 26016 18572 26022 18584
rect 26786 18572 26792 18624
rect 26844 18612 26850 18624
rect 27065 18615 27123 18621
rect 27065 18612 27077 18615
rect 26844 18584 27077 18612
rect 26844 18572 26850 18584
rect 27065 18581 27077 18584
rect 27111 18581 27123 18615
rect 27289 18612 27317 18643
rect 28074 18640 28080 18692
rect 28132 18680 28138 18692
rect 28905 18683 28963 18689
rect 28905 18680 28917 18683
rect 28132 18652 28917 18680
rect 28132 18640 28138 18652
rect 28905 18649 28917 18652
rect 28951 18649 28963 18683
rect 28905 18643 28963 18649
rect 29380 18624 29408 18720
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 30742 18748 30748 18760
rect 30703 18720 30748 18748
rect 30742 18708 30748 18720
rect 30800 18708 30806 18760
rect 31021 18751 31079 18757
rect 31021 18717 31033 18751
rect 31067 18748 31079 18751
rect 31662 18748 31668 18760
rect 31067 18720 31668 18748
rect 31067 18717 31079 18720
rect 31021 18711 31079 18717
rect 31662 18708 31668 18720
rect 31720 18708 31726 18760
rect 30650 18640 30656 18692
rect 30708 18680 30714 18692
rect 30837 18683 30895 18689
rect 30837 18680 30849 18683
rect 30708 18652 30849 18680
rect 30708 18640 30714 18652
rect 30837 18649 30849 18652
rect 30883 18680 30895 18683
rect 32490 18680 32496 18692
rect 30883 18652 32496 18680
rect 30883 18649 30895 18652
rect 30837 18643 30895 18649
rect 32490 18640 32496 18652
rect 32548 18640 32554 18692
rect 28442 18612 28448 18624
rect 27289 18584 28448 18612
rect 27065 18575 27123 18581
rect 28442 18572 28448 18584
rect 28500 18612 28506 18624
rect 29178 18612 29184 18624
rect 28500 18584 29184 18612
rect 28500 18572 28506 18584
rect 29178 18572 29184 18584
rect 29236 18572 29242 18624
rect 29362 18572 29368 18624
rect 29420 18572 29426 18624
rect 1104 18522 31992 18544
rect 1104 18470 8632 18522
rect 8684 18470 8696 18522
rect 8748 18470 8760 18522
rect 8812 18470 8824 18522
rect 8876 18470 8888 18522
rect 8940 18470 16314 18522
rect 16366 18470 16378 18522
rect 16430 18470 16442 18522
rect 16494 18470 16506 18522
rect 16558 18470 16570 18522
rect 16622 18470 23996 18522
rect 24048 18470 24060 18522
rect 24112 18470 24124 18522
rect 24176 18470 24188 18522
rect 24240 18470 24252 18522
rect 24304 18470 31678 18522
rect 31730 18470 31742 18522
rect 31794 18470 31806 18522
rect 31858 18470 31870 18522
rect 31922 18470 31934 18522
rect 31986 18470 31992 18522
rect 1104 18448 31992 18470
rect 10042 18408 10048 18420
rect 10003 18380 10048 18408
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 12897 18411 12955 18417
rect 12897 18377 12909 18411
rect 12943 18408 12955 18411
rect 15010 18408 15016 18420
rect 12943 18380 15016 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 15010 18368 15016 18380
rect 15068 18368 15074 18420
rect 15181 18411 15239 18417
rect 15181 18377 15193 18411
rect 15227 18408 15239 18411
rect 15470 18408 15476 18420
rect 15227 18380 15476 18408
rect 15227 18377 15239 18380
rect 15181 18371 15239 18377
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 15841 18411 15899 18417
rect 15841 18408 15853 18411
rect 15580 18380 15853 18408
rect 8389 18343 8447 18349
rect 8389 18309 8401 18343
rect 8435 18340 8447 18343
rect 11514 18340 11520 18352
rect 8435 18312 11520 18340
rect 8435 18309 8447 18312
rect 8389 18303 8447 18309
rect 11514 18300 11520 18312
rect 11572 18340 11578 18352
rect 11790 18340 11796 18352
rect 11572 18312 11796 18340
rect 11572 18300 11578 18312
rect 11790 18300 11796 18312
rect 11848 18340 11854 18352
rect 12253 18343 12311 18349
rect 11848 18312 12204 18340
rect 11848 18300 11854 18312
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 11238 18272 11244 18284
rect 9640 18244 11244 18272
rect 9640 18232 9646 18244
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 12176 18281 12204 18312
rect 12253 18309 12265 18343
rect 12299 18340 12311 18343
rect 14090 18340 14096 18352
rect 12299 18312 14096 18340
rect 12299 18309 12311 18312
rect 12253 18303 12311 18309
rect 14090 18300 14096 18312
rect 14148 18300 14154 18352
rect 14185 18343 14243 18349
rect 14185 18309 14197 18343
rect 14231 18340 14243 18343
rect 14274 18340 14280 18352
rect 14231 18312 14280 18340
rect 14231 18309 14243 18312
rect 14185 18303 14243 18309
rect 14274 18300 14280 18312
rect 14332 18300 14338 18352
rect 14458 18340 14464 18352
rect 14430 18315 14464 18340
rect 14415 18309 14464 18315
rect 12161 18275 12219 18281
rect 12161 18241 12173 18275
rect 12207 18241 12219 18275
rect 12802 18272 12808 18284
rect 12763 18244 12808 18272
rect 12161 18235 12219 18241
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 13630 18272 13636 18284
rect 13543 18244 13636 18272
rect 13630 18232 13636 18244
rect 13688 18272 13694 18284
rect 14415 18275 14427 18309
rect 14461 18300 14464 18309
rect 14516 18300 14522 18352
rect 14918 18300 14924 18352
rect 14976 18340 14982 18352
rect 15381 18343 15439 18349
rect 15381 18340 15393 18343
rect 14976 18312 15393 18340
rect 14976 18300 14982 18312
rect 15381 18309 15393 18312
rect 15427 18309 15439 18343
rect 15381 18303 15439 18309
rect 14461 18275 14473 18300
rect 13688 18244 14152 18272
rect 14415 18269 14473 18275
rect 13688 18232 13694 18244
rect 10870 18204 10876 18216
rect 9876 18176 10876 18204
rect 9876 18148 9904 18176
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 13998 18204 14004 18216
rect 12676 18176 14004 18204
rect 12676 18164 12682 18176
rect 13998 18164 14004 18176
rect 14056 18164 14062 18216
rect 6638 18096 6644 18148
rect 6696 18136 6702 18148
rect 8941 18139 8999 18145
rect 8941 18136 8953 18139
rect 6696 18108 8953 18136
rect 6696 18096 6702 18108
rect 8941 18105 8953 18108
rect 8987 18136 8999 18139
rect 9858 18136 9864 18148
rect 8987 18108 9864 18136
rect 8987 18105 8999 18108
rect 8941 18099 8999 18105
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 11054 18096 11060 18148
rect 11112 18136 11118 18148
rect 12250 18136 12256 18148
rect 11112 18108 12256 18136
rect 11112 18096 11118 18108
rect 12250 18096 12256 18108
rect 12308 18136 12314 18148
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 12308 18108 13645 18136
rect 12308 18096 12314 18108
rect 13633 18105 13645 18108
rect 13679 18136 13691 18139
rect 13906 18136 13912 18148
rect 13679 18108 13912 18136
rect 13679 18105 13691 18108
rect 13633 18099 13691 18105
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 14124 18136 14152 18244
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 15580 18272 15608 18380
rect 15841 18377 15853 18380
rect 15887 18377 15899 18411
rect 15841 18371 15899 18377
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 17218 18408 17224 18420
rect 16080 18380 17224 18408
rect 16080 18368 16086 18380
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 17497 18411 17555 18417
rect 17497 18377 17509 18411
rect 17543 18408 17555 18411
rect 17543 18380 17815 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 16301 18343 16359 18349
rect 14608 18244 15608 18272
rect 15665 18312 16151 18340
rect 14608 18232 14614 18244
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 15665 18204 15693 18312
rect 16022 18272 16028 18284
rect 15983 18244 16028 18272
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16123 18272 16151 18312
rect 16301 18309 16313 18343
rect 16347 18340 16359 18343
rect 16574 18340 16580 18352
rect 16347 18312 16580 18340
rect 16347 18309 16359 18312
rect 16301 18303 16359 18309
rect 16574 18300 16580 18312
rect 16632 18300 16638 18352
rect 16850 18300 16856 18352
rect 16908 18340 16914 18352
rect 17310 18340 17316 18352
rect 16908 18312 17316 18340
rect 16908 18300 16914 18312
rect 17310 18300 17316 18312
rect 17368 18300 17374 18352
rect 17512 18272 17540 18371
rect 17678 18340 17684 18352
rect 17639 18312 17684 18340
rect 17678 18300 17684 18312
rect 17736 18300 17742 18352
rect 16123 18244 17540 18272
rect 17589 18275 17647 18281
rect 17589 18241 17601 18275
rect 17635 18241 17647 18275
rect 17787 18272 17815 18380
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 21361 18411 21419 18417
rect 21361 18408 21373 18411
rect 18380 18380 21373 18408
rect 18380 18368 18386 18380
rect 21361 18377 21373 18380
rect 21407 18377 21419 18411
rect 21361 18371 21419 18377
rect 17865 18343 17923 18349
rect 17865 18309 17877 18343
rect 17911 18340 17923 18343
rect 17954 18340 17960 18352
rect 17911 18312 17960 18340
rect 17911 18309 17923 18312
rect 17865 18303 17923 18309
rect 17954 18300 17960 18312
rect 18012 18300 18018 18352
rect 18138 18300 18144 18352
rect 18196 18340 18202 18352
rect 19334 18340 19340 18352
rect 18196 18312 19340 18340
rect 18196 18300 18202 18312
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 19886 18340 19892 18352
rect 19847 18312 19892 18340
rect 19886 18300 19892 18312
rect 19944 18300 19950 18352
rect 19978 18300 19984 18352
rect 20036 18340 20042 18352
rect 21376 18340 21404 18371
rect 21450 18368 21456 18420
rect 21508 18408 21514 18420
rect 25317 18411 25375 18417
rect 25317 18408 25329 18411
rect 21508 18380 25329 18408
rect 21508 18368 21514 18380
rect 25317 18377 25329 18380
rect 25363 18377 25375 18411
rect 25317 18371 25375 18377
rect 25774 18368 25780 18420
rect 25832 18408 25838 18420
rect 26878 18408 26884 18420
rect 25832 18380 26884 18408
rect 25832 18368 25838 18380
rect 26878 18368 26884 18380
rect 26936 18368 26942 18420
rect 27175 18380 27659 18408
rect 21818 18340 21824 18352
rect 20036 18312 20378 18340
rect 21376 18312 21824 18340
rect 20036 18300 20042 18312
rect 21818 18300 21824 18312
rect 21876 18300 21882 18352
rect 22186 18300 22192 18352
rect 22244 18340 22250 18352
rect 22281 18343 22339 18349
rect 22281 18340 22293 18343
rect 22244 18312 22293 18340
rect 22244 18300 22250 18312
rect 22281 18309 22293 18312
rect 22327 18309 22339 18343
rect 22281 18303 22339 18309
rect 22738 18300 22744 18352
rect 22796 18300 22802 18352
rect 23566 18300 23572 18352
rect 23624 18340 23630 18352
rect 25869 18343 25927 18349
rect 23624 18312 25636 18340
rect 23624 18300 23630 18312
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 17787 18244 18613 18272
rect 17589 18235 17647 18241
rect 18601 18241 18613 18244
rect 18647 18272 18659 18275
rect 19150 18272 19156 18284
rect 18647 18244 19156 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 14240 18176 15693 18204
rect 14240 18164 14246 18176
rect 16114 18164 16120 18216
rect 16172 18204 16178 18216
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 16172 18176 16221 18204
rect 16172 18164 16178 18176
rect 16209 18173 16221 18176
rect 16255 18204 16267 18207
rect 16390 18204 16396 18216
rect 16255 18176 16396 18204
rect 16255 18173 16267 18176
rect 16209 18167 16267 18173
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 17604 18204 17632 18235
rect 19150 18232 19156 18244
rect 19208 18232 19214 18284
rect 19610 18272 19616 18284
rect 19571 18244 19616 18272
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 23750 18232 23756 18284
rect 23808 18272 23814 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 23808 18244 24225 18272
rect 23808 18232 23814 18244
rect 24213 18241 24225 18244
rect 24259 18272 24271 18275
rect 24394 18272 24400 18284
rect 24259 18244 24400 18272
rect 24259 18241 24271 18244
rect 24213 18235 24271 18241
rect 24394 18232 24400 18244
rect 24452 18232 24458 18284
rect 24673 18275 24731 18281
rect 24673 18241 24685 18275
rect 24719 18272 24731 18275
rect 25038 18272 25044 18284
rect 24719 18244 25044 18272
rect 24719 18241 24731 18244
rect 24673 18235 24731 18241
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25608 18281 25636 18312
rect 25869 18309 25881 18343
rect 25915 18340 25927 18343
rect 26142 18340 26148 18352
rect 25915 18312 26148 18340
rect 25915 18309 25927 18312
rect 25869 18303 25927 18309
rect 26142 18300 26148 18312
rect 26200 18300 26206 18352
rect 26234 18300 26240 18352
rect 26292 18340 26298 18352
rect 26292 18312 26556 18340
rect 26292 18300 26298 18312
rect 25593 18275 25651 18281
rect 25593 18241 25605 18275
rect 25639 18241 25651 18275
rect 25593 18235 25651 18241
rect 26421 18275 26479 18281
rect 26421 18241 26433 18275
rect 26467 18241 26479 18275
rect 26528 18272 26556 18312
rect 26694 18300 26700 18352
rect 26752 18340 26758 18352
rect 27175 18340 27203 18380
rect 27341 18343 27399 18349
rect 27341 18340 27353 18343
rect 26752 18312 27203 18340
rect 26752 18300 26758 18312
rect 26605 18275 26663 18281
rect 26605 18272 26617 18275
rect 26528 18244 26617 18272
rect 26421 18235 26479 18241
rect 26605 18241 26617 18244
rect 26651 18272 26663 18275
rect 26970 18272 26976 18284
rect 26651 18244 26976 18272
rect 26651 18241 26663 18244
rect 26605 18235 26663 18241
rect 17678 18204 17684 18216
rect 17604 18176 17684 18204
rect 17678 18164 17684 18176
rect 17736 18164 17742 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 17945 18176 18337 18204
rect 14458 18136 14464 18148
rect 14124 18108 14464 18136
rect 14458 18096 14464 18108
rect 14516 18096 14522 18148
rect 14553 18139 14611 18145
rect 14553 18105 14565 18139
rect 14599 18136 14611 18139
rect 17945 18136 17973 18176
rect 18325 18173 18337 18176
rect 18371 18173 18383 18207
rect 21634 18204 21640 18216
rect 18325 18167 18383 18173
rect 19260 18176 21640 18204
rect 14599 18108 17973 18136
rect 14599 18105 14611 18108
rect 14553 18099 14611 18105
rect 18046 18096 18052 18148
rect 18104 18136 18110 18148
rect 19260 18136 19288 18176
rect 21634 18164 21640 18176
rect 21692 18164 21698 18216
rect 22005 18207 22063 18213
rect 22005 18173 22017 18207
rect 22051 18204 22063 18207
rect 22370 18204 22376 18216
rect 22051 18176 22376 18204
rect 22051 18173 22063 18176
rect 22005 18167 22063 18173
rect 18104 18108 19288 18136
rect 18104 18096 18110 18108
rect 21082 18096 21088 18148
rect 21140 18136 21146 18148
rect 22020 18136 22048 18167
rect 22370 18164 22376 18176
rect 22428 18204 22434 18216
rect 23014 18204 23020 18216
rect 22428 18176 23020 18204
rect 22428 18164 22434 18176
rect 23014 18164 23020 18176
rect 23072 18164 23078 18216
rect 24581 18207 24639 18213
rect 24581 18173 24593 18207
rect 24627 18204 24639 18207
rect 25314 18204 25320 18216
rect 24627 18176 25320 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 25501 18207 25559 18213
rect 25501 18173 25513 18207
rect 25547 18204 25559 18207
rect 25774 18204 25780 18216
rect 25547 18176 25780 18204
rect 25547 18173 25559 18176
rect 25501 18167 25559 18173
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 25958 18204 25964 18216
rect 25919 18176 25964 18204
rect 25958 18164 25964 18176
rect 26016 18164 26022 18216
rect 26436 18204 26464 18235
rect 26970 18232 26976 18244
rect 27028 18232 27034 18284
rect 27175 18281 27203 18312
rect 27264 18312 27353 18340
rect 27157 18275 27215 18281
rect 27157 18241 27169 18275
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 26064 18176 26464 18204
rect 27264 18204 27292 18312
rect 27341 18309 27353 18312
rect 27387 18309 27399 18343
rect 27341 18303 27399 18309
rect 27430 18272 27436 18284
rect 27391 18244 27436 18272
rect 27430 18232 27436 18244
rect 27488 18232 27494 18284
rect 27525 18275 27583 18281
rect 27525 18241 27537 18275
rect 27571 18241 27583 18275
rect 27631 18272 27659 18380
rect 27706 18368 27712 18420
rect 27764 18408 27770 18420
rect 30190 18408 30196 18420
rect 27764 18380 30196 18408
rect 27764 18368 27770 18380
rect 30190 18368 30196 18380
rect 30248 18368 30254 18420
rect 30834 18368 30840 18420
rect 30892 18408 30898 18420
rect 31113 18411 31171 18417
rect 31113 18408 31125 18411
rect 30892 18380 31125 18408
rect 30892 18368 30898 18380
rect 31113 18377 31125 18380
rect 31159 18377 31171 18411
rect 31113 18371 31171 18377
rect 27890 18300 27896 18352
rect 27948 18340 27954 18352
rect 29181 18343 29239 18349
rect 27948 18312 28932 18340
rect 27948 18300 27954 18312
rect 27982 18272 27988 18284
rect 27631 18244 27988 18272
rect 27525 18235 27583 18241
rect 27540 18204 27568 18235
rect 27982 18232 27988 18244
rect 28040 18272 28046 18284
rect 28258 18272 28264 18284
rect 28040 18244 28264 18272
rect 28040 18232 28046 18244
rect 28258 18232 28264 18244
rect 28316 18232 28322 18284
rect 28442 18232 28448 18284
rect 28500 18272 28506 18284
rect 28537 18275 28595 18281
rect 28537 18272 28549 18275
rect 28500 18244 28549 18272
rect 28500 18232 28506 18244
rect 28537 18241 28549 18244
rect 28583 18241 28595 18275
rect 28537 18235 28595 18241
rect 28074 18204 28080 18216
rect 27264 18176 27476 18204
rect 27540 18176 28080 18204
rect 21140 18108 22048 18136
rect 21140 18096 21146 18108
rect 23474 18096 23480 18148
rect 23532 18136 23538 18148
rect 26064 18136 26092 18176
rect 23532 18108 26092 18136
rect 26421 18139 26479 18145
rect 23532 18096 23538 18108
rect 26421 18105 26433 18139
rect 26467 18136 26479 18139
rect 26510 18136 26516 18148
rect 26467 18108 26516 18136
rect 26467 18105 26479 18108
rect 26421 18099 26479 18105
rect 26510 18096 26516 18108
rect 26568 18096 26574 18148
rect 27448 18136 27476 18176
rect 28074 18164 28080 18176
rect 28132 18164 28138 18216
rect 28166 18164 28172 18216
rect 28224 18204 28230 18216
rect 28629 18207 28687 18213
rect 28224 18176 28269 18204
rect 28224 18164 28230 18176
rect 28629 18173 28641 18207
rect 28675 18204 28687 18207
rect 28810 18204 28816 18216
rect 28675 18176 28816 18204
rect 28675 18173 28687 18176
rect 28629 18167 28687 18173
rect 28810 18164 28816 18176
rect 28868 18164 28874 18216
rect 28904 18204 28932 18312
rect 29181 18309 29193 18343
rect 29227 18340 29239 18343
rect 32766 18340 32772 18352
rect 29227 18312 32772 18340
rect 29227 18309 29239 18312
rect 29181 18303 29239 18309
rect 32766 18300 32772 18312
rect 32824 18300 32830 18352
rect 28994 18232 29000 18284
rect 29052 18272 29058 18284
rect 29365 18275 29423 18281
rect 29365 18272 29377 18275
rect 29052 18244 29377 18272
rect 29052 18232 29058 18244
rect 29365 18241 29377 18244
rect 29411 18241 29423 18275
rect 29365 18235 29423 18241
rect 29178 18204 29184 18216
rect 28904 18176 29184 18204
rect 29178 18164 29184 18176
rect 29236 18164 29242 18216
rect 29380 18204 29408 18235
rect 29454 18232 29460 18284
rect 29512 18272 29518 18284
rect 29638 18272 29644 18284
rect 29512 18244 29557 18272
rect 29599 18244 29644 18272
rect 29512 18232 29518 18244
rect 29638 18232 29644 18244
rect 29696 18232 29702 18284
rect 29733 18275 29791 18281
rect 29733 18241 29745 18275
rect 29779 18272 29791 18275
rect 30006 18272 30012 18284
rect 29779 18244 30012 18272
rect 29779 18241 29791 18244
rect 29733 18235 29791 18241
rect 30006 18232 30012 18244
rect 30064 18232 30070 18284
rect 30190 18272 30196 18284
rect 30151 18244 30196 18272
rect 30190 18232 30196 18244
rect 30248 18232 30254 18284
rect 30466 18232 30472 18284
rect 30524 18272 30530 18284
rect 31113 18275 31171 18281
rect 31113 18272 31125 18275
rect 30524 18244 31125 18272
rect 30524 18232 30530 18244
rect 31113 18241 31125 18244
rect 31159 18241 31171 18275
rect 31113 18235 31171 18241
rect 31297 18275 31355 18281
rect 31297 18241 31309 18275
rect 31343 18272 31355 18275
rect 31662 18272 31668 18284
rect 31343 18244 31668 18272
rect 31343 18241 31355 18244
rect 31297 18235 31355 18241
rect 31662 18232 31668 18244
rect 31720 18232 31726 18284
rect 30282 18204 30288 18216
rect 29380 18176 30288 18204
rect 30282 18164 30288 18176
rect 30340 18164 30346 18216
rect 30377 18207 30435 18213
rect 30377 18173 30389 18207
rect 30423 18204 30435 18207
rect 32398 18204 32404 18216
rect 30423 18176 32404 18204
rect 30423 18173 30435 18176
rect 30377 18167 30435 18173
rect 32398 18164 32404 18176
rect 32456 18164 32462 18216
rect 27798 18136 27804 18148
rect 27448 18108 27804 18136
rect 27798 18096 27804 18108
rect 27856 18096 27862 18148
rect 29822 18136 29828 18148
rect 28460 18108 29828 18136
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 9490 18068 9496 18080
rect 9451 18040 9496 18068
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 10597 18071 10655 18077
rect 10597 18037 10609 18071
rect 10643 18068 10655 18071
rect 10870 18068 10876 18080
rect 10643 18040 10876 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11149 18071 11207 18077
rect 11149 18037 11161 18071
rect 11195 18068 11207 18071
rect 11238 18068 11244 18080
rect 11195 18040 11244 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11238 18028 11244 18040
rect 11296 18068 11302 18080
rect 12158 18068 12164 18080
rect 11296 18040 12164 18068
rect 11296 18028 11302 18040
rect 12158 18028 12164 18040
rect 12216 18068 12222 18080
rect 13722 18068 13728 18080
rect 12216 18040 13728 18068
rect 12216 18028 12222 18040
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14369 18071 14427 18077
rect 14369 18068 14381 18071
rect 13872 18040 14381 18068
rect 13872 18028 13878 18040
rect 14369 18037 14381 18040
rect 14415 18068 14427 18071
rect 14826 18068 14832 18080
rect 14415 18040 14832 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 15010 18068 15016 18080
rect 14971 18040 15016 18068
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 15148 18028 15154 18080
rect 15206 18077 15212 18080
rect 15206 18071 15255 18077
rect 15206 18037 15209 18071
rect 15243 18037 15255 18071
rect 15206 18031 15255 18037
rect 15206 18028 15212 18031
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 15654 18068 15660 18080
rect 15344 18040 15660 18068
rect 15344 18028 15350 18040
rect 15654 18028 15660 18040
rect 15712 18028 15718 18080
rect 15930 18028 15936 18080
rect 15988 18068 15994 18080
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15988 18040 16037 18068
rect 15988 18028 15994 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 17313 18071 17371 18077
rect 17313 18068 17325 18071
rect 16356 18040 17325 18068
rect 16356 18028 16362 18040
rect 17313 18037 17325 18040
rect 17359 18037 17371 18071
rect 17313 18031 17371 18037
rect 17402 18028 17408 18080
rect 17460 18068 17466 18080
rect 20346 18068 20352 18080
rect 17460 18040 20352 18068
rect 17460 18028 17466 18040
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 21818 18028 21824 18080
rect 21876 18068 21882 18080
rect 22922 18068 22928 18080
rect 21876 18040 22928 18068
rect 21876 18028 21882 18040
rect 22922 18028 22928 18040
rect 22980 18028 22986 18080
rect 23750 18068 23756 18080
rect 23711 18040 23756 18068
rect 23750 18028 23756 18040
rect 23808 18028 23814 18080
rect 24670 18068 24676 18080
rect 24631 18040 24676 18068
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 24857 18071 24915 18077
rect 24857 18037 24869 18071
rect 24903 18068 24915 18071
rect 28460 18068 28488 18108
rect 29822 18096 29828 18108
rect 29880 18096 29886 18148
rect 30742 18096 30748 18148
rect 30800 18136 30806 18148
rect 32214 18136 32220 18148
rect 30800 18108 32220 18136
rect 30800 18096 30806 18108
rect 32214 18096 32220 18108
rect 32272 18096 32278 18148
rect 24903 18040 28488 18068
rect 24903 18037 24915 18040
rect 24857 18031 24915 18037
rect 29270 18028 29276 18080
rect 29328 18068 29334 18080
rect 32306 18068 32312 18080
rect 29328 18040 32312 18068
rect 29328 18028 29334 18040
rect 32306 18028 32312 18040
rect 32364 18028 32370 18080
rect 1104 17978 31832 18000
rect 1104 17926 4791 17978
rect 4843 17926 4855 17978
rect 4907 17926 4919 17978
rect 4971 17926 4983 17978
rect 5035 17926 5047 17978
rect 5099 17926 12473 17978
rect 12525 17926 12537 17978
rect 12589 17926 12601 17978
rect 12653 17926 12665 17978
rect 12717 17926 12729 17978
rect 12781 17926 20155 17978
rect 20207 17926 20219 17978
rect 20271 17926 20283 17978
rect 20335 17926 20347 17978
rect 20399 17926 20411 17978
rect 20463 17926 27837 17978
rect 27889 17926 27901 17978
rect 27953 17926 27965 17978
rect 28017 17926 28029 17978
rect 28081 17926 28093 17978
rect 28145 17926 31832 17978
rect 1104 17904 31832 17926
rect 9309 17867 9367 17873
rect 9309 17833 9321 17867
rect 9355 17864 9367 17867
rect 9950 17864 9956 17876
rect 9355 17836 9956 17864
rect 9355 17833 9367 17836
rect 9309 17827 9367 17833
rect 9950 17824 9956 17836
rect 10008 17824 10014 17876
rect 12161 17867 12219 17873
rect 12161 17833 12173 17867
rect 12207 17864 12219 17867
rect 14550 17864 14556 17876
rect 12207 17836 14556 17864
rect 12207 17833 12219 17836
rect 12161 17827 12219 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 14737 17867 14795 17873
rect 14737 17833 14749 17867
rect 14783 17864 14795 17867
rect 15562 17864 15568 17876
rect 14783 17836 15240 17864
rect 14783 17833 14795 17836
rect 14737 17827 14795 17833
rect 15212 17808 15240 17836
rect 15396 17836 15568 17864
rect 15102 17796 15108 17808
rect 12360 17768 15108 17796
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 8619 17632 10885 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 10873 17629 10885 17632
rect 10919 17660 10931 17663
rect 11514 17660 11520 17672
rect 10919 17632 11520 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 12158 17660 12164 17672
rect 12119 17632 12164 17660
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 12360 17669 12388 17768
rect 15102 17756 15108 17768
rect 15160 17756 15166 17808
rect 15194 17756 15200 17808
rect 15252 17756 15258 17808
rect 12986 17688 12992 17740
rect 13044 17728 13050 17740
rect 15396 17728 15424 17836
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 15657 17867 15715 17873
rect 15657 17833 15669 17867
rect 15703 17864 15715 17867
rect 15930 17864 15936 17876
rect 15703 17836 15936 17864
rect 15703 17833 15715 17836
rect 15657 17827 15715 17833
rect 15930 17824 15936 17836
rect 15988 17864 15994 17876
rect 16666 17864 16672 17876
rect 15988 17836 16672 17864
rect 15988 17824 15994 17836
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 16850 17824 16856 17876
rect 16908 17864 16914 17876
rect 17954 17864 17960 17876
rect 16908 17836 17960 17864
rect 16908 17824 16914 17836
rect 17954 17824 17960 17836
rect 18012 17864 18018 17876
rect 22002 17864 22008 17876
rect 18012 17836 22008 17864
rect 18012 17824 18018 17836
rect 22002 17824 22008 17836
rect 22060 17864 22066 17876
rect 23017 17867 23075 17873
rect 23017 17864 23029 17867
rect 22060 17836 23029 17864
rect 22060 17824 22066 17836
rect 23017 17833 23029 17836
rect 23063 17833 23075 17867
rect 23017 17827 23075 17833
rect 23106 17824 23112 17876
rect 23164 17864 23170 17876
rect 25038 17864 25044 17876
rect 23164 17836 25044 17864
rect 23164 17824 23170 17836
rect 25038 17824 25044 17836
rect 25096 17824 25102 17876
rect 25498 17824 25504 17876
rect 25556 17864 25562 17876
rect 26878 17864 26884 17876
rect 25556 17836 26884 17864
rect 25556 17824 25562 17836
rect 26878 17824 26884 17836
rect 26936 17824 26942 17876
rect 28166 17864 28172 17876
rect 27724 17836 28028 17864
rect 28127 17836 28172 17864
rect 16114 17796 16120 17808
rect 15488 17768 16120 17796
rect 15488 17737 15516 17768
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 16224 17768 16436 17796
rect 13044 17700 15424 17728
rect 15473 17731 15531 17737
rect 13044 17688 13050 17700
rect 15473 17697 15485 17731
rect 15519 17697 15531 17731
rect 15473 17691 15531 17697
rect 15562 17688 15568 17740
rect 15620 17728 15626 17740
rect 16224 17728 16252 17768
rect 15620 17700 16252 17728
rect 16408 17728 16436 17768
rect 16574 17756 16580 17808
rect 16632 17796 16638 17808
rect 17586 17796 17592 17808
rect 16632 17768 17592 17796
rect 16632 17756 16638 17768
rect 17586 17756 17592 17768
rect 17644 17756 17650 17808
rect 19610 17796 19616 17808
rect 18892 17768 19616 17796
rect 18892 17737 18920 17768
rect 19610 17756 19616 17768
rect 19668 17796 19674 17808
rect 21082 17796 21088 17808
rect 19668 17768 21088 17796
rect 19668 17756 19674 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 22833 17799 22891 17805
rect 22833 17765 22845 17799
rect 22879 17765 22891 17799
rect 22833 17759 22891 17765
rect 18601 17731 18659 17737
rect 18601 17728 18613 17731
rect 16408 17700 18613 17728
rect 15620 17688 15626 17700
rect 18601 17697 18613 17700
rect 18647 17697 18659 17731
rect 18601 17691 18659 17697
rect 18877 17731 18935 17737
rect 18877 17697 18889 17731
rect 18923 17697 18935 17731
rect 18877 17691 18935 17697
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 22097 17731 22155 17737
rect 22097 17728 22109 17731
rect 19300 17700 22109 17728
rect 19300 17688 19306 17700
rect 22097 17697 22109 17700
rect 22143 17697 22155 17731
rect 22370 17728 22376 17740
rect 22331 17700 22376 17728
rect 22097 17691 22155 17697
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 22520 17700 22600 17728
rect 22520 17688 22526 17700
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17660 12863 17663
rect 15010 17660 15016 17672
rect 12851 17632 15016 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17660 15439 17663
rect 15746 17660 15752 17672
rect 15427 17632 15752 17660
rect 15427 17629 15439 17632
rect 15381 17623 15439 17629
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 16298 17669 16304 17672
rect 16275 17663 16304 17669
rect 16275 17660 16287 17663
rect 15896 17632 16287 17660
rect 15896 17620 15902 17632
rect 16275 17629 16287 17632
rect 16275 17623 16304 17629
rect 16298 17620 16304 17623
rect 16356 17620 16362 17672
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 16577 17663 16635 17669
rect 16577 17629 16589 17663
rect 16623 17660 16635 17663
rect 17310 17660 17316 17672
rect 16623 17632 17316 17660
rect 16623 17629 16635 17632
rect 16577 17623 16635 17629
rect 10965 17595 11023 17601
rect 10965 17561 10977 17595
rect 11011 17592 11023 17595
rect 13446 17592 13452 17604
rect 11011 17564 13452 17592
rect 11011 17561 11023 17564
rect 10965 17555 11023 17561
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 13630 17592 13636 17604
rect 13591 17564 13636 17592
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 14274 17552 14280 17604
rect 14332 17592 14338 17604
rect 14369 17595 14427 17601
rect 14369 17592 14381 17595
rect 14332 17564 14381 17592
rect 14332 17552 14338 17564
rect 14369 17561 14381 17564
rect 14415 17561 14427 17595
rect 14550 17592 14556 17604
rect 14511 17564 14556 17592
rect 14369 17555 14427 17561
rect 14550 17552 14556 17564
rect 14608 17552 14614 17604
rect 14660 17564 15424 17592
rect 9858 17524 9864 17536
rect 9819 17496 9864 17524
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 10410 17524 10416 17536
rect 10371 17496 10416 17524
rect 10410 17484 10416 17496
rect 10468 17484 10474 17536
rect 11606 17524 11612 17536
rect 11567 17496 11612 17524
rect 11606 17484 11612 17496
rect 11664 17484 11670 17536
rect 12986 17524 12992 17536
rect 12947 17496 12992 17524
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 13541 17527 13599 17533
rect 13541 17524 13553 17527
rect 13320 17496 13553 17524
rect 13320 17484 13326 17496
rect 13541 17493 13553 17496
rect 13587 17493 13599 17527
rect 13541 17487 13599 17493
rect 13722 17484 13728 17536
rect 13780 17524 13786 17536
rect 14660 17524 14688 17564
rect 15194 17524 15200 17536
rect 13780 17496 14688 17524
rect 15155 17496 15200 17524
rect 13780 17484 13786 17496
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 15396 17524 15424 17564
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 15657 17595 15715 17601
rect 15657 17592 15669 17595
rect 15620 17564 15669 17592
rect 15620 17552 15626 17564
rect 15657 17561 15669 17564
rect 15703 17561 15715 17595
rect 15657 17555 15715 17561
rect 15930 17552 15936 17604
rect 15988 17592 15994 17604
rect 16408 17592 16436 17623
rect 15988 17564 16436 17592
rect 16500 17592 16528 17623
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 19392 17632 19441 17660
rect 19392 17620 19398 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 19429 17623 19487 17629
rect 19536 17632 19625 17660
rect 16758 17592 16764 17604
rect 16500 17564 16764 17592
rect 15988 17552 15994 17564
rect 16758 17552 16764 17564
rect 16816 17552 16822 17604
rect 16942 17552 16948 17604
rect 17000 17592 17006 17604
rect 19536 17592 19564 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 19720 17592 19748 17623
rect 19794 17620 19800 17672
rect 19852 17660 19858 17672
rect 20714 17660 20720 17672
rect 19852 17632 20720 17660
rect 19852 17620 19858 17632
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 22572 17660 22600 17700
rect 22646 17688 22652 17740
rect 22704 17728 22710 17740
rect 22848 17728 22876 17759
rect 23566 17756 23572 17808
rect 23624 17796 23630 17808
rect 23624 17768 25452 17796
rect 23624 17756 23630 17768
rect 22704 17700 22876 17728
rect 22704 17688 22710 17700
rect 22922 17688 22928 17740
rect 22980 17728 22986 17740
rect 23477 17731 23535 17737
rect 23477 17728 23489 17731
rect 22980 17700 23489 17728
rect 22980 17688 22986 17700
rect 23477 17697 23489 17700
rect 23523 17697 23535 17731
rect 23477 17691 23535 17697
rect 23676 17700 25084 17728
rect 23017 17663 23075 17669
rect 23017 17660 23029 17663
rect 22572 17632 23029 17660
rect 23017 17629 23029 17632
rect 23063 17629 23075 17663
rect 23017 17623 23075 17629
rect 23385 17663 23443 17669
rect 23385 17629 23397 17663
rect 23431 17629 23443 17663
rect 23385 17623 23443 17629
rect 17000 17564 17434 17592
rect 18248 17564 19564 17592
rect 19628 17564 19748 17592
rect 17000 17552 17006 17564
rect 18248 17536 18276 17564
rect 16117 17527 16175 17533
rect 16117 17524 16129 17527
rect 15396 17496 16129 17524
rect 16117 17493 16129 17496
rect 16163 17493 16175 17527
rect 16117 17487 16175 17493
rect 16206 17484 16212 17536
rect 16264 17524 16270 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 16264 17496 17141 17524
rect 16264 17484 16270 17496
rect 17129 17493 17141 17496
rect 17175 17524 17187 17527
rect 17678 17524 17684 17536
rect 17175 17496 17684 17524
rect 17175 17493 17187 17496
rect 17129 17487 17187 17493
rect 17678 17484 17684 17496
rect 17736 17524 17742 17536
rect 17954 17524 17960 17536
rect 17736 17496 17960 17524
rect 17736 17484 17742 17496
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 18230 17484 18236 17536
rect 18288 17484 18294 17536
rect 19518 17484 19524 17536
rect 19576 17524 19582 17536
rect 19628 17524 19656 17564
rect 20162 17552 20168 17604
rect 20220 17592 20226 17604
rect 20806 17592 20812 17604
rect 20220 17564 20812 17592
rect 20220 17552 20226 17564
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 23400 17592 23428 17623
rect 22572 17564 23428 17592
rect 19576 17496 19656 17524
rect 19576 17484 19582 17496
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 20073 17527 20131 17533
rect 20073 17524 20085 17527
rect 19760 17496 20085 17524
rect 19760 17484 19766 17496
rect 20073 17493 20085 17496
rect 20119 17493 20131 17527
rect 20622 17524 20628 17536
rect 20583 17496 20628 17524
rect 20073 17487 20131 17493
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 22572 17524 22600 17564
rect 20772 17496 22600 17524
rect 20772 17484 20778 17496
rect 22646 17484 22652 17536
rect 22704 17524 22710 17536
rect 23676 17524 23704 17700
rect 25056 17669 25084 17700
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17629 24915 17663
rect 24857 17623 24915 17629
rect 24949 17663 25007 17669
rect 24949 17629 24961 17663
rect 24995 17629 25007 17663
rect 24949 17623 25007 17629
rect 25041 17663 25099 17669
rect 25041 17629 25053 17663
rect 25087 17629 25099 17663
rect 25222 17660 25228 17672
rect 25183 17632 25228 17660
rect 25041 17623 25099 17629
rect 24578 17524 24584 17536
rect 22704 17496 23704 17524
rect 24539 17496 24584 17524
rect 22704 17484 22710 17496
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 24872 17524 24900 17623
rect 24964 17592 24992 17623
rect 25222 17620 25228 17632
rect 25280 17620 25286 17672
rect 25424 17660 25452 17768
rect 25590 17756 25596 17808
rect 25648 17796 25654 17808
rect 25685 17799 25743 17805
rect 25685 17796 25697 17799
rect 25648 17768 25697 17796
rect 25648 17756 25654 17768
rect 25685 17765 25697 17768
rect 25731 17765 25743 17799
rect 27724 17796 27752 17836
rect 25685 17759 25743 17765
rect 25792 17768 27752 17796
rect 28000 17796 28028 17836
rect 28166 17824 28172 17836
rect 28224 17824 28230 17876
rect 30466 17864 30472 17876
rect 28276 17836 30472 17864
rect 28276 17796 28304 17836
rect 30466 17824 30472 17836
rect 30524 17824 30530 17876
rect 28000 17768 28304 17796
rect 25792 17740 25820 17768
rect 28350 17756 28356 17808
rect 28408 17796 28414 17808
rect 30742 17796 30748 17808
rect 28408 17768 30748 17796
rect 28408 17756 28414 17768
rect 30742 17756 30748 17768
rect 30800 17756 30806 17808
rect 25498 17688 25504 17740
rect 25556 17728 25562 17740
rect 25774 17728 25780 17740
rect 25556 17700 25780 17728
rect 25556 17688 25562 17700
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 26510 17728 26516 17740
rect 26200 17700 26516 17728
rect 26200 17688 26206 17700
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 27614 17728 27620 17740
rect 26896 17700 27620 17728
rect 26050 17660 26056 17672
rect 25424 17632 26056 17660
rect 26050 17620 26056 17632
rect 26108 17620 26114 17672
rect 26896 17669 26924 17700
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 27706 17688 27712 17740
rect 27764 17728 27770 17740
rect 28997 17731 29055 17737
rect 27764 17700 27809 17728
rect 27764 17688 27770 17700
rect 28997 17697 29009 17731
rect 29043 17728 29055 17731
rect 29546 17728 29552 17740
rect 29043 17700 29552 17728
rect 29043 17697 29055 17700
rect 28997 17691 29055 17697
rect 29546 17688 29552 17700
rect 29604 17688 29610 17740
rect 29730 17688 29736 17740
rect 29788 17688 29794 17740
rect 30009 17731 30067 17737
rect 30009 17697 30021 17731
rect 30055 17728 30067 17731
rect 31294 17728 31300 17740
rect 30055 17700 31300 17728
rect 30055 17697 30067 17700
rect 30009 17691 30067 17697
rect 31294 17688 31300 17700
rect 31352 17688 31358 17740
rect 26881 17663 26939 17669
rect 26881 17629 26893 17663
rect 26927 17629 26939 17663
rect 26881 17623 26939 17629
rect 27249 17663 27307 17669
rect 27249 17629 27261 17663
rect 27295 17660 27307 17663
rect 27430 17660 27436 17672
rect 27295 17632 27436 17660
rect 27295 17629 27307 17632
rect 27249 17623 27307 17629
rect 27430 17620 27436 17632
rect 27488 17620 27494 17672
rect 28074 17660 28080 17672
rect 28035 17632 28080 17660
rect 28074 17620 28080 17632
rect 28132 17620 28138 17672
rect 29086 17620 29092 17672
rect 29144 17660 29150 17672
rect 29181 17663 29239 17669
rect 29181 17660 29193 17663
rect 29144 17632 29193 17660
rect 29144 17620 29150 17632
rect 29181 17629 29193 17632
rect 29227 17660 29239 17663
rect 29748 17660 29776 17688
rect 30193 17663 30251 17669
rect 30193 17660 30205 17663
rect 29227 17632 30205 17660
rect 29227 17629 29239 17632
rect 29181 17623 29239 17629
rect 30193 17629 30205 17632
rect 30239 17629 30251 17663
rect 30193 17623 30251 17629
rect 30466 17620 30472 17672
rect 30524 17660 30530 17672
rect 30653 17663 30711 17669
rect 30653 17660 30665 17663
rect 30524 17632 30665 17660
rect 30524 17620 30530 17632
rect 30653 17629 30665 17632
rect 30699 17629 30711 17663
rect 30653 17623 30711 17629
rect 30742 17620 30748 17672
rect 30800 17660 30806 17672
rect 30837 17663 30895 17669
rect 30837 17660 30849 17663
rect 30800 17632 30849 17660
rect 30800 17620 30806 17632
rect 30837 17629 30849 17632
rect 30883 17629 30895 17663
rect 30837 17623 30895 17629
rect 25774 17592 25780 17604
rect 24964 17564 25780 17592
rect 25774 17552 25780 17564
rect 25832 17552 25838 17604
rect 25869 17595 25927 17601
rect 25869 17561 25881 17595
rect 25915 17592 25927 17595
rect 26142 17592 26148 17604
rect 25915 17564 26148 17592
rect 25915 17561 25927 17564
rect 25869 17555 25927 17561
rect 26142 17552 26148 17564
rect 26200 17552 26206 17604
rect 26234 17552 26240 17604
rect 26292 17592 26298 17604
rect 26292 17564 26337 17592
rect 26292 17552 26298 17564
rect 26786 17552 26792 17604
rect 26844 17552 26850 17604
rect 26970 17592 26976 17604
rect 26931 17564 26976 17592
rect 26970 17552 26976 17564
rect 27028 17552 27034 17604
rect 27065 17595 27123 17601
rect 27065 17561 27077 17595
rect 27111 17561 27123 17595
rect 27065 17555 27123 17561
rect 25958 17524 25964 17536
rect 24872 17496 25964 17524
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 26694 17524 26700 17536
rect 26655 17496 26700 17524
rect 26694 17484 26700 17496
rect 26752 17484 26758 17536
rect 26804 17524 26832 17552
rect 27080 17524 27108 17555
rect 27522 17552 27528 17604
rect 27580 17592 27586 17604
rect 29362 17592 29368 17604
rect 27580 17564 29368 17592
rect 27580 17552 27586 17564
rect 29362 17552 29368 17564
rect 29420 17552 29426 17604
rect 29730 17552 29736 17604
rect 29788 17592 29794 17604
rect 31570 17592 31576 17604
rect 29788 17564 31576 17592
rect 29788 17552 29794 17564
rect 31570 17552 31576 17564
rect 31628 17552 31634 17604
rect 26804 17496 27108 17524
rect 27893 17527 27951 17533
rect 27893 17493 27905 17527
rect 27939 17524 27951 17527
rect 28258 17524 28264 17536
rect 27939 17496 28264 17524
rect 27939 17493 27951 17496
rect 27893 17487 27951 17493
rect 28258 17484 28264 17496
rect 28316 17484 28322 17536
rect 28534 17484 28540 17536
rect 28592 17524 28598 17536
rect 29270 17524 29276 17536
rect 28592 17496 29276 17524
rect 28592 17484 28598 17496
rect 29270 17484 29276 17496
rect 29328 17484 29334 17536
rect 30006 17484 30012 17536
rect 30064 17524 30070 17536
rect 31021 17527 31079 17533
rect 31021 17524 31033 17527
rect 30064 17496 31033 17524
rect 30064 17484 30070 17496
rect 31021 17493 31033 17496
rect 31067 17493 31079 17527
rect 31021 17487 31079 17493
rect 31294 17484 31300 17536
rect 31352 17524 31358 17536
rect 31662 17524 31668 17536
rect 31352 17496 31668 17524
rect 31352 17484 31358 17496
rect 31662 17484 31668 17496
rect 31720 17484 31726 17536
rect 1104 17434 31992 17456
rect 1104 17382 8632 17434
rect 8684 17382 8696 17434
rect 8748 17382 8760 17434
rect 8812 17382 8824 17434
rect 8876 17382 8888 17434
rect 8940 17382 16314 17434
rect 16366 17382 16378 17434
rect 16430 17382 16442 17434
rect 16494 17382 16506 17434
rect 16558 17382 16570 17434
rect 16622 17382 23996 17434
rect 24048 17382 24060 17434
rect 24112 17382 24124 17434
rect 24176 17382 24188 17434
rect 24240 17382 24252 17434
rect 24304 17382 31678 17434
rect 31730 17382 31742 17434
rect 31794 17382 31806 17434
rect 31858 17382 31870 17434
rect 31922 17382 31934 17434
rect 31986 17382 31992 17434
rect 1104 17360 31992 17382
rect 9953 17323 10011 17329
rect 9953 17289 9965 17323
rect 9999 17320 10011 17323
rect 10962 17320 10968 17332
rect 9999 17292 10968 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 13630 17280 13636 17332
rect 13688 17320 13694 17332
rect 13688 17292 14044 17320
rect 13688 17280 13694 17292
rect 12529 17255 12587 17261
rect 12529 17221 12541 17255
rect 12575 17252 12587 17255
rect 12894 17252 12900 17264
rect 12575 17224 12900 17252
rect 12575 17221 12587 17224
rect 12529 17215 12587 17221
rect 12894 17212 12900 17224
rect 12952 17212 12958 17264
rect 13081 17255 13139 17261
rect 13081 17221 13093 17255
rect 13127 17252 13139 17255
rect 13170 17252 13176 17264
rect 13127 17224 13176 17252
rect 13127 17221 13139 17224
rect 13081 17215 13139 17221
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 13262 17212 13268 17264
rect 13320 17261 13326 17264
rect 13320 17255 13339 17261
rect 13327 17221 13339 17255
rect 13320 17215 13339 17221
rect 13909 17255 13967 17261
rect 13909 17221 13921 17255
rect 13955 17221 13967 17255
rect 14016 17252 14044 17292
rect 14090 17280 14096 17332
rect 14148 17329 14154 17332
rect 14148 17323 14167 17329
rect 14155 17289 14167 17323
rect 14829 17323 14887 17329
rect 14829 17320 14841 17323
rect 14148 17283 14167 17289
rect 14200 17292 14841 17320
rect 14148 17280 14154 17283
rect 14200 17252 14228 17292
rect 14829 17289 14841 17292
rect 14875 17289 14887 17323
rect 14829 17283 14887 17289
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 16301 17323 16359 17329
rect 15252 17292 16252 17320
rect 15252 17280 15258 17292
rect 14016 17224 14228 17252
rect 13909 17215 13967 17221
rect 13320 17212 13326 17215
rect 10962 17184 10968 17196
rect 10923 17156 10968 17184
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 11330 17144 11336 17196
rect 11388 17184 11394 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11388 17156 11713 17184
rect 11388 17144 11394 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 12342 17184 12348 17196
rect 12303 17156 12348 17184
rect 11701 17147 11759 17153
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 12618 17184 12624 17196
rect 12579 17156 12624 17184
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 13924 17184 13952 17215
rect 15470 17212 15476 17264
rect 15528 17252 15534 17264
rect 16224 17252 16252 17292
rect 16301 17289 16313 17323
rect 16347 17320 16359 17323
rect 16942 17320 16948 17332
rect 16347 17292 16948 17320
rect 16347 17289 16359 17292
rect 16301 17283 16359 17289
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 17129 17323 17187 17329
rect 17129 17289 17141 17323
rect 17175 17320 17187 17323
rect 17175 17292 17254 17320
rect 17175 17289 17187 17292
rect 17129 17283 17187 17289
rect 17226 17252 17254 17292
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 18966 17320 18972 17332
rect 17552 17292 18972 17320
rect 17552 17280 17558 17292
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 19484 17292 21097 17320
rect 19484 17280 19490 17292
rect 21085 17289 21097 17292
rect 21131 17289 21143 17323
rect 23934 17320 23940 17332
rect 21085 17283 21143 17289
rect 21252 17292 23940 17320
rect 17402 17252 17408 17264
rect 15528 17224 15976 17252
rect 16224 17224 17172 17252
rect 17226 17224 17408 17252
rect 15528 17212 15534 17224
rect 14642 17184 14648 17196
rect 13924 17156 14648 17184
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17184 14795 17187
rect 14918 17184 14924 17196
rect 14783 17156 14924 17184
rect 14783 17153 14795 17156
rect 14737 17147 14795 17153
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15378 17184 15384 17196
rect 15068 17156 15384 17184
rect 15068 17144 15074 17156
rect 15378 17144 15384 17156
rect 15436 17184 15442 17196
rect 15948 17193 15976 17224
rect 15657 17190 15715 17193
rect 15580 17187 15715 17190
rect 15580 17184 15669 17187
rect 15436 17162 15669 17184
rect 15436 17156 15608 17162
rect 15436 17144 15442 17156
rect 15657 17153 15669 17162
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 15820 17187 15878 17193
rect 15820 17153 15832 17187
rect 15866 17184 15878 17187
rect 15933 17187 15991 17193
rect 15866 17153 15884 17184
rect 15820 17147 15884 17153
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17184 16083 17187
rect 16666 17184 16672 17196
rect 16071 17156 16672 17184
rect 16071 17153 16083 17156
rect 16025 17147 16083 17153
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17116 9459 17119
rect 11514 17116 11520 17128
rect 9447 17088 11520 17116
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17116 11851 17119
rect 15105 17119 15163 17125
rect 11839 17088 15056 17116
rect 11839 17085 11851 17088
rect 11793 17079 11851 17085
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 11057 17051 11115 17057
rect 9732 17020 10548 17048
rect 9732 17008 9738 17020
rect 10520 16992 10548 17020
rect 11057 17017 11069 17051
rect 11103 17048 11115 17051
rect 12250 17048 12256 17060
rect 11103 17020 12256 17048
rect 11103 17017 11115 17020
rect 11057 17011 11115 17017
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 13170 17008 13176 17060
rect 13228 17048 13234 17060
rect 13449 17051 13507 17057
rect 13449 17048 13461 17051
rect 13228 17020 13461 17048
rect 13228 17008 13234 17020
rect 13449 17017 13461 17020
rect 13495 17017 13507 17051
rect 15028 17048 15056 17088
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15286 17116 15292 17128
rect 15151 17088 15292 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 15856 17116 15884 17147
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 17144 17193 17172 17224
rect 17402 17212 17408 17224
rect 17460 17212 17466 17264
rect 17770 17212 17776 17264
rect 17828 17252 17834 17264
rect 18322 17252 18328 17264
rect 17828 17224 18328 17252
rect 17828 17212 17834 17224
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 20349 17255 20407 17261
rect 20349 17221 20361 17255
rect 20395 17252 20407 17255
rect 20622 17252 20628 17264
rect 20395 17224 20628 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 20622 17212 20628 17224
rect 20680 17212 20686 17264
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 21252 17261 21280 17292
rect 23934 17280 23940 17292
rect 23992 17280 23998 17332
rect 24486 17280 24492 17332
rect 24544 17320 24550 17332
rect 27157 17323 27215 17329
rect 27157 17320 27169 17323
rect 24544 17292 27169 17320
rect 24544 17280 24550 17292
rect 27157 17289 27169 17292
rect 27203 17289 27215 17323
rect 28166 17320 28172 17332
rect 27157 17283 27215 17289
rect 27264 17292 28172 17320
rect 21237 17255 21295 17261
rect 21237 17252 21249 17255
rect 20864 17224 21249 17252
rect 20864 17212 20870 17224
rect 21237 17221 21249 17224
rect 21283 17221 21295 17255
rect 21237 17215 21295 17221
rect 21453 17255 21511 17261
rect 21453 17221 21465 17255
rect 21499 17252 21511 17255
rect 21726 17252 21732 17264
rect 21499 17224 21732 17252
rect 21499 17221 21511 17224
rect 21453 17215 21511 17221
rect 21726 17212 21732 17224
rect 21784 17212 21790 17264
rect 22922 17212 22928 17264
rect 22980 17212 22986 17264
rect 23569 17255 23627 17261
rect 23569 17221 23581 17255
rect 23615 17252 23627 17255
rect 24670 17252 24676 17264
rect 23615 17224 24676 17252
rect 23615 17221 23627 17224
rect 23569 17215 23627 17221
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 25038 17212 25044 17264
rect 25096 17212 25102 17264
rect 26510 17212 26516 17264
rect 26568 17252 26574 17264
rect 26694 17252 26700 17264
rect 26568 17224 26700 17252
rect 26568 17212 26574 17224
rect 26694 17212 26700 17224
rect 26752 17212 26758 17264
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16766 17156 16865 17184
rect 16482 17116 16488 17128
rect 15856 17088 16488 17116
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 16766 17116 16794 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17153 17187 17187
rect 21082 17184 21088 17196
rect 17129 17147 17187 17153
rect 17226 17156 19274 17184
rect 20640 17156 21088 17184
rect 17226 17116 17254 17156
rect 16632 17088 16794 17116
rect 16868 17088 17254 17116
rect 16632 17076 16638 17088
rect 15028 17020 15700 17048
rect 13449 17011 13507 17017
rect 15672 16992 15700 17020
rect 15838 17008 15844 17060
rect 15896 17048 15902 17060
rect 16868 17048 16896 17088
rect 17402 17076 17408 17128
rect 17460 17116 17466 17128
rect 17862 17116 17868 17128
rect 17460 17088 17868 17116
rect 17460 17076 17466 17088
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18414 17125 18420 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 18012 17088 18153 17116
rect 18012 17076 18018 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18371 17119 18420 17125
rect 18371 17116 18383 17119
rect 18141 17079 18199 17085
rect 18248 17088 18383 17116
rect 17034 17048 17040 17060
rect 15896 17020 16896 17048
rect 16995 17020 17040 17048
rect 15896 17008 15902 17020
rect 17034 17008 17040 17020
rect 17092 17008 17098 17060
rect 18248 17048 18276 17088
rect 18371 17085 18383 17088
rect 18417 17085 18420 17119
rect 18371 17079 18420 17085
rect 18414 17076 18420 17079
rect 18472 17076 18478 17128
rect 18506 17076 18512 17128
rect 18564 17116 18570 17128
rect 20640 17125 20668 17156
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17184 23903 17187
rect 24026 17184 24032 17196
rect 23891 17156 24032 17184
rect 23891 17153 23903 17156
rect 23845 17147 23903 17153
rect 24026 17144 24032 17156
rect 24084 17144 24090 17196
rect 27264 17184 27292 17292
rect 28166 17280 28172 17292
rect 28224 17280 28230 17332
rect 28534 17280 28540 17332
rect 28592 17320 28598 17332
rect 28629 17323 28687 17329
rect 28629 17320 28641 17323
rect 28592 17292 28641 17320
rect 28592 17280 28598 17292
rect 28629 17289 28641 17292
rect 28675 17289 28687 17323
rect 28629 17283 28687 17289
rect 28902 17280 28908 17332
rect 28960 17280 28966 17332
rect 29178 17280 29184 17332
rect 29236 17320 29242 17332
rect 30377 17323 30435 17329
rect 29236 17292 30328 17320
rect 29236 17280 29242 17292
rect 27430 17252 27436 17264
rect 25792 17156 27292 17184
rect 27367 17224 27436 17252
rect 20625 17119 20683 17125
rect 18564 17088 20576 17116
rect 18564 17076 18570 17088
rect 17604 17020 18276 17048
rect 20548 17048 20576 17088
rect 20625 17085 20637 17119
rect 20671 17085 20683 17119
rect 22830 17116 22836 17128
rect 20625 17079 20683 17085
rect 20732 17088 22836 17116
rect 20732 17048 20760 17088
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 23014 17076 23020 17128
rect 23072 17116 23078 17128
rect 24305 17119 24363 17125
rect 23072 17088 23796 17116
rect 23072 17076 23078 17088
rect 20548 17020 20760 17048
rect 10502 16980 10508 16992
rect 10463 16952 10508 16980
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 12158 16940 12164 16992
rect 12216 16980 12222 16992
rect 12345 16983 12403 16989
rect 12345 16980 12357 16983
rect 12216 16952 12357 16980
rect 12216 16940 12222 16952
rect 12345 16949 12357 16952
rect 12391 16949 12403 16983
rect 12345 16943 12403 16949
rect 13265 16983 13323 16989
rect 13265 16949 13277 16983
rect 13311 16980 13323 16983
rect 13722 16980 13728 16992
rect 13311 16952 13728 16980
rect 13311 16949 13323 16952
rect 13265 16943 13323 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 14274 16980 14280 16992
rect 14235 16952 14280 16980
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 15013 16983 15071 16989
rect 15013 16949 15025 16983
rect 15059 16980 15071 16983
rect 15102 16980 15108 16992
rect 15059 16952 15108 16980
rect 15059 16949 15071 16952
rect 15013 16943 15071 16949
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 15252 16952 15297 16980
rect 15252 16940 15258 16952
rect 15654 16940 15660 16992
rect 15712 16940 15718 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 17604 16980 17632 17020
rect 20806 17008 20812 17060
rect 20864 17048 20870 17060
rect 21174 17048 21180 17060
rect 20864 17020 21180 17048
rect 20864 17008 20870 17020
rect 21174 17008 21180 17020
rect 21232 17008 21238 17060
rect 21634 17008 21640 17060
rect 21692 17048 21698 17060
rect 23768 17048 23796 17088
rect 24305 17085 24317 17119
rect 24351 17085 24363 17119
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24305 17079 24363 17085
rect 24412 17088 24593 17116
rect 24320 17048 24348 17079
rect 21692 17020 22600 17048
rect 23768 17020 24348 17048
rect 21692 17008 21698 17020
rect 16080 16952 17632 16980
rect 16080 16940 16086 16952
rect 17678 16940 17684 16992
rect 17736 16980 17742 16992
rect 18138 16980 18144 16992
rect 17736 16952 18144 16980
rect 17736 16940 17742 16952
rect 18138 16940 18144 16952
rect 18196 16940 18202 16992
rect 18322 16940 18328 16992
rect 18380 16980 18386 16992
rect 18877 16983 18935 16989
rect 18877 16980 18889 16983
rect 18380 16952 18889 16980
rect 18380 16940 18386 16952
rect 18877 16949 18889 16952
rect 18923 16949 18935 16983
rect 18877 16943 18935 16949
rect 19058 16940 19064 16992
rect 19116 16980 19122 16992
rect 21269 16983 21327 16989
rect 21269 16980 21281 16983
rect 19116 16952 21281 16980
rect 19116 16940 19122 16952
rect 21269 16949 21281 16952
rect 21315 16949 21327 16983
rect 21269 16943 21327 16949
rect 21450 16940 21456 16992
rect 21508 16980 21514 16992
rect 22002 16980 22008 16992
rect 21508 16952 22008 16980
rect 21508 16940 21514 16952
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22097 16983 22155 16989
rect 22097 16949 22109 16983
rect 22143 16980 22155 16983
rect 22462 16980 22468 16992
rect 22143 16952 22468 16980
rect 22143 16949 22155 16952
rect 22097 16943 22155 16949
rect 22462 16940 22468 16952
rect 22520 16940 22526 16992
rect 22572 16980 22600 17020
rect 24412 16980 24440 17088
rect 24581 17085 24593 17088
rect 24627 17085 24639 17119
rect 24581 17079 24639 17085
rect 25314 17076 25320 17128
rect 25372 17116 25378 17128
rect 25792 17116 25820 17156
rect 26050 17116 26056 17128
rect 25372 17088 25820 17116
rect 26011 17088 26056 17116
rect 25372 17076 25378 17088
rect 26050 17076 26056 17088
rect 26108 17076 26114 17128
rect 26694 17076 26700 17128
rect 26752 17116 26758 17128
rect 27367 17116 27395 17224
rect 27430 17212 27436 17224
rect 27488 17212 27494 17264
rect 27706 17212 27712 17264
rect 27764 17252 27770 17264
rect 28721 17255 28779 17261
rect 28721 17252 28733 17255
rect 27764 17224 28733 17252
rect 27764 17212 27770 17224
rect 28721 17221 28733 17224
rect 28767 17252 28779 17255
rect 28920 17252 28948 17280
rect 28767 17224 28948 17252
rect 29549 17255 29607 17261
rect 28767 17221 28779 17224
rect 28721 17215 28779 17221
rect 29319 17221 29377 17227
rect 27525 17187 27583 17193
rect 27525 17153 27537 17187
rect 27571 17153 27583 17187
rect 27525 17147 27583 17153
rect 26752 17088 27395 17116
rect 27433 17119 27491 17125
rect 26752 17076 26758 17088
rect 27433 17085 27445 17119
rect 27479 17085 27491 17119
rect 27540 17116 27568 17147
rect 28350 17144 28356 17196
rect 28408 17184 28414 17196
rect 28445 17187 28503 17193
rect 28445 17184 28457 17187
rect 28408 17156 28457 17184
rect 28408 17144 28414 17156
rect 28445 17153 28457 17156
rect 28491 17184 28503 17187
rect 29178 17184 29184 17196
rect 28491 17156 29184 17184
rect 28491 17153 28503 17156
rect 28445 17147 28503 17153
rect 29178 17144 29184 17156
rect 29236 17144 29242 17196
rect 29319 17187 29331 17221
rect 29365 17196 29377 17221
rect 29549 17221 29561 17255
rect 29595 17252 29607 17255
rect 30006 17252 30012 17264
rect 29595 17224 29684 17252
rect 29967 17224 30012 17252
rect 29595 17221 29607 17224
rect 29549 17215 29607 17221
rect 29365 17187 29368 17196
rect 29319 17181 29368 17187
rect 29334 17156 29368 17181
rect 29362 17144 29368 17156
rect 29420 17144 29426 17196
rect 29454 17116 29460 17128
rect 27540 17088 29460 17116
rect 27433 17079 27491 17085
rect 25590 17008 25596 17060
rect 25648 17048 25654 17060
rect 25648 17020 26372 17048
rect 25648 17008 25654 17020
rect 22572 16952 24440 16980
rect 26344 16980 26372 17020
rect 26510 17008 26516 17060
rect 26568 17048 26574 17060
rect 27448 17048 27476 17079
rect 29454 17076 29460 17088
rect 29512 17076 29518 17128
rect 29656 17116 29684 17224
rect 30006 17212 30012 17224
rect 30064 17212 30070 17264
rect 30300 17252 30328 17292
rect 30377 17289 30389 17323
rect 30423 17320 30435 17323
rect 30466 17320 30472 17332
rect 30423 17292 30472 17320
rect 30423 17289 30435 17292
rect 30377 17283 30435 17289
rect 30466 17280 30472 17292
rect 30524 17280 30530 17332
rect 30989 17255 31047 17261
rect 30989 17252 31001 17255
rect 30300 17224 31001 17252
rect 30989 17221 31001 17224
rect 31035 17221 31047 17255
rect 30989 17215 31047 17221
rect 31205 17255 31263 17261
rect 31205 17221 31217 17255
rect 31251 17221 31263 17255
rect 31205 17215 31263 17221
rect 29822 17144 29828 17196
rect 29880 17184 29886 17196
rect 30193 17187 30251 17193
rect 30193 17184 30205 17187
rect 29880 17156 30205 17184
rect 29880 17144 29886 17156
rect 30193 17153 30205 17156
rect 30239 17153 30251 17187
rect 30193 17147 30251 17153
rect 30466 17144 30472 17196
rect 30524 17184 30530 17196
rect 31220 17184 31248 17215
rect 30524 17156 31248 17184
rect 30524 17144 30530 17156
rect 32122 17116 32128 17128
rect 29656 17088 32128 17116
rect 32122 17076 32128 17088
rect 32180 17076 32186 17128
rect 27522 17048 27528 17060
rect 26568 17020 26613 17048
rect 27448 17020 27528 17048
rect 26568 17008 26574 17020
rect 27522 17008 27528 17020
rect 27580 17008 27586 17060
rect 28258 17048 28264 17060
rect 28219 17020 28264 17048
rect 28258 17008 28264 17020
rect 28316 17048 28322 17060
rect 28994 17048 29000 17060
rect 28316 17020 29000 17048
rect 28316 17008 28322 17020
rect 28994 17008 29000 17020
rect 29052 17008 29058 17060
rect 29178 17048 29184 17060
rect 29139 17020 29184 17048
rect 29178 17008 29184 17020
rect 29236 17008 29242 17060
rect 29365 16983 29423 16989
rect 29365 16980 29377 16983
rect 26344 16952 29377 16980
rect 29365 16949 29377 16952
rect 29411 16949 29423 16983
rect 29365 16943 29423 16949
rect 30466 16940 30472 16992
rect 30524 16980 30530 16992
rect 30837 16983 30895 16989
rect 30837 16980 30849 16983
rect 30524 16952 30849 16980
rect 30524 16940 30530 16952
rect 30837 16949 30849 16952
rect 30883 16949 30895 16983
rect 30837 16943 30895 16949
rect 31021 16983 31079 16989
rect 31021 16949 31033 16983
rect 31067 16980 31079 16983
rect 31662 16980 31668 16992
rect 31067 16952 31668 16980
rect 31067 16949 31079 16952
rect 31021 16943 31079 16949
rect 31662 16940 31668 16952
rect 31720 16940 31726 16992
rect 1104 16890 31832 16912
rect 1104 16838 4791 16890
rect 4843 16838 4855 16890
rect 4907 16838 4919 16890
rect 4971 16838 4983 16890
rect 5035 16838 5047 16890
rect 5099 16838 12473 16890
rect 12525 16838 12537 16890
rect 12589 16838 12601 16890
rect 12653 16838 12665 16890
rect 12717 16838 12729 16890
rect 12781 16838 20155 16890
rect 20207 16838 20219 16890
rect 20271 16838 20283 16890
rect 20335 16838 20347 16890
rect 20399 16838 20411 16890
rect 20463 16838 27837 16890
rect 27889 16838 27901 16890
rect 27953 16838 27965 16890
rect 28017 16838 28029 16890
rect 28081 16838 28093 16890
rect 28145 16838 31832 16890
rect 1104 16816 31832 16838
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 11112 16748 11157 16776
rect 11112 16736 11118 16748
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 13446 16776 13452 16788
rect 11664 16748 13452 16776
rect 11664 16736 11670 16748
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 15286 16776 15292 16788
rect 15247 16748 15292 16776
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15838 16736 15844 16788
rect 15896 16776 15902 16788
rect 16206 16776 16212 16788
rect 15896 16748 16212 16776
rect 15896 16736 15902 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16669 16779 16727 16785
rect 16669 16745 16681 16779
rect 16715 16776 16727 16779
rect 16715 16748 19472 16776
rect 16715 16745 16727 16748
rect 16669 16739 16727 16745
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 10410 16708 10416 16720
rect 9916 16680 10416 16708
rect 9916 16668 9922 16680
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 12986 16708 12992 16720
rect 12947 16680 12992 16708
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 13722 16708 13728 16720
rect 13683 16680 13728 16708
rect 13722 16668 13728 16680
rect 13780 16668 13786 16720
rect 14553 16711 14611 16717
rect 14553 16677 14565 16711
rect 14599 16677 14611 16711
rect 14553 16671 14611 16677
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10962 16640 10968 16652
rect 9999 16612 10968 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11606 16640 11612 16652
rect 11567 16612 11612 16640
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 12158 16640 12164 16652
rect 11716 16612 12164 16640
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 11716 16581 11744 16612
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 12820 16612 14412 16640
rect 12820 16581 12848 16612
rect 11517 16575 11575 16581
rect 11517 16572 11529 16575
rect 11296 16544 11529 16572
rect 11296 16532 11302 16544
rect 11517 16541 11529 16544
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 11695 16575 11753 16581
rect 11695 16541 11707 16575
rect 11741 16541 11753 16575
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 11695 16535 11753 16541
rect 12176 16544 12357 16572
rect 12176 16436 12204 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 12805 16575 12863 16581
rect 12805 16541 12817 16575
rect 12851 16541 12863 16575
rect 12805 16535 12863 16541
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16541 13047 16575
rect 13354 16572 13360 16584
rect 12989 16535 13047 16541
rect 13188 16544 13360 16572
rect 12253 16507 12311 16513
rect 12253 16473 12265 16507
rect 12299 16504 12311 16507
rect 12618 16504 12624 16516
rect 12299 16476 12624 16504
rect 12299 16473 12311 16476
rect 12253 16467 12311 16473
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 12710 16464 12716 16516
rect 12768 16504 12774 16516
rect 13004 16504 13032 16535
rect 12768 16476 13032 16504
rect 12768 16464 12774 16476
rect 12986 16436 12992 16448
rect 12176 16408 12992 16436
rect 12986 16396 12992 16408
rect 13044 16436 13050 16448
rect 13188 16436 13216 16544
rect 13354 16532 13360 16544
rect 13412 16572 13418 16584
rect 13449 16575 13507 16581
rect 13449 16572 13461 16575
rect 13412 16544 13461 16572
rect 13412 16532 13418 16544
rect 13449 16541 13461 16544
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 14182 16532 14188 16584
rect 14240 16572 14246 16584
rect 14384 16581 14412 16612
rect 14277 16575 14335 16581
rect 14277 16572 14289 16575
rect 14240 16544 14289 16572
rect 14240 16532 14246 16544
rect 14277 16541 14289 16544
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16572 14427 16575
rect 14458 16572 14464 16584
rect 14415 16544 14464 16572
rect 14415 16541 14427 16544
rect 14369 16535 14427 16541
rect 14458 16532 14464 16544
rect 14516 16532 14522 16584
rect 14568 16572 14596 16671
rect 15194 16668 15200 16720
rect 15252 16708 15258 16720
rect 18874 16708 18880 16720
rect 15252 16680 16414 16708
rect 18835 16680 18880 16708
rect 15252 16668 15258 16680
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 16386 16640 16414 16680
rect 18874 16668 18880 16680
rect 18932 16668 18938 16720
rect 19444 16708 19472 16748
rect 19794 16736 19800 16788
rect 19852 16776 19858 16788
rect 21177 16779 21235 16785
rect 19852 16748 21128 16776
rect 19852 16736 19858 16748
rect 21100 16708 21128 16748
rect 21177 16745 21189 16779
rect 21223 16776 21235 16779
rect 21450 16776 21456 16788
rect 21223 16748 21456 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 21542 16736 21548 16788
rect 21600 16776 21606 16788
rect 23474 16776 23480 16788
rect 21600 16748 23480 16776
rect 21600 16736 21606 16748
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 23934 16776 23940 16788
rect 23895 16748 23940 16776
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 26418 16776 26424 16788
rect 24084 16748 26424 16776
rect 24084 16736 24090 16748
rect 26418 16736 26424 16748
rect 26476 16736 26482 16788
rect 26878 16736 26884 16788
rect 26936 16776 26942 16788
rect 28442 16776 28448 16788
rect 26936 16748 28448 16776
rect 26936 16736 26942 16748
rect 28442 16736 28448 16748
rect 28500 16776 28506 16788
rect 28905 16779 28963 16785
rect 28905 16776 28917 16779
rect 28500 16748 28917 16776
rect 28500 16736 28506 16748
rect 28905 16745 28917 16748
rect 28951 16776 28963 16779
rect 29917 16779 29975 16785
rect 29917 16776 29929 16779
rect 28951 16748 29929 16776
rect 28951 16745 28963 16748
rect 28905 16739 28963 16745
rect 29917 16745 29929 16748
rect 29963 16745 29975 16779
rect 31294 16776 31300 16788
rect 29917 16739 29975 16745
rect 31220 16748 31300 16776
rect 22002 16708 22008 16720
rect 19444 16680 19564 16708
rect 21100 16680 22008 16708
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 15160 16612 16344 16640
rect 16386 16612 17417 16640
rect 15160 16600 15166 16612
rect 14826 16572 14832 16584
rect 14568 16544 14832 16572
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 15010 16572 15016 16584
rect 14971 16544 15016 16572
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 15194 16532 15200 16584
rect 15252 16572 15258 16584
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 15252 16544 15301 16572
rect 15252 16532 15258 16544
rect 15289 16541 15301 16544
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 15396 16572 15792 16582
rect 15930 16572 15936 16584
rect 15396 16554 15936 16572
rect 13725 16507 13783 16513
rect 13725 16473 13737 16507
rect 13771 16473 13783 16507
rect 13725 16467 13783 16473
rect 14553 16507 14611 16513
rect 14553 16473 14565 16507
rect 14599 16504 14611 16507
rect 14642 16504 14648 16516
rect 14599 16476 14648 16504
rect 14599 16473 14611 16476
rect 14553 16467 14611 16473
rect 13044 16408 13216 16436
rect 13044 16396 13050 16408
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 13541 16439 13599 16445
rect 13541 16436 13553 16439
rect 13412 16408 13553 16436
rect 13412 16396 13418 16408
rect 13541 16405 13553 16408
rect 13587 16405 13599 16439
rect 13740 16436 13768 16467
rect 14642 16464 14648 16476
rect 14700 16504 14706 16516
rect 15396 16504 15424 16554
rect 15764 16544 15936 16554
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16022 16532 16028 16584
rect 16080 16572 16086 16584
rect 16206 16572 16212 16584
rect 16080 16544 16125 16572
rect 16167 16544 16212 16572
rect 16080 16532 16086 16544
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16316 16581 16344 16612
rect 17405 16609 17417 16612
rect 17451 16609 17463 16643
rect 17405 16603 17463 16609
rect 17954 16600 17960 16652
rect 18012 16640 18018 16652
rect 19536 16640 19564 16680
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 25590 16708 25596 16720
rect 23492 16680 25596 16708
rect 23492 16652 23520 16680
rect 25590 16668 25596 16680
rect 25648 16668 25654 16720
rect 26326 16668 26332 16720
rect 26384 16708 26390 16720
rect 28258 16708 28264 16720
rect 26384 16680 28264 16708
rect 26384 16668 26390 16680
rect 23109 16643 23167 16649
rect 23109 16640 23121 16643
rect 18012 16612 19288 16640
rect 19536 16612 23121 16640
rect 18012 16600 18018 16612
rect 19260 16584 19288 16612
rect 23109 16609 23121 16612
rect 23155 16609 23167 16643
rect 23109 16603 23167 16609
rect 23474 16600 23480 16652
rect 23532 16600 23538 16652
rect 23768 16612 25268 16640
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16541 16359 16575
rect 16301 16535 16359 16541
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16572 16451 16575
rect 16574 16572 16580 16584
rect 16439 16544 16580 16572
rect 16439 16541 16451 16544
rect 16393 16535 16451 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16942 16572 16948 16584
rect 16724 16544 16948 16572
rect 16724 16532 16730 16544
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17126 16572 17132 16584
rect 17087 16544 17132 16572
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 19242 16572 19248 16584
rect 19155 16544 19248 16572
rect 19242 16532 19248 16544
rect 19300 16572 19306 16584
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 19300 16544 19441 16572
rect 19300 16532 19306 16544
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 21358 16532 21364 16584
rect 21416 16572 21422 16584
rect 23385 16575 23443 16581
rect 21416 16544 21772 16572
rect 21416 16532 21422 16544
rect 17678 16504 17684 16516
rect 14700 16476 15424 16504
rect 16290 16476 17684 16504
rect 14700 16464 14706 16476
rect 14366 16436 14372 16448
rect 13740 16408 14372 16436
rect 13541 16399 13599 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 14458 16396 14464 16448
rect 14516 16436 14522 16448
rect 15470 16436 15476 16448
rect 14516 16408 15476 16436
rect 14516 16396 14522 16408
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15565 16439 15623 16445
rect 15565 16405 15577 16439
rect 15611 16436 15623 16439
rect 15654 16436 15660 16448
rect 15611 16408 15660 16436
rect 15611 16405 15623 16408
rect 15565 16399 15623 16405
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 16022 16396 16028 16448
rect 16080 16436 16086 16448
rect 16290 16436 16318 16476
rect 17678 16464 17684 16476
rect 17736 16464 17742 16516
rect 17954 16464 17960 16516
rect 18012 16464 18018 16516
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19705 16507 19763 16513
rect 19705 16504 19717 16507
rect 19392 16476 19717 16504
rect 19392 16464 19398 16476
rect 19705 16473 19717 16476
rect 19751 16473 19763 16507
rect 19705 16467 19763 16473
rect 19794 16464 19800 16516
rect 19852 16504 19858 16516
rect 21450 16504 21456 16516
rect 19852 16476 20194 16504
rect 21284 16476 21456 16504
rect 19852 16464 19858 16476
rect 16080 16408 16318 16436
rect 16080 16396 16086 16408
rect 16482 16396 16488 16448
rect 16540 16436 16546 16448
rect 21284 16436 21312 16476
rect 21450 16464 21456 16476
rect 21508 16464 21514 16516
rect 16540 16408 21312 16436
rect 16540 16396 16546 16408
rect 21358 16396 21364 16448
rect 21416 16436 21422 16448
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 21416 16408 21649 16436
rect 21416 16396 21422 16408
rect 21637 16405 21649 16408
rect 21683 16405 21695 16439
rect 21744 16436 21772 16544
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 23658 16572 23664 16584
rect 23431 16544 23664 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 23658 16532 23664 16544
rect 23716 16532 23722 16584
rect 21818 16464 21824 16516
rect 21876 16504 21882 16516
rect 21876 16476 21942 16504
rect 21876 16464 21882 16476
rect 22830 16464 22836 16516
rect 22888 16504 22894 16516
rect 23768 16504 23796 16612
rect 25240 16584 25268 16612
rect 25314 16600 25320 16652
rect 25372 16640 25378 16652
rect 25685 16643 25743 16649
rect 25685 16640 25697 16643
rect 25372 16612 25697 16640
rect 25372 16600 25378 16612
rect 25685 16609 25697 16612
rect 25731 16609 25743 16643
rect 25685 16603 25743 16609
rect 25774 16600 25780 16652
rect 25832 16640 25838 16652
rect 25869 16643 25927 16649
rect 25869 16640 25881 16643
rect 25832 16612 25881 16640
rect 25832 16600 25838 16612
rect 25869 16609 25881 16612
rect 25915 16609 25927 16643
rect 26050 16640 26056 16652
rect 26011 16612 26056 16640
rect 25869 16603 25927 16609
rect 26050 16600 26056 16612
rect 26108 16600 26114 16652
rect 26142 16600 26148 16652
rect 26200 16640 26206 16652
rect 26697 16643 26755 16649
rect 26200 16612 26245 16640
rect 26200 16600 26206 16612
rect 26697 16609 26709 16643
rect 26743 16640 26755 16643
rect 26970 16640 26976 16652
rect 26743 16612 26976 16640
rect 26743 16609 26755 16612
rect 26697 16603 26755 16609
rect 26970 16600 26976 16612
rect 27028 16600 27034 16652
rect 27264 16649 27292 16680
rect 28258 16668 28264 16680
rect 28316 16668 28322 16720
rect 31220 16708 31248 16748
rect 31294 16736 31300 16748
rect 31352 16736 31358 16788
rect 28748 16680 31248 16708
rect 27249 16643 27307 16649
rect 27249 16609 27261 16643
rect 27295 16609 27307 16643
rect 27249 16603 27307 16609
rect 27430 16600 27436 16652
rect 27488 16640 27494 16652
rect 28748 16640 28776 16680
rect 27488 16612 28776 16640
rect 29012 16612 30144 16640
rect 27488 16600 27494 16612
rect 29012 16584 29040 16612
rect 24854 16582 24860 16584
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16541 23903 16575
rect 24780 16572 24860 16582
rect 24767 16544 24860 16572
rect 23845 16535 23903 16541
rect 22888 16476 23796 16504
rect 22888 16464 22894 16476
rect 23860 16436 23888 16535
rect 24486 16464 24492 16516
rect 24544 16504 24550 16516
rect 24780 16504 24808 16544
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 24544 16476 24808 16504
rect 24964 16504 24992 16535
rect 25038 16532 25044 16584
rect 25096 16572 25102 16584
rect 25096 16544 25141 16572
rect 25096 16532 25102 16544
rect 25222 16532 25228 16584
rect 25280 16572 25286 16584
rect 25958 16572 25964 16584
rect 25280 16544 25325 16572
rect 25919 16544 25964 16572
rect 25280 16532 25286 16544
rect 25958 16532 25964 16544
rect 26016 16532 26022 16584
rect 26602 16532 26608 16584
rect 26660 16572 26666 16584
rect 27065 16575 27123 16581
rect 27065 16572 27077 16575
rect 26660 16544 27077 16572
rect 26660 16532 26666 16544
rect 27065 16541 27077 16544
rect 27111 16572 27123 16575
rect 27706 16572 27712 16584
rect 27111 16544 27712 16572
rect 27111 16541 27123 16544
rect 27065 16535 27123 16541
rect 27706 16532 27712 16544
rect 27764 16532 27770 16584
rect 28169 16575 28227 16581
rect 28169 16541 28181 16575
rect 28215 16541 28227 16575
rect 28994 16572 29000 16584
rect 28955 16544 29000 16572
rect 28169 16535 28227 16541
rect 24964 16476 25268 16504
rect 24544 16464 24550 16476
rect 21744 16408 23888 16436
rect 21637 16399 21695 16405
rect 24026 16396 24032 16448
rect 24084 16436 24090 16448
rect 24581 16439 24639 16445
rect 24581 16436 24593 16439
rect 24084 16408 24593 16436
rect 24084 16396 24090 16408
rect 24581 16405 24593 16408
rect 24627 16405 24639 16439
rect 25240 16436 25268 16476
rect 25314 16464 25320 16516
rect 25372 16504 25378 16516
rect 27893 16507 27951 16513
rect 27893 16504 27905 16507
rect 25372 16476 27905 16504
rect 25372 16464 25378 16476
rect 27893 16473 27905 16476
rect 27939 16473 27951 16507
rect 27893 16467 27951 16473
rect 26878 16436 26884 16448
rect 25240 16408 26884 16436
rect 24581 16399 24639 16405
rect 26878 16396 26884 16408
rect 26936 16396 26942 16448
rect 27062 16436 27068 16448
rect 27023 16408 27068 16436
rect 27062 16396 27068 16408
rect 27120 16396 27126 16448
rect 27430 16396 27436 16448
rect 27488 16436 27494 16448
rect 28184 16436 28212 16535
rect 28994 16532 29000 16544
rect 29052 16532 29058 16584
rect 29089 16575 29147 16581
rect 29089 16541 29101 16575
rect 29135 16572 29147 16575
rect 29178 16572 29184 16584
rect 29135 16544 29184 16572
rect 29135 16541 29147 16544
rect 29089 16535 29147 16541
rect 29178 16532 29184 16544
rect 29236 16532 29242 16584
rect 28810 16464 28816 16516
rect 28868 16504 28874 16516
rect 30116 16513 30144 16612
rect 30650 16532 30656 16584
rect 30708 16532 30714 16584
rect 29885 16507 29943 16513
rect 29885 16504 29897 16507
rect 28868 16476 29897 16504
rect 28868 16464 28874 16476
rect 29885 16473 29897 16476
rect 29931 16473 29943 16507
rect 29885 16467 29943 16473
rect 30101 16507 30159 16513
rect 30101 16473 30113 16507
rect 30147 16473 30159 16507
rect 30668 16504 30696 16532
rect 30101 16467 30159 16473
rect 30392 16476 30696 16504
rect 30745 16507 30803 16513
rect 30392 16448 30420 16476
rect 30745 16473 30757 16507
rect 30791 16504 30803 16507
rect 31294 16504 31300 16516
rect 30791 16476 31300 16504
rect 30791 16473 30803 16476
rect 30745 16467 30803 16473
rect 31294 16464 31300 16476
rect 31352 16464 31358 16516
rect 28442 16436 28448 16448
rect 27488 16408 28448 16436
rect 27488 16396 27494 16408
rect 28442 16396 28448 16408
rect 28500 16396 28506 16448
rect 28721 16439 28779 16445
rect 28721 16405 28733 16439
rect 28767 16436 28779 16439
rect 29638 16436 29644 16448
rect 28767 16408 29644 16436
rect 28767 16405 28779 16408
rect 28721 16399 28779 16405
rect 29638 16396 29644 16408
rect 29696 16396 29702 16448
rect 29730 16396 29736 16448
rect 29788 16436 29794 16448
rect 29788 16408 29833 16436
rect 29788 16396 29794 16408
rect 30374 16396 30380 16448
rect 30432 16396 30438 16448
rect 30650 16436 30656 16448
rect 30611 16408 30656 16436
rect 30650 16396 30656 16408
rect 30708 16396 30714 16448
rect 1104 16346 31992 16368
rect 1104 16294 8632 16346
rect 8684 16294 8696 16346
rect 8748 16294 8760 16346
rect 8812 16294 8824 16346
rect 8876 16294 8888 16346
rect 8940 16294 16314 16346
rect 16366 16294 16378 16346
rect 16430 16294 16442 16346
rect 16494 16294 16506 16346
rect 16558 16294 16570 16346
rect 16622 16294 23996 16346
rect 24048 16294 24060 16346
rect 24112 16294 24124 16346
rect 24176 16294 24188 16346
rect 24240 16294 24252 16346
rect 24304 16294 31678 16346
rect 31730 16294 31742 16346
rect 31794 16294 31806 16346
rect 31858 16294 31870 16346
rect 31922 16294 31934 16346
rect 31986 16294 31992 16346
rect 1104 16272 31992 16294
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10928 16204 11069 16232
rect 10928 16192 10934 16204
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 11057 16195 11115 16201
rect 12161 16235 12219 16241
rect 12161 16201 12173 16235
rect 12207 16232 12219 16235
rect 12342 16232 12348 16244
rect 12207 16204 12348 16232
rect 12207 16201 12219 16204
rect 12161 16195 12219 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 14182 16192 14188 16244
rect 14240 16232 14246 16244
rect 14734 16232 14740 16244
rect 14240 16204 14740 16232
rect 14240 16192 14246 16204
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 15010 16192 15016 16244
rect 15068 16232 15074 16244
rect 16301 16235 16359 16241
rect 16301 16232 16313 16235
rect 15068 16204 16313 16232
rect 15068 16192 15074 16204
rect 16301 16201 16313 16204
rect 16347 16201 16359 16235
rect 16301 16195 16359 16201
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 16850 16232 16856 16244
rect 16448 16204 16856 16232
rect 16448 16192 16454 16204
rect 16850 16192 16856 16204
rect 16908 16192 16914 16244
rect 17862 16232 17868 16244
rect 16960 16204 17868 16232
rect 10597 16167 10655 16173
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 11238 16164 11244 16176
rect 10643 16136 11244 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 12713 16167 12771 16173
rect 12713 16133 12725 16167
rect 12759 16164 12771 16167
rect 16758 16164 16764 16176
rect 12759 16136 16764 16164
rect 12759 16133 12771 16136
rect 12713 16127 12771 16133
rect 16758 16124 16764 16136
rect 16816 16124 16822 16176
rect 16960 16173 16988 16204
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18138 16232 18144 16244
rect 17972 16204 18144 16232
rect 16945 16167 17003 16173
rect 16945 16133 16957 16167
rect 16991 16133 17003 16167
rect 17972 16164 18000 16204
rect 18138 16192 18144 16204
rect 18196 16232 18202 16244
rect 18874 16232 18880 16244
rect 18196 16204 18880 16232
rect 18196 16192 18202 16204
rect 18874 16192 18880 16204
rect 18932 16192 18938 16244
rect 19150 16192 19156 16244
rect 19208 16232 19214 16244
rect 20530 16232 20536 16244
rect 19208 16204 20392 16232
rect 20491 16204 20536 16232
rect 19208 16192 19214 16204
rect 16945 16127 17003 16133
rect 17604 16136 18000 16164
rect 11330 16056 11336 16108
rect 11388 16096 11394 16108
rect 12621 16099 12679 16105
rect 12621 16096 12633 16099
rect 11388 16068 12633 16096
rect 11388 16056 11394 16068
rect 12621 16065 12633 16068
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 13044 16068 13277 16096
rect 13044 16056 13050 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13449 16099 13507 16105
rect 13449 16096 13461 16099
rect 13412 16068 13461 16096
rect 13412 16056 13418 16068
rect 13449 16065 13461 16068
rect 13495 16096 13507 16099
rect 13814 16096 13820 16108
rect 13495 16068 13820 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14185 16099 14243 16105
rect 13964 16068 14009 16096
rect 13964 16056 13970 16068
rect 14185 16065 14197 16099
rect 14231 16096 14243 16099
rect 14550 16096 14556 16108
rect 14231 16068 14556 16096
rect 14231 16065 14243 16068
rect 14185 16059 14243 16065
rect 14550 16056 14556 16068
rect 14608 16096 14614 16108
rect 14829 16099 14887 16105
rect 14829 16096 14841 16099
rect 14608 16068 14841 16096
rect 14608 16056 14614 16068
rect 14829 16065 14841 16068
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15194 16096 15200 16108
rect 15059 16068 15200 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 14936 16028 14964 16059
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 16025 16099 16083 16105
rect 16025 16096 16037 16099
rect 15804 16068 16037 16096
rect 15804 16056 15810 16068
rect 16025 16065 16037 16068
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 16142 16099 16200 16105
rect 16142 16065 16154 16099
rect 16188 16096 16200 16099
rect 17604 16096 17632 16136
rect 19058 16124 19064 16176
rect 19116 16164 19122 16176
rect 19116 16136 19550 16164
rect 19116 16124 19122 16136
rect 17770 16096 17776 16108
rect 16188 16068 16896 16096
rect 16188 16065 16200 16068
rect 16142 16059 16200 16065
rect 15286 16028 15292 16040
rect 14936 16000 15292 16028
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 15654 16028 15660 16040
rect 15615 16000 15660 16028
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 15838 15988 15844 16040
rect 15896 16028 15902 16040
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15896 16000 15945 16028
rect 15896 15988 15902 16000
rect 15933 15997 15945 16000
rect 15979 15997 15991 16031
rect 16040 16028 16068 16059
rect 16666 16028 16672 16040
rect 16040 16000 16672 16028
rect 15933 15991 15991 15997
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 16868 16028 16896 16068
rect 16960 16068 17632 16096
rect 17731 16068 17776 16096
rect 16960 16028 16988 16068
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 18046 16056 18052 16108
rect 18104 16096 18110 16108
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 18104 16068 18153 16096
rect 18104 16056 18110 16068
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 18233 16099 18291 16105
rect 18233 16065 18245 16099
rect 18279 16096 18291 16099
rect 18322 16096 18328 16108
rect 18279 16068 18328 16096
rect 18279 16065 18291 16068
rect 18233 16059 18291 16065
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 20364 16096 20392 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 23290 16192 23296 16244
rect 23348 16232 23354 16244
rect 23753 16235 23811 16241
rect 23348 16204 23612 16232
rect 23348 16192 23354 16204
rect 20622 16124 20628 16176
rect 20680 16164 20686 16176
rect 21453 16167 21511 16173
rect 21453 16164 21465 16167
rect 20680 16136 21465 16164
rect 20680 16124 20686 16136
rect 21453 16133 21465 16136
rect 21499 16133 21511 16167
rect 22278 16164 22284 16176
rect 22239 16136 22284 16164
rect 21453 16127 21511 16133
rect 22278 16124 22284 16136
rect 22336 16124 22342 16176
rect 22554 16124 22560 16176
rect 22612 16164 22618 16176
rect 22612 16136 22770 16164
rect 22612 16124 22618 16136
rect 20993 16099 21051 16105
rect 20993 16096 21005 16099
rect 20364 16068 21005 16096
rect 20993 16065 21005 16068
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 16868 16000 16988 16028
rect 17126 15988 17132 16040
rect 17184 16028 17190 16040
rect 18690 16028 18696 16040
rect 17184 16000 18696 16028
rect 17184 15988 17190 16000
rect 18690 15988 18696 16000
rect 18748 16028 18754 16040
rect 18785 16031 18843 16037
rect 18785 16028 18797 16031
rect 18748 16000 18797 16028
rect 18748 15988 18754 16000
rect 18785 15997 18797 16000
rect 18831 15997 18843 16031
rect 19058 16028 19064 16040
rect 19019 16000 19064 16028
rect 18785 15991 18843 15997
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 19150 15988 19156 16040
rect 19208 16028 19214 16040
rect 20254 16028 20260 16040
rect 19208 16000 20260 16028
rect 19208 15988 19214 16000
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 21100 16028 21128 16059
rect 21174 16056 21180 16108
rect 21232 16096 21238 16108
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 21232 16068 21281 16096
rect 21232 16056 21238 16068
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 21269 16059 21327 16065
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 23584 16096 23612 16204
rect 23753 16201 23765 16235
rect 23799 16201 23811 16235
rect 23753 16195 23811 16201
rect 23768 16164 23796 16195
rect 24026 16192 24032 16244
rect 24084 16232 24090 16244
rect 24854 16232 24860 16244
rect 24084 16204 24860 16232
rect 24084 16192 24090 16204
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 26050 16192 26056 16244
rect 26108 16232 26114 16244
rect 28261 16235 28319 16241
rect 28261 16232 28273 16235
rect 26108 16204 28273 16232
rect 26108 16192 26114 16204
rect 28261 16201 28273 16204
rect 28307 16201 28319 16235
rect 28261 16195 28319 16201
rect 28350 16192 28356 16244
rect 28408 16232 28414 16244
rect 29273 16235 29331 16241
rect 29273 16232 29285 16235
rect 28408 16204 29285 16232
rect 28408 16192 28414 16204
rect 29273 16201 29285 16204
rect 29319 16232 29331 16235
rect 29914 16232 29920 16244
rect 29319 16204 29920 16232
rect 29319 16201 29331 16204
rect 29273 16195 29331 16201
rect 29914 16192 29920 16204
rect 29972 16192 29978 16244
rect 30098 16192 30104 16244
rect 30156 16232 30162 16244
rect 31205 16235 31263 16241
rect 31205 16232 31217 16235
rect 30156 16204 31217 16232
rect 30156 16192 30162 16204
rect 31205 16201 31217 16204
rect 31251 16201 31263 16235
rect 31205 16195 31263 16201
rect 31294 16192 31300 16244
rect 31352 16232 31358 16244
rect 31662 16232 31668 16244
rect 31352 16204 31668 16232
rect 31352 16192 31358 16204
rect 31662 16192 31668 16204
rect 31720 16192 31726 16244
rect 23934 16164 23940 16176
rect 23768 16136 23940 16164
rect 23934 16124 23940 16136
rect 23992 16124 23998 16176
rect 24489 16167 24547 16173
rect 24489 16164 24501 16167
rect 24044 16136 24501 16164
rect 24044 16096 24072 16136
rect 24489 16133 24501 16136
rect 24535 16133 24547 16167
rect 24489 16127 24547 16133
rect 25038 16124 25044 16176
rect 25096 16124 25102 16176
rect 26142 16124 26148 16176
rect 26200 16164 26206 16176
rect 26200 16136 27844 16164
rect 26200 16124 26206 16136
rect 23584 16068 24072 16096
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 21008 16000 21128 16028
rect 21361 16031 21419 16037
rect 14090 15960 14096 15972
rect 14051 15932 14096 15960
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 14182 15920 14188 15972
rect 14240 15960 14246 15972
rect 15197 15963 15255 15969
rect 14240 15932 14285 15960
rect 14240 15920 14246 15932
rect 15197 15929 15209 15963
rect 15243 15960 15255 15963
rect 15378 15960 15384 15972
rect 15243 15932 15384 15960
rect 15243 15929 15255 15932
rect 15197 15923 15255 15929
rect 15378 15920 15384 15932
rect 15436 15920 15442 15972
rect 15488 15960 15516 15988
rect 16206 15960 16212 15972
rect 15488 15932 16212 15960
rect 16206 15920 16212 15932
rect 16264 15920 16270 15972
rect 16574 15920 16580 15972
rect 16632 15960 16638 15972
rect 16632 15932 17356 15960
rect 16632 15920 16638 15932
rect 13354 15892 13360 15904
rect 13315 15864 13360 15892
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14645 15895 14703 15901
rect 14645 15861 14657 15895
rect 14691 15892 14703 15895
rect 15470 15892 15476 15904
rect 14691 15864 15476 15892
rect 14691 15861 14703 15864
rect 14645 15855 14703 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 15838 15852 15844 15904
rect 15896 15892 15902 15904
rect 16114 15892 16120 15904
rect 15896 15864 16120 15892
rect 15896 15852 15902 15864
rect 16114 15852 16120 15864
rect 16172 15892 16178 15904
rect 16666 15892 16672 15904
rect 16172 15864 16672 15892
rect 16172 15852 16178 15864
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17218 15892 17224 15904
rect 16908 15864 17224 15892
rect 16908 15852 16914 15864
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 17328 15892 17356 15932
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 17589 15963 17647 15969
rect 17589 15960 17601 15963
rect 17552 15932 17601 15960
rect 17552 15920 17558 15932
rect 17589 15929 17601 15932
rect 17635 15929 17647 15963
rect 17589 15923 17647 15929
rect 18322 15920 18328 15972
rect 18380 15960 18386 15972
rect 21008 15960 21036 16000
rect 21361 15997 21373 16031
rect 21407 16028 21419 16031
rect 21542 16028 21548 16040
rect 21407 16000 21548 16028
rect 21407 15997 21419 16000
rect 21361 15991 21419 15997
rect 21542 15988 21548 16000
rect 21600 15988 21606 16040
rect 22370 15988 22376 16040
rect 22428 16028 22434 16040
rect 23750 16028 23756 16040
rect 22428 16000 23756 16028
rect 22428 15988 22434 16000
rect 23750 15988 23756 16000
rect 23808 16028 23814 16040
rect 24213 16031 24271 16037
rect 24213 16028 24225 16031
rect 23808 16000 24225 16028
rect 23808 15988 23814 16000
rect 24213 15997 24225 16000
rect 24259 15997 24271 16031
rect 26436 16028 26464 16059
rect 26510 16056 26516 16108
rect 26568 16096 26574 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 26568 16068 27169 16096
rect 26568 16056 26574 16068
rect 27157 16065 27169 16068
rect 27203 16096 27215 16099
rect 27430 16096 27436 16108
rect 27203 16068 27436 16096
rect 27203 16065 27215 16068
rect 27157 16059 27215 16065
rect 27430 16056 27436 16068
rect 27488 16056 27494 16108
rect 27816 16094 27844 16136
rect 27890 16124 27896 16176
rect 27948 16164 27954 16176
rect 29638 16164 29644 16176
rect 27948 16136 28212 16164
rect 27948 16124 27954 16136
rect 28184 16105 28212 16136
rect 28828 16136 29644 16164
rect 28077 16099 28135 16105
rect 28077 16096 28089 16099
rect 27934 16094 28089 16096
rect 27816 16068 28089 16094
rect 27816 16066 27962 16068
rect 28077 16065 28089 16068
rect 28123 16065 28135 16099
rect 28077 16059 28135 16065
rect 28169 16099 28227 16105
rect 28169 16065 28181 16099
rect 28215 16065 28227 16099
rect 28169 16059 28227 16065
rect 24213 15991 24271 15997
rect 24320 16000 26464 16028
rect 18380 15932 18644 15960
rect 18380 15920 18386 15932
rect 17678 15892 17684 15904
rect 17328 15864 17684 15892
rect 17678 15852 17684 15864
rect 17736 15852 17742 15904
rect 17865 15895 17923 15901
rect 17865 15861 17877 15895
rect 17911 15892 17923 15895
rect 18506 15892 18512 15904
rect 17911 15864 18512 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 18616 15892 18644 15932
rect 20180 15932 21036 15960
rect 20180 15892 20208 15932
rect 23382 15920 23388 15972
rect 23440 15960 23446 15972
rect 23566 15960 23572 15972
rect 23440 15932 23572 15960
rect 23440 15920 23446 15932
rect 23566 15920 23572 15932
rect 23624 15920 23630 15972
rect 23658 15920 23664 15972
rect 23716 15960 23722 15972
rect 24320 15960 24348 16000
rect 26602 15988 26608 16040
rect 26660 16028 26666 16040
rect 27341 16031 27399 16037
rect 27341 16028 27353 16031
rect 26660 16000 27353 16028
rect 26660 15988 26666 16000
rect 27341 15997 27353 16000
rect 27387 15997 27399 16031
rect 28445 16031 28503 16037
rect 28445 16028 28457 16031
rect 27341 15991 27399 15997
rect 28000 16000 28457 16028
rect 26513 15963 26571 15969
rect 26513 15960 26525 15963
rect 23716 15932 24348 15960
rect 25516 15932 26525 15960
rect 23716 15920 23722 15932
rect 18616 15864 20208 15892
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 25516 15892 25544 15932
rect 26513 15929 26525 15932
rect 26559 15929 26571 15963
rect 26513 15923 26571 15929
rect 27062 15920 27068 15972
rect 27120 15960 27126 15972
rect 27890 15960 27896 15972
rect 27120 15932 27896 15960
rect 27120 15920 27126 15932
rect 27890 15920 27896 15932
rect 27948 15920 27954 15972
rect 20312 15864 25544 15892
rect 20312 15852 20318 15864
rect 25590 15852 25596 15904
rect 25648 15892 25654 15904
rect 25961 15895 26019 15901
rect 25961 15892 25973 15895
rect 25648 15864 25973 15892
rect 25648 15852 25654 15864
rect 25961 15861 25973 15864
rect 26007 15861 26019 15895
rect 25961 15855 26019 15861
rect 26234 15852 26240 15904
rect 26292 15892 26298 15904
rect 28000 15892 28028 16000
rect 28445 15997 28457 16000
rect 28491 15997 28503 16031
rect 28445 15991 28503 15997
rect 28074 15920 28080 15972
rect 28132 15960 28138 15972
rect 28169 15963 28227 15969
rect 28169 15960 28181 15963
rect 28132 15932 28181 15960
rect 28132 15920 28138 15932
rect 28169 15929 28181 15932
rect 28215 15929 28227 15963
rect 28169 15923 28227 15929
rect 26292 15864 28028 15892
rect 28828 15892 28856 16136
rect 29638 16124 29644 16136
rect 29696 16164 29702 16176
rect 30009 16167 30067 16173
rect 30009 16164 30021 16167
rect 29696 16136 30021 16164
rect 29696 16124 29702 16136
rect 30009 16133 30021 16136
rect 30055 16133 30067 16167
rect 30009 16127 30067 16133
rect 30561 16167 30619 16173
rect 30561 16133 30573 16167
rect 30607 16164 30619 16167
rect 30742 16164 30748 16176
rect 30607 16136 30748 16164
rect 30607 16133 30619 16136
rect 30561 16127 30619 16133
rect 30742 16124 30748 16136
rect 30800 16124 30806 16176
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16096 29147 16099
rect 29178 16096 29184 16108
rect 29135 16068 29184 16096
rect 29135 16065 29147 16068
rect 29089 16059 29147 16065
rect 29178 16056 29184 16068
rect 29236 16056 29242 16108
rect 29270 16056 29276 16108
rect 29328 16096 29334 16108
rect 29733 16099 29791 16105
rect 29733 16096 29745 16099
rect 29328 16068 29745 16096
rect 29328 16056 29334 16068
rect 29733 16065 29745 16068
rect 29779 16065 29791 16099
rect 29733 16059 29791 16065
rect 29825 16099 29883 16105
rect 29825 16065 29837 16099
rect 29871 16096 29883 16099
rect 29914 16096 29920 16108
rect 29871 16068 29920 16096
rect 29871 16065 29883 16068
rect 29825 16059 29883 16065
rect 28905 16031 28963 16037
rect 28905 15997 28917 16031
rect 28951 15997 28963 16031
rect 28905 15991 28963 15997
rect 28920 15960 28948 15991
rect 29362 15988 29368 16040
rect 29420 15988 29426 16040
rect 29748 16028 29776 16059
rect 29914 16056 29920 16068
rect 29972 16056 29978 16108
rect 30190 16028 30196 16040
rect 29748 16000 30196 16028
rect 30190 15988 30196 16000
rect 30248 15988 30254 16040
rect 29380 15960 29408 15988
rect 28920 15932 29408 15960
rect 29638 15920 29644 15972
rect 29696 15960 29702 15972
rect 30742 15960 30748 15972
rect 29696 15932 30748 15960
rect 29696 15920 29702 15932
rect 30742 15920 30748 15932
rect 30800 15920 30806 15972
rect 29086 15892 29092 15904
rect 28828 15864 29092 15892
rect 26292 15852 26298 15864
rect 29086 15852 29092 15864
rect 29144 15852 29150 15904
rect 29362 15852 29368 15904
rect 29420 15892 29426 15904
rect 29733 15895 29791 15901
rect 29733 15892 29745 15895
rect 29420 15864 29745 15892
rect 29420 15852 29426 15864
rect 29733 15861 29745 15864
rect 29779 15861 29791 15895
rect 29733 15855 29791 15861
rect 1104 15802 31832 15824
rect 1104 15750 4791 15802
rect 4843 15750 4855 15802
rect 4907 15750 4919 15802
rect 4971 15750 4983 15802
rect 5035 15750 5047 15802
rect 5099 15750 12473 15802
rect 12525 15750 12537 15802
rect 12589 15750 12601 15802
rect 12653 15750 12665 15802
rect 12717 15750 12729 15802
rect 12781 15750 20155 15802
rect 20207 15750 20219 15802
rect 20271 15750 20283 15802
rect 20335 15750 20347 15802
rect 20399 15750 20411 15802
rect 20463 15750 27837 15802
rect 27889 15750 27901 15802
rect 27953 15750 27965 15802
rect 28017 15750 28029 15802
rect 28081 15750 28093 15802
rect 28145 15750 31832 15802
rect 1104 15728 31832 15750
rect 11330 15688 11336 15700
rect 11291 15660 11336 15688
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 11790 15688 11796 15700
rect 11751 15660 11796 15688
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 14829 15691 14887 15697
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 14918 15688 14924 15700
rect 14875 15660 14924 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 15160 15660 15301 15688
rect 15160 15648 15166 15660
rect 15289 15657 15301 15660
rect 15335 15657 15347 15691
rect 15289 15651 15347 15657
rect 15473 15691 15531 15697
rect 15473 15657 15485 15691
rect 15519 15688 15531 15691
rect 15838 15688 15844 15700
rect 15519 15660 15844 15688
rect 15519 15657 15531 15660
rect 15473 15651 15531 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 15930 15648 15936 15700
rect 15988 15688 15994 15700
rect 16298 15688 16304 15700
rect 15988 15660 16304 15688
rect 15988 15648 15994 15660
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16482 15688 16488 15700
rect 16443 15660 16488 15688
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 16669 15691 16727 15697
rect 16669 15657 16681 15691
rect 16715 15688 16727 15691
rect 16715 15660 16794 15688
rect 16715 15657 16727 15660
rect 16669 15651 16727 15657
rect 11238 15580 11244 15632
rect 11296 15620 11302 15632
rect 12345 15623 12403 15629
rect 12345 15620 12357 15623
rect 11296 15592 12357 15620
rect 11296 15580 11302 15592
rect 12345 15589 12357 15592
rect 12391 15589 12403 15623
rect 12345 15583 12403 15589
rect 13633 15623 13691 15629
rect 13633 15589 13645 15623
rect 13679 15620 13691 15623
rect 15562 15620 15568 15632
rect 13679 15592 15568 15620
rect 13679 15589 13691 15592
rect 13633 15583 13691 15589
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 16114 15620 16120 15632
rect 15660 15592 16120 15620
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 15660 15552 15688 15592
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 16766 15620 16794 15660
rect 17034 15648 17040 15700
rect 17092 15688 17098 15700
rect 17092 15660 18825 15688
rect 17092 15648 17098 15660
rect 17586 15620 17592 15632
rect 16766 15592 17592 15620
rect 17586 15580 17592 15592
rect 17644 15580 17650 15632
rect 18797 15620 18825 15660
rect 18966 15648 18972 15700
rect 19024 15688 19030 15700
rect 19024 15660 20760 15688
rect 19024 15648 19030 15660
rect 19150 15620 19156 15632
rect 18797 15592 19156 15620
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 19426 15580 19432 15632
rect 19484 15580 19490 15632
rect 13136 15524 13584 15552
rect 13136 15512 13142 15524
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 11790 15444 11796 15496
rect 11848 15484 11854 15496
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 11848 15456 12909 15484
rect 11848 15444 11854 15456
rect 12897 15453 12909 15456
rect 12943 15484 12955 15487
rect 13262 15484 13268 15496
rect 12943 15456 13268 15484
rect 12943 15453 12955 15456
rect 12897 15447 12955 15453
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 13556 15493 13584 15524
rect 14752 15524 15688 15552
rect 14752 15493 14780 15524
rect 15930 15512 15936 15564
rect 15988 15552 15994 15564
rect 16393 15555 16451 15561
rect 16393 15552 16405 15555
rect 15988 15524 16405 15552
rect 15988 15512 15994 15524
rect 16393 15521 16405 15524
rect 16439 15521 16451 15555
rect 16393 15515 16451 15521
rect 16942 15512 16948 15564
rect 17000 15552 17006 15564
rect 19058 15552 19064 15564
rect 17000 15524 19064 15552
rect 17000 15512 17006 15524
rect 19058 15512 19064 15524
rect 19116 15512 19122 15564
rect 19444 15552 19472 15580
rect 20070 15552 20076 15564
rect 19444 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 20732 15552 20760 15660
rect 20898 15648 20904 15700
rect 20956 15688 20962 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20956 15660 21189 15688
rect 20956 15648 20962 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 21177 15651 21235 15657
rect 21450 15648 21456 15700
rect 21508 15688 21514 15700
rect 24670 15688 24676 15700
rect 21508 15660 24676 15688
rect 21508 15648 21514 15660
rect 24670 15648 24676 15660
rect 24728 15648 24734 15700
rect 25958 15648 25964 15700
rect 26016 15688 26022 15700
rect 27062 15688 27068 15700
rect 26016 15660 27068 15688
rect 26016 15648 26022 15660
rect 27062 15648 27068 15660
rect 27120 15648 27126 15700
rect 27890 15688 27896 15700
rect 27851 15660 27896 15688
rect 27890 15648 27896 15660
rect 27948 15648 27954 15700
rect 28077 15691 28135 15697
rect 28077 15688 28089 15691
rect 28000 15660 28089 15688
rect 23106 15580 23112 15632
rect 23164 15620 23170 15632
rect 23164 15592 23520 15620
rect 23164 15580 23170 15592
rect 21913 15555 21971 15561
rect 21913 15552 21925 15555
rect 20732 15524 21925 15552
rect 21913 15521 21925 15524
rect 21959 15521 21971 15555
rect 23492 15552 23520 15592
rect 23566 15580 23572 15632
rect 23624 15620 23630 15632
rect 23937 15623 23995 15629
rect 23937 15620 23949 15623
rect 23624 15592 23949 15620
rect 23624 15580 23630 15592
rect 23937 15589 23949 15592
rect 23983 15589 23995 15623
rect 23937 15583 23995 15589
rect 27430 15580 27436 15632
rect 27488 15620 27494 15632
rect 28000 15620 28028 15660
rect 28077 15657 28089 15660
rect 28123 15688 28135 15691
rect 28810 15688 28816 15700
rect 28123 15660 28816 15688
rect 28123 15657 28135 15660
rect 28077 15651 28135 15657
rect 28810 15648 28816 15660
rect 28868 15648 28874 15700
rect 28994 15648 29000 15700
rect 29052 15688 29058 15700
rect 30561 15691 30619 15697
rect 30561 15688 30573 15691
rect 29052 15660 30573 15688
rect 29052 15648 29058 15660
rect 30561 15657 30573 15660
rect 30607 15657 30619 15691
rect 30561 15651 30619 15657
rect 27488 15592 28028 15620
rect 27488 15580 27494 15592
rect 28258 15580 28264 15632
rect 28316 15620 28322 15632
rect 29086 15620 29092 15632
rect 28316 15592 29092 15620
rect 28316 15580 28322 15592
rect 29086 15580 29092 15592
rect 29144 15580 29150 15632
rect 29917 15623 29975 15629
rect 29917 15589 29929 15623
rect 29963 15620 29975 15623
rect 30190 15620 30196 15632
rect 29963 15592 30196 15620
rect 29963 15589 29975 15592
rect 29917 15583 29975 15589
rect 30190 15580 30196 15592
rect 30248 15580 30254 15632
rect 23492 15524 26004 15552
rect 21913 15515 21971 15521
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 10870 15376 10876 15428
rect 10928 15416 10934 15428
rect 13078 15416 13084 15428
rect 10928 15388 13084 15416
rect 10928 15376 10934 15388
rect 13078 15376 13084 15388
rect 13136 15376 13142 15428
rect 14553 15419 14611 15425
rect 14553 15385 14565 15419
rect 14599 15385 14611 15419
rect 14844 15416 14872 15447
rect 15010 15444 15016 15496
rect 15068 15484 15074 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15068 15456 16129 15484
rect 15068 15444 15074 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 16574 15484 16580 15496
rect 16264 15456 16580 15484
rect 16264 15444 16270 15456
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15484 18935 15487
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 18923 15456 19441 15484
rect 18923 15453 18935 15456
rect 18877 15447 18935 15453
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 21637 15487 21695 15493
rect 21637 15453 21649 15487
rect 21683 15453 21695 15487
rect 21637 15447 21695 15453
rect 15654 15416 15660 15428
rect 14844 15388 15660 15416
rect 14553 15379 14611 15385
rect 12986 15348 12992 15360
rect 12947 15320 12992 15348
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 14568 15348 14596 15379
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 16482 15376 16488 15428
rect 16540 15416 16546 15428
rect 16540 15388 17254 15416
rect 16540 15376 16546 15388
rect 15457 15351 15515 15357
rect 15457 15348 15469 15351
rect 14568 15320 15469 15348
rect 15457 15317 15469 15320
rect 15503 15348 15515 15351
rect 15562 15348 15568 15360
rect 15503 15320 15568 15348
rect 15503 15317 15515 15320
rect 15457 15311 15515 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 15672 15348 15700 15376
rect 17126 15348 17132 15360
rect 15672 15320 17132 15348
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 17226 15348 17254 15388
rect 17586 15376 17592 15428
rect 17644 15376 17650 15428
rect 18601 15419 18659 15425
rect 18601 15385 18613 15419
rect 18647 15385 18659 15419
rect 18601 15379 18659 15385
rect 17862 15348 17868 15360
rect 17226 15320 17868 15348
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18616 15348 18644 15379
rect 18690 15376 18696 15428
rect 18748 15416 18754 15428
rect 18892 15416 18920 15447
rect 18748 15388 18920 15416
rect 19444 15416 19472 15447
rect 19610 15416 19616 15428
rect 19444 15388 19616 15416
rect 18748 15376 18754 15388
rect 19610 15376 19616 15388
rect 19668 15376 19674 15428
rect 19702 15376 19708 15428
rect 19760 15416 19766 15428
rect 19760 15388 19805 15416
rect 19760 15376 19766 15388
rect 20714 15376 20720 15428
rect 20772 15376 20778 15428
rect 21652 15416 21680 15447
rect 23750 15444 23756 15496
rect 23808 15484 23814 15496
rect 23845 15487 23903 15493
rect 23845 15484 23857 15487
rect 23808 15456 23857 15484
rect 23808 15444 23814 15456
rect 23845 15453 23857 15456
rect 23891 15453 23903 15487
rect 23845 15447 23903 15453
rect 24486 15444 24492 15496
rect 24544 15484 24550 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24544 15456 24593 15484
rect 24544 15444 24550 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 25976 15470 26004 15524
rect 26786 15512 26792 15564
rect 26844 15552 26850 15564
rect 26844 15524 27200 15552
rect 26844 15512 26850 15524
rect 24581 15447 24639 15453
rect 26878 15444 26884 15496
rect 26936 15484 26942 15496
rect 27172 15493 27200 15524
rect 27522 15512 27528 15564
rect 27580 15552 27586 15564
rect 28537 15555 28595 15561
rect 27580 15524 28396 15552
rect 27580 15512 27586 15524
rect 26973 15487 27031 15493
rect 26973 15484 26985 15487
rect 26936 15456 26985 15484
rect 26936 15444 26942 15456
rect 26973 15453 26985 15456
rect 27019 15453 27031 15487
rect 26973 15447 27031 15453
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15453 27215 15487
rect 27157 15447 27215 15453
rect 27249 15487 27307 15493
rect 27249 15453 27261 15487
rect 27295 15484 27307 15487
rect 28258 15484 28264 15496
rect 27295 15456 28264 15484
rect 27295 15453 27307 15456
rect 27249 15447 27307 15453
rect 28258 15444 28264 15456
rect 28316 15444 28322 15496
rect 28368 15428 28396 15524
rect 28537 15521 28549 15555
rect 28583 15552 28595 15555
rect 28626 15552 28632 15564
rect 28583 15524 28632 15552
rect 28583 15521 28595 15524
rect 28537 15515 28595 15521
rect 28626 15512 28632 15524
rect 28684 15512 28690 15564
rect 29454 15444 29460 15496
rect 29512 15484 29518 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29512 15456 29745 15484
rect 29512 15444 29518 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 22002 15416 22008 15428
rect 21652 15388 22008 15416
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 24857 15419 24915 15425
rect 24857 15416 24869 15419
rect 22244 15388 22402 15416
rect 23308 15388 24869 15416
rect 22244 15376 22250 15388
rect 18874 15348 18880 15360
rect 18616 15320 18880 15348
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 23308 15348 23336 15388
rect 24857 15385 24869 15388
rect 24903 15385 24915 15419
rect 24857 15379 24915 15385
rect 27709 15419 27767 15425
rect 27709 15385 27721 15419
rect 27755 15416 27767 15419
rect 27798 15416 27804 15428
rect 27755 15388 27804 15416
rect 27755 15385 27767 15388
rect 27709 15379 27767 15385
rect 27798 15376 27804 15388
rect 27856 15376 27862 15428
rect 28350 15376 28356 15428
rect 28408 15416 28414 15428
rect 28721 15419 28779 15425
rect 28721 15416 28733 15419
rect 28408 15388 28733 15416
rect 28408 15376 28414 15388
rect 28721 15385 28733 15388
rect 28767 15385 28779 15419
rect 28721 15379 28779 15385
rect 28905 15419 28963 15425
rect 28905 15385 28917 15419
rect 28951 15416 28963 15419
rect 30466 15416 30472 15428
rect 28951 15388 30472 15416
rect 28951 15385 28963 15388
rect 28905 15379 28963 15385
rect 30466 15376 30472 15388
rect 30524 15376 30530 15428
rect 30650 15416 30656 15428
rect 30611 15388 30656 15416
rect 30650 15376 30656 15388
rect 30708 15376 30714 15428
rect 19484 15320 23336 15348
rect 23385 15351 23443 15357
rect 19484 15308 19490 15320
rect 23385 15317 23397 15351
rect 23431 15348 23443 15351
rect 26142 15348 26148 15360
rect 23431 15320 26148 15348
rect 23431 15317 23443 15320
rect 23385 15311 23443 15317
rect 26142 15308 26148 15320
rect 26200 15308 26206 15360
rect 26326 15348 26332 15360
rect 26287 15320 26332 15348
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 26786 15348 26792 15360
rect 26747 15320 26792 15348
rect 26786 15308 26792 15320
rect 26844 15308 26850 15360
rect 27919 15351 27977 15357
rect 27919 15317 27931 15351
rect 27965 15348 27977 15351
rect 28442 15348 28448 15360
rect 27965 15320 28448 15348
rect 27965 15317 27977 15320
rect 27919 15311 27977 15317
rect 28442 15308 28448 15320
rect 28500 15308 28506 15360
rect 28626 15308 28632 15360
rect 28684 15348 28690 15360
rect 29178 15348 29184 15360
rect 28684 15320 29184 15348
rect 28684 15308 28690 15320
rect 29178 15308 29184 15320
rect 29236 15308 29242 15360
rect 29914 15308 29920 15360
rect 29972 15348 29978 15360
rect 31205 15351 31263 15357
rect 31205 15348 31217 15351
rect 29972 15320 31217 15348
rect 29972 15308 29978 15320
rect 31205 15317 31217 15320
rect 31251 15348 31263 15351
rect 31662 15348 31668 15360
rect 31251 15320 31668 15348
rect 31251 15317 31263 15320
rect 31205 15311 31263 15317
rect 31662 15308 31668 15320
rect 31720 15308 31726 15360
rect 1104 15258 31992 15280
rect 1104 15206 8632 15258
rect 8684 15206 8696 15258
rect 8748 15206 8760 15258
rect 8812 15206 8824 15258
rect 8876 15206 8888 15258
rect 8940 15206 16314 15258
rect 16366 15206 16378 15258
rect 16430 15206 16442 15258
rect 16494 15206 16506 15258
rect 16558 15206 16570 15258
rect 16622 15206 23996 15258
rect 24048 15206 24060 15258
rect 24112 15206 24124 15258
rect 24176 15206 24188 15258
rect 24240 15206 24252 15258
rect 24304 15206 31678 15258
rect 31730 15206 31742 15258
rect 31794 15206 31806 15258
rect 31858 15206 31870 15258
rect 31922 15206 31934 15258
rect 31986 15206 31992 15258
rect 1104 15184 31992 15206
rect 11330 15104 11336 15156
rect 11388 15144 11394 15156
rect 11977 15147 12035 15153
rect 11977 15144 11989 15147
rect 11388 15116 11989 15144
rect 11388 15104 11394 15116
rect 11977 15113 11989 15116
rect 12023 15144 12035 15147
rect 12158 15144 12164 15156
rect 12023 15116 12164 15144
rect 12023 15113 12035 15116
rect 11977 15107 12035 15113
rect 12158 15104 12164 15116
rect 12216 15144 12222 15156
rect 12216 15116 14504 15144
rect 12216 15104 12222 15116
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 12989 15079 13047 15085
rect 12989 15076 13001 15079
rect 12400 15048 13001 15076
rect 12400 15036 12406 15048
rect 12989 15045 13001 15048
rect 13035 15076 13047 15079
rect 13906 15076 13912 15088
rect 13035 15048 13912 15076
rect 13035 15045 13047 15048
rect 12989 15039 13047 15045
rect 13906 15036 13912 15048
rect 13964 15036 13970 15088
rect 14476 15017 14504 15116
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15194 15144 15200 15156
rect 14792 15116 15200 15144
rect 14792 15104 14798 15116
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 15378 15104 15384 15156
rect 15436 15144 15442 15156
rect 17494 15144 17500 15156
rect 15436 15116 17500 15144
rect 15436 15104 15442 15116
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 18322 15104 18328 15156
rect 18380 15144 18386 15156
rect 18380 15116 20668 15144
rect 18380 15104 18386 15116
rect 15102 15076 15108 15088
rect 15063 15048 15108 15076
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 15712 15048 18722 15076
rect 15712 15036 15718 15048
rect 19794 15036 19800 15088
rect 19852 15076 19858 15088
rect 19852 15048 20208 15076
rect 19852 15036 19858 15048
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 14977 13875 15011
rect 13817 14971 13875 14977
rect 14461 15011 14519 15017
rect 14461 14977 14473 15011
rect 14507 14977 14519 15011
rect 15286 15008 15292 15020
rect 15247 14980 15292 15008
rect 14461 14971 14519 14977
rect 13832 14940 13860 14971
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15436 14980 15481 15008
rect 15436 14968 15442 14980
rect 15562 14968 15568 15020
rect 15620 15008 15626 15020
rect 16945 15011 17003 15017
rect 15620 14980 16344 15008
rect 15620 14968 15626 14980
rect 16316 14952 16344 14980
rect 16945 14977 16957 15011
rect 16991 15008 17003 15011
rect 17402 15008 17408 15020
rect 16991 14980 17408 15008
rect 16991 14977 17003 14980
rect 16945 14971 17003 14977
rect 17402 14968 17408 14980
rect 17460 14968 17466 15020
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 15008 17647 15011
rect 17862 15008 17868 15020
rect 17635 14980 17868 15008
rect 17635 14977 17647 14980
rect 17589 14971 17647 14977
rect 17862 14968 17868 14980
rect 17920 15008 17926 15020
rect 18598 15008 18604 15020
rect 17920 14980 18604 15008
rect 17920 14968 17926 14980
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 15841 14943 15899 14949
rect 15841 14940 15853 14943
rect 13832 14912 15853 14940
rect 15841 14909 15853 14912
rect 15887 14909 15899 14943
rect 16114 14940 16120 14952
rect 15841 14903 15899 14909
rect 15948 14912 16120 14940
rect 14553 14875 14611 14881
rect 14553 14841 14565 14875
rect 14599 14872 14611 14875
rect 14918 14872 14924 14884
rect 14599 14844 14924 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 15194 14832 15200 14884
rect 15252 14872 15258 14884
rect 15948 14872 15976 14912
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 16298 14940 16304 14952
rect 16259 14912 16304 14940
rect 16298 14900 16304 14912
rect 16356 14900 16362 14952
rect 16482 14900 16488 14952
rect 16540 14940 16546 14952
rect 17678 14940 17684 14952
rect 16540 14912 17540 14940
rect 17639 14912 17684 14940
rect 16540 14900 16546 14912
rect 15252 14844 15976 14872
rect 16025 14875 16083 14881
rect 15252 14832 15258 14844
rect 16025 14841 16037 14875
rect 16071 14872 16083 14875
rect 17310 14872 17316 14884
rect 16071 14844 17316 14872
rect 16071 14841 16083 14844
rect 16025 14835 16083 14841
rect 17310 14832 17316 14844
rect 17368 14832 17374 14884
rect 17512 14872 17540 14912
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 17880 14912 18920 14940
rect 17880 14872 17908 14912
rect 17512 14844 17908 14872
rect 17957 14875 18015 14881
rect 17957 14841 17969 14875
rect 18003 14872 18015 14875
rect 18782 14872 18788 14884
rect 18003 14844 18788 14872
rect 18003 14841 18015 14844
rect 17957 14835 18015 14841
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 13998 14804 14004 14816
rect 13959 14776 14004 14804
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 15105 14807 15163 14813
rect 15105 14804 15117 14807
rect 14700 14776 15117 14804
rect 14700 14764 14706 14776
rect 15105 14773 15117 14776
rect 15151 14773 15163 14807
rect 15105 14767 15163 14773
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 16482 14804 16488 14816
rect 15896 14776 16488 14804
rect 15896 14764 15902 14776
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 17770 14804 17776 14816
rect 16724 14776 17776 14804
rect 16724 14764 16730 14776
rect 17770 14764 17776 14776
rect 17828 14804 17834 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 17828 14776 18429 14804
rect 17828 14764 17834 14776
rect 18417 14773 18429 14776
rect 18463 14773 18475 14807
rect 18892 14804 18920 14912
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 20180 14949 20208 15048
rect 20640 15008 20668 15116
rect 21726 15104 21732 15156
rect 21784 15144 21790 15156
rect 22830 15144 22836 15156
rect 21784 15116 22836 15144
rect 21784 15104 21790 15116
rect 22830 15104 22836 15116
rect 22888 15104 22894 15156
rect 24762 15104 24768 15156
rect 24820 15144 24826 15156
rect 26513 15147 26571 15153
rect 26513 15144 26525 15147
rect 24820 15116 26525 15144
rect 24820 15104 24826 15116
rect 26513 15113 26525 15116
rect 26559 15113 26571 15147
rect 26513 15107 26571 15113
rect 27525 15147 27583 15153
rect 27525 15113 27537 15147
rect 27571 15144 27583 15147
rect 28626 15144 28632 15156
rect 27571 15116 28632 15144
rect 27571 15113 27583 15116
rect 27525 15107 27583 15113
rect 28626 15104 28632 15116
rect 28684 15104 28690 15156
rect 28810 15104 28816 15156
rect 28868 15144 28874 15156
rect 30006 15144 30012 15156
rect 28868 15116 30012 15144
rect 28868 15104 28874 15116
rect 30006 15104 30012 15116
rect 30064 15104 30070 15156
rect 30098 15104 30104 15156
rect 30156 15144 30162 15156
rect 30558 15144 30564 15156
rect 30156 15116 30564 15144
rect 30156 15104 30162 15116
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 23382 15076 23388 15088
rect 23046 15048 23388 15076
rect 23382 15036 23388 15048
rect 23440 15036 23446 15088
rect 23477 15079 23535 15085
rect 23477 15045 23489 15079
rect 23523 15076 23535 15079
rect 24578 15076 24584 15088
rect 23523 15048 24584 15076
rect 23523 15045 23535 15048
rect 23477 15039 23535 15045
rect 24578 15036 24584 15048
rect 24636 15036 24642 15088
rect 25222 15036 25228 15088
rect 25280 15036 25286 15088
rect 25958 15036 25964 15088
rect 26016 15076 26022 15088
rect 26234 15076 26240 15088
rect 26016 15048 26240 15076
rect 26016 15036 26022 15048
rect 26234 15036 26240 15048
rect 26292 15036 26298 15088
rect 27798 15036 27804 15088
rect 27856 15076 27862 15088
rect 30190 15076 30196 15088
rect 27856 15048 30196 15076
rect 27856 15036 27862 15048
rect 30190 15036 30196 15048
rect 30248 15036 30254 15088
rect 30466 15036 30472 15088
rect 30524 15076 30530 15088
rect 30837 15079 30895 15085
rect 30837 15076 30849 15079
rect 30524 15048 30849 15076
rect 30524 15036 30530 15048
rect 30837 15045 30849 15048
rect 30883 15045 30895 15079
rect 30837 15039 30895 15045
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 20640 14980 21189 15008
rect 21177 14977 21189 14980
rect 21223 14977 21235 15011
rect 26421 15011 26479 15017
rect 26421 15008 26433 15011
rect 21177 14971 21235 14977
rect 25700 14980 26433 15008
rect 25700 14952 25728 14980
rect 26421 14977 26433 14980
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 26605 15011 26663 15017
rect 26605 14977 26617 15011
rect 26651 15006 26663 15011
rect 27341 15011 27399 15017
rect 26651 14978 26740 15006
rect 26651 14977 26663 14978
rect 26605 14971 26663 14977
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19576 14912 19901 14940
rect 19576 14900 19582 14912
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 19889 14903 19947 14909
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14909 20223 14943
rect 21450 14940 21456 14952
rect 21411 14912 21456 14940
rect 20165 14903 20223 14909
rect 20180 14872 20208 14903
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 21542 14900 21548 14952
rect 21600 14940 21606 14952
rect 22005 14943 22063 14949
rect 22005 14940 22017 14943
rect 21600 14912 22017 14940
rect 21600 14900 21606 14912
rect 22005 14909 22017 14912
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 22738 14900 22744 14952
rect 22796 14940 22802 14952
rect 23753 14943 23811 14949
rect 23753 14940 23765 14943
rect 22796 14912 23765 14940
rect 22796 14900 22802 14912
rect 23753 14909 23765 14912
rect 23799 14909 23811 14943
rect 23753 14903 23811 14909
rect 24213 14943 24271 14949
rect 24213 14909 24225 14943
rect 24259 14909 24271 14943
rect 24213 14903 24271 14909
rect 24489 14943 24547 14949
rect 24489 14909 24501 14943
rect 24535 14940 24547 14943
rect 24578 14940 24584 14952
rect 24535 14912 24584 14940
rect 24535 14909 24547 14912
rect 24489 14903 24547 14909
rect 20806 14872 20812 14884
rect 20180 14844 20812 14872
rect 20806 14832 20812 14844
rect 20864 14872 20870 14884
rect 22370 14872 22376 14884
rect 20864 14844 22376 14872
rect 20864 14832 20870 14844
rect 22370 14832 22376 14844
rect 22428 14832 22434 14884
rect 24228 14872 24256 14903
rect 24578 14900 24584 14912
rect 24636 14900 24642 14952
rect 25498 14900 25504 14952
rect 25556 14940 25562 14952
rect 25682 14940 25688 14952
rect 25556 14912 25688 14940
rect 25556 14900 25562 14912
rect 25682 14900 25688 14912
rect 25740 14900 25746 14952
rect 25958 14900 25964 14952
rect 26016 14940 26022 14952
rect 26016 14912 26464 14940
rect 26016 14900 26022 14912
rect 23676 14844 24256 14872
rect 26436 14872 26464 14912
rect 26712 14872 26740 14978
rect 27341 14977 27353 15011
rect 27387 15008 27399 15011
rect 27706 15008 27712 15020
rect 27387 14980 27712 15008
rect 27387 14977 27399 14980
rect 27341 14971 27399 14977
rect 27706 14968 27712 14980
rect 27764 15008 27770 15020
rect 27982 15008 27988 15020
rect 27764 14980 27988 15008
rect 27764 14968 27770 14980
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 28077 15014 28135 15017
rect 28077 15011 28212 15014
rect 28077 14977 28089 15011
rect 28123 14998 28212 15011
rect 28123 14986 28396 14998
rect 28123 14977 28135 14986
rect 28077 14971 28135 14977
rect 28184 14970 28396 14986
rect 27157 14943 27215 14949
rect 27157 14909 27169 14943
rect 27203 14940 27215 14943
rect 27890 14940 27896 14952
rect 27203 14912 27896 14940
rect 27203 14909 27215 14912
rect 27157 14903 27215 14909
rect 27890 14900 27896 14912
rect 27948 14900 27954 14952
rect 28368 14940 28396 14970
rect 28626 14968 28632 15020
rect 28684 15008 28690 15020
rect 28813 15011 28871 15017
rect 28813 15008 28825 15011
rect 28684 14980 28825 15008
rect 28684 14968 28690 14980
rect 28813 14977 28825 14980
rect 28859 14977 28871 15011
rect 29638 15008 29644 15020
rect 29599 14980 29644 15008
rect 28813 14971 28871 14977
rect 29638 14968 29644 14980
rect 29696 14968 29702 15020
rect 29730 14968 29736 15020
rect 29788 15008 29794 15020
rect 30285 15011 30343 15017
rect 30285 15008 30297 15011
rect 29788 14980 30297 15008
rect 29788 14968 29794 14980
rect 30285 14977 30297 14980
rect 30331 15008 30343 15011
rect 30745 15011 30803 15017
rect 30745 15008 30757 15011
rect 30331 14980 30757 15008
rect 30331 14977 30343 14980
rect 30285 14971 30343 14977
rect 30745 14977 30757 14980
rect 30791 15008 30803 15011
rect 32398 15008 32404 15020
rect 30791 14980 32404 15008
rect 30791 14977 30803 14980
rect 30745 14971 30803 14977
rect 32398 14968 32404 14980
rect 32456 14968 32462 15020
rect 28442 14940 28448 14952
rect 28368 14912 28448 14940
rect 28442 14900 28448 14912
rect 28500 14900 28506 14952
rect 29549 14943 29607 14949
rect 29549 14909 29561 14943
rect 29595 14940 29607 14943
rect 29595 14912 29868 14940
rect 29595 14909 29607 14912
rect 29549 14903 29607 14909
rect 26436 14844 26740 14872
rect 23676 14816 23704 14844
rect 19702 14804 19708 14816
rect 18892 14776 19708 14804
rect 18417 14767 18475 14773
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 20070 14764 20076 14816
rect 20128 14804 20134 14816
rect 21726 14804 21732 14816
rect 20128 14776 21732 14804
rect 20128 14764 20134 14776
rect 21726 14764 21732 14776
rect 21784 14764 21790 14816
rect 22002 14764 22008 14816
rect 22060 14804 22066 14816
rect 22278 14804 22284 14816
rect 22060 14776 22284 14804
rect 22060 14764 22066 14776
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 23658 14764 23664 14816
rect 23716 14764 23722 14816
rect 24228 14804 24256 14844
rect 26878 14832 26884 14884
rect 26936 14872 26942 14884
rect 28626 14872 28632 14884
rect 26936 14844 28632 14872
rect 26936 14832 26942 14844
rect 28626 14832 28632 14844
rect 28684 14832 28690 14884
rect 29178 14872 29184 14884
rect 28736 14844 29184 14872
rect 24486 14804 24492 14816
rect 24228 14776 24492 14804
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 25961 14807 26019 14813
rect 25961 14773 25973 14807
rect 26007 14804 26019 14807
rect 26050 14804 26056 14816
rect 26007 14776 26056 14804
rect 26007 14773 26019 14776
rect 25961 14767 26019 14773
rect 26050 14764 26056 14776
rect 26108 14764 26114 14816
rect 27614 14764 27620 14816
rect 27672 14804 27678 14816
rect 28077 14807 28135 14813
rect 28077 14804 28089 14807
rect 27672 14776 28089 14804
rect 27672 14764 27678 14776
rect 28077 14773 28089 14776
rect 28123 14773 28135 14807
rect 28077 14767 28135 14773
rect 28166 14764 28172 14816
rect 28224 14804 28230 14816
rect 28736 14804 28764 14844
rect 29178 14832 29184 14844
rect 29236 14832 29242 14884
rect 29840 14872 29868 14912
rect 30006 14900 30012 14952
rect 30064 14940 30070 14952
rect 30193 14943 30251 14949
rect 30193 14940 30205 14943
rect 30064 14912 30205 14940
rect 30064 14900 30070 14912
rect 30193 14909 30205 14912
rect 30239 14909 30251 14943
rect 30193 14903 30251 14909
rect 29840 14844 30052 14872
rect 30024 14816 30052 14844
rect 28224 14776 28764 14804
rect 28905 14807 28963 14813
rect 28224 14764 28230 14776
rect 28905 14773 28917 14807
rect 28951 14804 28963 14807
rect 29086 14804 29092 14816
rect 28951 14776 29092 14804
rect 28951 14773 28963 14776
rect 28905 14767 28963 14773
rect 29086 14764 29092 14776
rect 29144 14804 29150 14816
rect 29914 14804 29920 14816
rect 29144 14776 29920 14804
rect 29144 14764 29150 14776
rect 29914 14764 29920 14776
rect 29972 14764 29978 14816
rect 30006 14764 30012 14816
rect 30064 14764 30070 14816
rect 1104 14714 31832 14736
rect 1104 14662 4791 14714
rect 4843 14662 4855 14714
rect 4907 14662 4919 14714
rect 4971 14662 4983 14714
rect 5035 14662 5047 14714
rect 5099 14662 12473 14714
rect 12525 14662 12537 14714
rect 12589 14662 12601 14714
rect 12653 14662 12665 14714
rect 12717 14662 12729 14714
rect 12781 14662 20155 14714
rect 20207 14662 20219 14714
rect 20271 14662 20283 14714
rect 20335 14662 20347 14714
rect 20399 14662 20411 14714
rect 20463 14662 27837 14714
rect 27889 14662 27901 14714
rect 27953 14662 27965 14714
rect 28017 14662 28029 14714
rect 28081 14662 28093 14714
rect 28145 14662 31832 14714
rect 1104 14640 31832 14662
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 14645 14603 14703 14609
rect 11020 14572 14596 14600
rect 11020 14560 11026 14572
rect 12158 14492 12164 14544
rect 12216 14532 12222 14544
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 12216 14504 13645 14532
rect 12216 14492 12222 14504
rect 13633 14501 13645 14504
rect 13679 14532 13691 14535
rect 14366 14532 14372 14544
rect 13679 14504 14372 14532
rect 13679 14501 13691 14504
rect 13633 14495 13691 14501
rect 14366 14492 14372 14504
rect 14424 14492 14430 14544
rect 14568 14532 14596 14572
rect 14645 14569 14657 14603
rect 14691 14600 14703 14603
rect 15470 14600 15476 14612
rect 14691 14572 15476 14600
rect 14691 14569 14703 14572
rect 14645 14563 14703 14569
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 17034 14600 17040 14612
rect 15856 14572 17040 14600
rect 15856 14532 15884 14572
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 17310 14600 17316 14612
rect 17271 14572 17316 14600
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 18046 14600 18052 14612
rect 17420 14572 18052 14600
rect 14568 14504 15884 14532
rect 15933 14535 15991 14541
rect 15933 14501 15945 14535
rect 15979 14532 15991 14535
rect 16942 14532 16948 14544
rect 15979 14504 16948 14532
rect 15979 14501 15991 14504
rect 15933 14495 15991 14501
rect 16942 14492 16948 14504
rect 17000 14492 17006 14544
rect 13078 14464 13084 14476
rect 13039 14436 13084 14464
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 13780 14436 15792 14464
rect 13780 14424 13786 14436
rect 14458 14396 14464 14408
rect 14419 14368 14464 14396
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 14642 14396 14648 14408
rect 14603 14368 14648 14396
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15764 14405 15792 14436
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 17420 14464 17448 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 20438 14600 20444 14612
rect 18288 14572 20444 14600
rect 18288 14560 18294 14572
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 21174 14600 21180 14612
rect 20916 14572 21180 14600
rect 18598 14532 18604 14544
rect 17604 14504 18604 14532
rect 17604 14473 17632 14504
rect 18598 14492 18604 14504
rect 18656 14492 18662 14544
rect 18874 14532 18880 14544
rect 18835 14504 18880 14532
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 19242 14492 19248 14544
rect 19300 14532 19306 14544
rect 20916 14532 20944 14572
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 21450 14560 21456 14612
rect 21508 14600 21514 14612
rect 24581 14603 24639 14609
rect 24581 14600 24593 14603
rect 21508 14572 24593 14600
rect 21508 14560 21514 14572
rect 24581 14569 24593 14572
rect 24627 14569 24639 14603
rect 24581 14563 24639 14569
rect 25406 14560 25412 14612
rect 25464 14600 25470 14612
rect 26786 14600 26792 14612
rect 25464 14572 25636 14600
rect 26747 14572 26792 14600
rect 25464 14560 25470 14572
rect 19300 14504 20944 14532
rect 19300 14492 19306 14504
rect 22370 14492 22376 14544
rect 22428 14532 22434 14544
rect 25133 14535 25191 14541
rect 25133 14532 25145 14535
rect 22428 14504 25145 14532
rect 22428 14492 22434 14504
rect 25133 14501 25145 14504
rect 25179 14532 25191 14535
rect 25498 14532 25504 14544
rect 25179 14504 25504 14532
rect 25179 14501 25191 14504
rect 25133 14495 25191 14501
rect 25498 14492 25504 14504
rect 25556 14492 25562 14544
rect 25608 14532 25636 14572
rect 26786 14560 26792 14572
rect 26844 14560 26850 14612
rect 27154 14560 27160 14612
rect 27212 14600 27218 14612
rect 28813 14603 28871 14609
rect 28813 14600 28825 14603
rect 27212 14572 28825 14600
rect 27212 14560 27218 14572
rect 28813 14569 28825 14572
rect 28859 14569 28871 14603
rect 30466 14600 30472 14612
rect 30427 14572 30472 14600
rect 28813 14563 28871 14569
rect 30466 14560 30472 14572
rect 30524 14560 30530 14612
rect 31297 14603 31355 14609
rect 31297 14569 31309 14603
rect 31343 14600 31355 14603
rect 31386 14600 31392 14612
rect 31343 14572 31392 14600
rect 31343 14569 31355 14572
rect 31297 14563 31355 14569
rect 31386 14560 31392 14572
rect 31444 14560 31450 14612
rect 26878 14532 26884 14544
rect 25608 14504 26884 14532
rect 26878 14492 26884 14504
rect 26936 14492 26942 14544
rect 27709 14535 27767 14541
rect 27709 14501 27721 14535
rect 27755 14532 27767 14535
rect 27798 14532 27804 14544
rect 27755 14504 27804 14532
rect 27755 14501 27767 14504
rect 27709 14495 27767 14501
rect 27798 14492 27804 14504
rect 27856 14492 27862 14544
rect 27890 14492 27896 14544
rect 27948 14532 27954 14544
rect 28442 14532 28448 14544
rect 27948 14504 28448 14532
rect 27948 14492 27954 14504
rect 28442 14492 28448 14504
rect 28500 14492 28506 14544
rect 16356 14436 17448 14464
rect 17589 14467 17647 14473
rect 16356 14424 16362 14436
rect 15105 14399 15163 14405
rect 15105 14398 15117 14399
rect 14936 14370 15117 14398
rect 14366 14288 14372 14340
rect 14424 14328 14430 14340
rect 14936 14328 14964 14370
rect 15105 14365 15117 14370
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16114 14396 16120 14408
rect 15979 14368 16120 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16408 14405 16436 14436
rect 17589 14433 17601 14467
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14464 17739 14467
rect 17862 14464 17868 14476
rect 17727 14436 17868 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 18104 14436 18429 14464
rect 18104 14424 18110 14436
rect 18417 14433 18429 14436
rect 18463 14464 18475 14467
rect 18463 14436 19564 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14365 16451 14399
rect 16666 14396 16672 14408
rect 16627 14368 16672 14396
rect 16393 14359 16451 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 16942 14396 16948 14408
rect 16816 14368 16948 14396
rect 16816 14356 16822 14368
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17310 14396 17316 14408
rect 17092 14368 17316 14396
rect 17092 14356 17098 14368
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 17773 14399 17831 14405
rect 17552 14368 17597 14396
rect 17552 14356 17558 14368
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 18230 14396 18236 14408
rect 17819 14368 18236 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 18555 14368 19441 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 14424 14300 14964 14328
rect 15197 14331 15255 14337
rect 14424 14288 14430 14300
rect 15197 14297 15209 14331
rect 15243 14328 15255 14331
rect 15562 14328 15568 14340
rect 15243 14300 15568 14328
rect 15243 14297 15255 14300
rect 15197 14291 15255 14297
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 15838 14288 15844 14340
rect 15896 14328 15902 14340
rect 16298 14328 16304 14340
rect 15896 14300 16304 14328
rect 15896 14288 15902 14300
rect 16298 14288 16304 14300
rect 16356 14288 16362 14340
rect 16485 14331 16543 14337
rect 16485 14297 16497 14331
rect 16531 14328 16543 14331
rect 17126 14328 17132 14340
rect 16531 14300 17132 14328
rect 16531 14297 16543 14300
rect 16485 14291 16543 14297
rect 17126 14288 17132 14300
rect 17184 14328 17190 14340
rect 18524 14328 18552 14359
rect 17184 14300 18552 14328
rect 19536 14328 19564 14436
rect 19610 14424 19616 14476
rect 19668 14464 19674 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19668 14436 19993 14464
rect 19668 14424 19674 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 21358 14464 21364 14476
rect 19981 14427 20039 14433
rect 20272 14436 21364 14464
rect 19702 14396 19708 14408
rect 19663 14368 19708 14396
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 19797 14331 19855 14337
rect 19797 14328 19809 14331
rect 19536 14300 19809 14328
rect 17184 14288 17190 14300
rect 19797 14297 19809 14300
rect 19843 14297 19855 14331
rect 19797 14291 19855 14297
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 16758 14260 16764 14272
rect 13412 14232 16764 14260
rect 13412 14220 13418 14232
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 16853 14263 16911 14269
rect 16853 14229 16865 14263
rect 16899 14260 16911 14263
rect 19150 14260 19156 14272
rect 16899 14232 19156 14260
rect 16899 14229 16911 14232
rect 16853 14223 16911 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19613 14263 19671 14269
rect 19613 14229 19625 14263
rect 19659 14260 19671 14263
rect 19702 14260 19708 14272
rect 19659 14232 19708 14260
rect 19659 14229 19671 14232
rect 19613 14223 19671 14229
rect 19702 14220 19708 14232
rect 19760 14260 19766 14272
rect 20272 14260 20300 14436
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 21913 14467 21971 14473
rect 21913 14433 21925 14467
rect 21959 14464 21971 14467
rect 23014 14464 23020 14476
rect 21959 14436 23020 14464
rect 21959 14433 21971 14436
rect 21913 14427 21971 14433
rect 23014 14424 23020 14436
rect 23072 14424 23078 14476
rect 24762 14424 24768 14476
rect 24820 14464 24826 14476
rect 26145 14467 26203 14473
rect 26145 14464 26157 14467
rect 24820 14436 26157 14464
rect 24820 14424 24826 14436
rect 26145 14433 26157 14436
rect 26191 14433 26203 14467
rect 26145 14427 26203 14433
rect 26970 14424 26976 14476
rect 27028 14464 27034 14476
rect 28626 14464 28632 14476
rect 27028 14436 27568 14464
rect 27028 14424 27034 14436
rect 22189 14399 22247 14405
rect 22189 14365 22201 14399
rect 22235 14396 22247 14399
rect 22738 14396 22744 14408
rect 22235 14368 22744 14396
rect 22235 14365 22247 14368
rect 22189 14359 22247 14365
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 23201 14399 23259 14405
rect 23201 14365 23213 14399
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14396 23535 14399
rect 25593 14399 25651 14405
rect 25593 14396 25605 14399
rect 23523 14368 25605 14396
rect 23523 14365 23535 14368
rect 23477 14359 23535 14365
rect 25593 14365 25605 14368
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 25961 14399 26019 14405
rect 25961 14365 25973 14399
rect 26007 14396 26019 14399
rect 26050 14396 26056 14408
rect 26007 14368 26056 14396
rect 26007 14365 26019 14368
rect 25961 14359 26019 14365
rect 21450 14288 21456 14340
rect 21508 14288 21514 14340
rect 22830 14288 22836 14340
rect 22888 14328 22894 14340
rect 23216 14328 23244 14359
rect 26050 14356 26056 14368
rect 26108 14356 26114 14408
rect 27430 14396 27436 14408
rect 27391 14368 27436 14396
rect 27430 14356 27436 14368
rect 27488 14356 27494 14408
rect 27540 14405 27568 14436
rect 27724 14436 28632 14464
rect 27724 14405 27752 14436
rect 28626 14424 28632 14436
rect 28684 14424 28690 14476
rect 27525 14399 27583 14405
rect 27525 14365 27537 14399
rect 27571 14365 27583 14399
rect 27525 14359 27583 14365
rect 27709 14399 27767 14405
rect 27709 14365 27721 14399
rect 27755 14365 27767 14399
rect 27709 14359 27767 14365
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14396 28411 14399
rect 28994 14396 29000 14408
rect 28399 14368 28580 14396
rect 28955 14368 29000 14396
rect 28399 14365 28411 14368
rect 28353 14359 28411 14365
rect 22888 14300 24072 14328
rect 22888 14288 22894 14300
rect 19760 14232 20300 14260
rect 19760 14220 19766 14232
rect 20346 14220 20352 14272
rect 20404 14260 20410 14272
rect 20441 14263 20499 14269
rect 20441 14260 20453 14263
rect 20404 14232 20453 14260
rect 20404 14220 20410 14232
rect 20441 14229 20453 14232
rect 20487 14260 20499 14263
rect 21082 14260 21088 14272
rect 20487 14232 21088 14260
rect 20487 14229 20499 14232
rect 20441 14223 20499 14229
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 21174 14220 21180 14272
rect 21232 14260 21238 14272
rect 22002 14260 22008 14272
rect 21232 14232 22008 14260
rect 21232 14220 21238 14232
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 23474 14220 23480 14272
rect 23532 14260 23538 14272
rect 23937 14263 23995 14269
rect 23937 14260 23949 14263
rect 23532 14232 23949 14260
rect 23532 14220 23538 14232
rect 23937 14229 23949 14232
rect 23983 14229 23995 14263
rect 24044 14260 24072 14300
rect 24118 14288 24124 14340
rect 24176 14328 24182 14340
rect 24949 14331 25007 14337
rect 24949 14328 24961 14331
rect 24176 14300 24961 14328
rect 24176 14288 24182 14300
rect 24949 14297 24961 14300
rect 24995 14297 25007 14331
rect 24949 14291 25007 14297
rect 25038 14288 25044 14340
rect 25096 14328 25102 14340
rect 26786 14337 26792 14340
rect 25869 14331 25927 14337
rect 25869 14328 25881 14331
rect 25096 14300 25881 14328
rect 25096 14288 25102 14300
rect 25869 14297 25881 14300
rect 25915 14328 25927 14331
rect 26773 14331 26792 14337
rect 25915 14300 26740 14328
rect 25915 14297 25927 14300
rect 25869 14291 25927 14297
rect 24765 14263 24823 14269
rect 24765 14260 24777 14263
rect 24044 14232 24777 14260
rect 23937 14223 23995 14229
rect 24765 14229 24777 14232
rect 24811 14229 24823 14263
rect 24765 14223 24823 14229
rect 24854 14220 24860 14272
rect 24912 14260 24918 14272
rect 24912 14232 24957 14260
rect 24912 14220 24918 14232
rect 25682 14220 25688 14272
rect 25740 14260 25746 14272
rect 25777 14263 25835 14269
rect 25777 14260 25789 14263
rect 25740 14232 25789 14260
rect 25740 14220 25746 14232
rect 25777 14229 25789 14232
rect 25823 14229 25835 14263
rect 25777 14223 25835 14229
rect 26050 14220 26056 14272
rect 26108 14260 26114 14272
rect 26605 14263 26663 14269
rect 26605 14260 26617 14263
rect 26108 14232 26617 14260
rect 26108 14220 26114 14232
rect 26605 14229 26617 14232
rect 26651 14229 26663 14263
rect 26712 14260 26740 14300
rect 26773 14297 26785 14331
rect 26773 14291 26792 14297
rect 26786 14288 26792 14291
rect 26844 14288 26850 14340
rect 26878 14288 26884 14340
rect 26936 14328 26942 14340
rect 26973 14331 27031 14337
rect 26973 14328 26985 14331
rect 26936 14300 26985 14328
rect 26936 14288 26942 14300
rect 26973 14297 26985 14300
rect 27019 14297 27031 14331
rect 26973 14291 27031 14297
rect 27982 14260 27988 14272
rect 26712 14232 27988 14260
rect 26605 14223 26663 14229
rect 27982 14220 27988 14232
rect 28040 14220 28046 14272
rect 28184 14260 28212 14359
rect 28261 14331 28319 14337
rect 28261 14297 28273 14331
rect 28307 14328 28319 14331
rect 28442 14328 28448 14340
rect 28307 14300 28448 14328
rect 28307 14297 28319 14300
rect 28261 14291 28319 14297
rect 28442 14288 28448 14300
rect 28500 14288 28506 14340
rect 28552 14328 28580 14368
rect 28994 14356 29000 14368
rect 29052 14356 29058 14408
rect 29638 14356 29644 14408
rect 29696 14396 29702 14408
rect 29733 14399 29791 14405
rect 29733 14396 29745 14399
rect 29696 14368 29745 14396
rect 29696 14356 29702 14368
rect 29733 14365 29745 14368
rect 29779 14365 29791 14399
rect 29733 14359 29791 14365
rect 29822 14356 29828 14408
rect 29880 14356 29886 14408
rect 30558 14356 30564 14408
rect 30616 14396 30622 14408
rect 30653 14399 30711 14405
rect 30653 14396 30665 14399
rect 30616 14368 30665 14396
rect 30616 14356 30622 14368
rect 30653 14365 30665 14368
rect 30699 14396 30711 14399
rect 31018 14396 31024 14408
rect 30699 14368 31024 14396
rect 30699 14365 30711 14368
rect 30653 14359 30711 14365
rect 31018 14356 31024 14368
rect 31076 14356 31082 14408
rect 29270 14328 29276 14340
rect 28552 14300 29276 14328
rect 29270 14288 29276 14300
rect 29328 14328 29334 14340
rect 29840 14328 29868 14356
rect 29328 14300 29868 14328
rect 29328 14288 29334 14300
rect 28810 14260 28816 14272
rect 28184 14232 28816 14260
rect 28810 14220 28816 14232
rect 28868 14220 28874 14272
rect 29822 14260 29828 14272
rect 29783 14232 29828 14260
rect 29822 14220 29828 14232
rect 29880 14220 29886 14272
rect 1104 14170 31992 14192
rect 1104 14118 8632 14170
rect 8684 14118 8696 14170
rect 8748 14118 8760 14170
rect 8812 14118 8824 14170
rect 8876 14118 8888 14170
rect 8940 14118 16314 14170
rect 16366 14118 16378 14170
rect 16430 14118 16442 14170
rect 16494 14118 16506 14170
rect 16558 14118 16570 14170
rect 16622 14118 23996 14170
rect 24048 14118 24060 14170
rect 24112 14118 24124 14170
rect 24176 14118 24188 14170
rect 24240 14118 24252 14170
rect 24304 14118 31678 14170
rect 31730 14118 31742 14170
rect 31794 14118 31806 14170
rect 31858 14118 31870 14170
rect 31922 14118 31934 14170
rect 31986 14118 31992 14170
rect 1104 14096 31992 14118
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 13354 14056 13360 14068
rect 13136 14028 13360 14056
rect 13136 14016 13142 14028
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14090 14016 14096 14068
rect 14148 14056 14154 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 14148 14028 15577 14056
rect 14148 14016 14154 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 16209 14059 16267 14065
rect 16209 14025 16221 14059
rect 16255 14056 16267 14059
rect 16255 14028 16574 14056
rect 16255 14025 16267 14028
rect 16209 14019 16267 14025
rect 14366 13988 14372 14000
rect 14327 13960 14372 13988
rect 14366 13948 14372 13960
rect 14424 13988 14430 14000
rect 15194 13988 15200 14000
rect 14424 13960 15200 13988
rect 14424 13948 14430 13960
rect 15194 13948 15200 13960
rect 15252 13988 15258 14000
rect 15252 13960 16160 13988
rect 15252 13948 15258 13960
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 14516 13892 15485 13920
rect 14516 13880 14522 13892
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 15654 13920 15660 13932
rect 15615 13892 15660 13920
rect 15473 13883 15531 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 14921 13855 14979 13861
rect 14921 13852 14933 13855
rect 14792 13824 14933 13852
rect 14792 13812 14798 13824
rect 14921 13821 14933 13824
rect 14967 13821 14979 13855
rect 15488 13852 15516 13883
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 16132 13929 16160 13960
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16390 13920 16396 13932
rect 16163 13892 16396 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 16546 13920 16574 14028
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 16816 14028 17141 14056
rect 16816 14016 16822 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17129 14019 17187 14025
rect 18230 14016 18236 14068
rect 18288 14056 18294 14068
rect 21085 14059 21143 14065
rect 21085 14056 21097 14059
rect 18288 14028 21097 14056
rect 18288 14016 18294 14028
rect 21085 14025 21097 14028
rect 21131 14025 21143 14059
rect 21085 14019 21143 14025
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 23658 14056 23664 14068
rect 22060 14028 23664 14056
rect 22060 14016 22066 14028
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 23753 14059 23811 14065
rect 23753 14025 23765 14059
rect 23799 14056 23811 14059
rect 23842 14056 23848 14068
rect 23799 14028 23848 14056
rect 23799 14025 23811 14028
rect 23753 14019 23811 14025
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 25435 14059 25493 14065
rect 25435 14025 25447 14059
rect 25481 14056 25493 14059
rect 27614 14056 27620 14068
rect 25481 14028 27620 14056
rect 25481 14025 25493 14028
rect 25435 14019 25493 14025
rect 27614 14016 27620 14028
rect 27672 14016 27678 14068
rect 27893 14059 27951 14065
rect 27893 14025 27905 14059
rect 27939 14056 27951 14059
rect 28626 14056 28632 14068
rect 27939 14028 28632 14056
rect 27939 14025 27951 14028
rect 27893 14019 27951 14025
rect 28626 14016 28632 14028
rect 28684 14016 28690 14068
rect 28718 14016 28724 14068
rect 28776 14056 28782 14068
rect 30006 14056 30012 14068
rect 28776 14028 30012 14056
rect 28776 14016 28782 14028
rect 30006 14016 30012 14028
rect 30064 14016 30070 14068
rect 17218 13988 17224 14000
rect 17179 13960 17224 13988
rect 17218 13948 17224 13960
rect 17276 13948 17282 14000
rect 19426 13988 19432 14000
rect 18432 13960 19432 13988
rect 16546 13892 16804 13920
rect 16776 13864 16804 13892
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17402 13920 17408 13932
rect 17184 13892 17229 13920
rect 17363 13892 17408 13920
rect 17184 13880 17190 13892
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17862 13880 17868 13932
rect 17920 13920 17926 13932
rect 18046 13920 18052 13932
rect 17920 13892 18052 13920
rect 17920 13880 17926 13892
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 16666 13852 16672 13864
rect 15488 13824 16672 13852
rect 14921 13815 14979 13821
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 16758 13812 16764 13864
rect 16816 13812 16822 13864
rect 18141 13855 18199 13861
rect 16868 13824 17172 13852
rect 13998 13744 14004 13796
rect 14056 13784 14062 13796
rect 16868 13784 16896 13824
rect 14056 13756 16896 13784
rect 17144 13784 17172 13824
rect 18141 13821 18153 13855
rect 18187 13852 18199 13855
rect 18322 13852 18328 13864
rect 18187 13824 18328 13852
rect 18187 13821 18199 13824
rect 18141 13815 18199 13821
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 18432 13861 18460 13960
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 19610 13948 19616 14000
rect 19668 13948 19674 14000
rect 20530 13948 20536 14000
rect 20588 13988 20594 14000
rect 21237 13991 21295 13997
rect 21237 13988 21249 13991
rect 20588 13960 21249 13988
rect 20588 13948 20594 13960
rect 21237 13957 21249 13960
rect 21283 13957 21295 13991
rect 21237 13951 21295 13957
rect 21453 13991 21511 13997
rect 21453 13957 21465 13991
rect 21499 13988 21511 13991
rect 21726 13988 21732 14000
rect 21499 13960 21732 13988
rect 21499 13957 21511 13960
rect 21453 13951 21511 13957
rect 21726 13948 21732 13960
rect 21784 13948 21790 14000
rect 25225 13991 25283 13997
rect 23506 13960 25176 13988
rect 18690 13880 18696 13932
rect 18748 13920 18754 13932
rect 18877 13923 18935 13929
rect 18877 13920 18889 13923
rect 18748 13892 18889 13920
rect 18748 13880 18754 13892
rect 18877 13889 18889 13892
rect 18923 13889 18935 13923
rect 22002 13920 22008 13932
rect 21963 13892 22008 13920
rect 18877 13883 18935 13889
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 23842 13920 23848 13932
rect 23584 13892 23848 13920
rect 18417 13855 18475 13861
rect 18417 13821 18429 13855
rect 18463 13821 18475 13855
rect 19153 13855 19211 13861
rect 19153 13852 19165 13855
rect 18417 13815 18475 13821
rect 18524 13824 19165 13852
rect 18524 13784 18552 13824
rect 19153 13821 19165 13824
rect 19199 13821 19211 13855
rect 19153 13815 19211 13821
rect 20438 13812 20444 13864
rect 20496 13852 20502 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20496 13824 20637 13852
rect 20496 13812 20502 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 21726 13812 21732 13864
rect 21784 13852 21790 13864
rect 23584 13852 23612 13892
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 24581 13923 24639 13929
rect 24581 13920 24593 13923
rect 24452 13892 24593 13920
rect 24452 13880 24458 13892
rect 24581 13889 24593 13892
rect 24627 13920 24639 13923
rect 24762 13920 24768 13932
rect 24627 13892 24768 13920
rect 24627 13889 24639 13892
rect 24581 13883 24639 13889
rect 24762 13880 24768 13892
rect 24820 13880 24826 13932
rect 21784 13824 23612 13852
rect 21784 13812 21790 13824
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23716 13824 24225 13852
rect 23716 13812 23722 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 24489 13855 24547 13861
rect 24489 13821 24501 13855
rect 24535 13821 24547 13855
rect 25148 13852 25176 13960
rect 25225 13957 25237 13991
rect 25271 13988 25283 13991
rect 26053 13991 26111 13997
rect 25271 13960 25452 13988
rect 25271 13957 25283 13960
rect 25225 13951 25283 13957
rect 25424 13932 25452 13960
rect 26053 13957 26065 13991
rect 26099 13988 26111 13991
rect 26418 13988 26424 14000
rect 26099 13960 26424 13988
rect 26099 13957 26111 13960
rect 26053 13951 26111 13957
rect 26418 13948 26424 13960
rect 26476 13948 26482 14000
rect 28994 13988 29000 14000
rect 26804 13960 29000 13988
rect 25406 13880 25412 13932
rect 25464 13880 25470 13932
rect 25498 13880 25504 13932
rect 25556 13920 25562 13932
rect 26142 13920 26148 13932
rect 25556 13892 26148 13920
rect 25556 13880 25562 13892
rect 26142 13880 26148 13892
rect 26200 13880 26206 13932
rect 26237 13923 26295 13929
rect 26237 13889 26249 13923
rect 26283 13920 26295 13923
rect 26694 13920 26700 13932
rect 26283 13892 26700 13920
rect 26283 13889 26295 13892
rect 26237 13883 26295 13889
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 26804 13852 26832 13960
rect 28994 13948 29000 13960
rect 29052 13948 29058 14000
rect 26878 13880 26884 13932
rect 26936 13920 26942 13932
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 26936 13892 27169 13920
rect 26936 13880 26942 13892
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 27341 13923 27399 13929
rect 27341 13889 27353 13923
rect 27387 13889 27399 13923
rect 27798 13920 27804 13932
rect 27759 13892 27804 13920
rect 27341 13883 27399 13889
rect 27246 13852 27252 13864
rect 25148 13824 25544 13852
rect 24489 13815 24547 13821
rect 17144 13756 18552 13784
rect 14056 13744 14062 13756
rect 20806 13744 20812 13796
rect 20864 13784 20870 13796
rect 20990 13784 20996 13796
rect 20864 13756 20996 13784
rect 20864 13744 20870 13756
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 23382 13744 23388 13796
rect 23440 13784 23446 13796
rect 24504 13784 24532 13815
rect 24762 13784 24768 13796
rect 23440 13756 24768 13784
rect 23440 13744 23446 13756
rect 24762 13744 24768 13756
rect 24820 13744 24826 13796
rect 25038 13744 25044 13796
rect 25096 13744 25102 13796
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 18414 13716 18420 13728
rect 15436 13688 18420 13716
rect 15436 13676 15442 13688
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 21269 13719 21327 13725
rect 21269 13716 21281 13719
rect 19208 13688 21281 13716
rect 19208 13676 19214 13688
rect 21269 13685 21281 13688
rect 21315 13685 21327 13719
rect 21269 13679 21327 13685
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 22262 13719 22320 13725
rect 22262 13716 22274 13719
rect 21416 13688 22274 13716
rect 21416 13676 21422 13688
rect 22262 13685 22274 13688
rect 22308 13685 22320 13719
rect 22262 13679 22320 13685
rect 24210 13676 24216 13728
rect 24268 13716 24274 13728
rect 25056 13716 25084 13744
rect 25406 13716 25412 13728
rect 24268 13688 25084 13716
rect 25367 13688 25412 13716
rect 24268 13676 24274 13688
rect 25406 13676 25412 13688
rect 25464 13676 25470 13728
rect 25516 13716 25544 13824
rect 25608 13824 26832 13852
rect 27207 13824 27252 13852
rect 25608 13793 25636 13824
rect 27246 13812 27252 13824
rect 27304 13812 27310 13864
rect 25593 13787 25651 13793
rect 25593 13753 25605 13787
rect 25639 13753 25651 13787
rect 25593 13747 25651 13753
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 26786 13784 26792 13796
rect 26292 13756 26792 13784
rect 26292 13744 26298 13756
rect 26786 13744 26792 13756
rect 26844 13784 26850 13796
rect 27356 13784 27384 13883
rect 27798 13880 27804 13892
rect 27856 13880 27862 13932
rect 27985 13923 28043 13929
rect 27985 13889 27997 13923
rect 28031 13920 28043 13923
rect 28074 13920 28080 13932
rect 28031 13892 28080 13920
rect 28031 13889 28043 13892
rect 27985 13883 28043 13889
rect 28074 13880 28080 13892
rect 28132 13880 28138 13932
rect 28442 13920 28448 13932
rect 28403 13892 28448 13920
rect 28442 13880 28448 13892
rect 28500 13880 28506 13932
rect 28629 13923 28687 13929
rect 28629 13889 28641 13923
rect 28675 13889 28687 13923
rect 28629 13883 28687 13889
rect 26844 13756 27384 13784
rect 26844 13744 26850 13756
rect 27982 13744 27988 13796
rect 28040 13784 28046 13796
rect 28644 13784 28672 13883
rect 28902 13880 28908 13932
rect 28960 13920 28966 13932
rect 28960 13892 29224 13920
rect 28960 13880 28966 13892
rect 29196 13852 29224 13892
rect 29270 13880 29276 13932
rect 29328 13920 29334 13932
rect 29730 13920 29736 13932
rect 29328 13892 29736 13920
rect 29328 13880 29334 13892
rect 29730 13880 29736 13892
rect 29788 13880 29794 13932
rect 30653 13923 30711 13929
rect 30653 13889 30665 13923
rect 30699 13920 30711 13923
rect 30834 13920 30840 13932
rect 30699 13892 30840 13920
rect 30699 13889 30711 13892
rect 30653 13883 30711 13889
rect 30834 13880 30840 13892
rect 30892 13880 30898 13932
rect 31297 13923 31355 13929
rect 31297 13889 31309 13923
rect 31343 13920 31355 13923
rect 31478 13920 31484 13932
rect 31343 13892 31484 13920
rect 31343 13889 31355 13892
rect 31297 13883 31355 13889
rect 31478 13880 31484 13892
rect 31536 13880 31542 13932
rect 30009 13855 30067 13861
rect 30009 13852 30021 13855
rect 29196 13824 30021 13852
rect 30009 13821 30021 13824
rect 30055 13821 30067 13855
rect 30009 13815 30067 13821
rect 28040 13756 28672 13784
rect 28040 13744 28046 13756
rect 25682 13716 25688 13728
rect 25516 13688 25688 13716
rect 25682 13676 25688 13688
rect 25740 13676 25746 13728
rect 25958 13676 25964 13728
rect 26016 13716 26022 13728
rect 27890 13716 27896 13728
rect 26016 13688 27896 13716
rect 26016 13676 26022 13688
rect 27890 13676 27896 13688
rect 27948 13676 27954 13728
rect 28445 13719 28503 13725
rect 28445 13685 28457 13719
rect 28491 13716 28503 13719
rect 28994 13716 29000 13728
rect 28491 13688 29000 13716
rect 28491 13685 28503 13688
rect 28445 13679 28503 13685
rect 28994 13676 29000 13688
rect 29052 13676 29058 13728
rect 29178 13716 29184 13728
rect 29139 13688 29184 13716
rect 29178 13676 29184 13688
rect 29236 13676 29242 13728
rect 1104 13626 31832 13648
rect 1104 13574 4791 13626
rect 4843 13574 4855 13626
rect 4907 13574 4919 13626
rect 4971 13574 4983 13626
rect 5035 13574 5047 13626
rect 5099 13574 12473 13626
rect 12525 13574 12537 13626
rect 12589 13574 12601 13626
rect 12653 13574 12665 13626
rect 12717 13574 12729 13626
rect 12781 13574 20155 13626
rect 20207 13574 20219 13626
rect 20271 13574 20283 13626
rect 20335 13574 20347 13626
rect 20399 13574 20411 13626
rect 20463 13574 27837 13626
rect 27889 13574 27901 13626
rect 27953 13574 27965 13626
rect 28017 13574 28029 13626
rect 28081 13574 28093 13626
rect 28145 13574 31832 13626
rect 1104 13552 31832 13574
rect 15194 13512 15200 13524
rect 15155 13484 15200 13512
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 16298 13512 16304 13524
rect 15344 13484 16304 13512
rect 15344 13472 15350 13484
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 17865 13515 17923 13521
rect 16408 13484 17730 13512
rect 14826 13404 14832 13456
rect 14884 13444 14890 13456
rect 16408 13444 16436 13484
rect 14884 13416 16436 13444
rect 16485 13447 16543 13453
rect 14884 13404 14890 13416
rect 16485 13413 16497 13447
rect 16531 13444 16543 13447
rect 16942 13444 16948 13456
rect 16531 13416 16948 13444
rect 16531 13413 16543 13416
rect 16485 13407 16543 13413
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 15838 13376 15844 13388
rect 15799 13348 15844 13376
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 16022 13336 16028 13388
rect 16080 13336 16086 13388
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 15927 13311 15985 13317
rect 15927 13277 15939 13311
rect 15973 13302 15985 13311
rect 16040 13302 16068 13336
rect 17702 13324 17730 13484
rect 17865 13481 17877 13515
rect 17911 13512 17923 13515
rect 19242 13512 19248 13524
rect 17911 13484 19248 13512
rect 17911 13481 17923 13484
rect 17865 13475 17923 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 25041 13515 25099 13521
rect 19392 13484 23704 13512
rect 19392 13472 19398 13484
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 19610 13444 19616 13456
rect 18840 13416 19616 13444
rect 18840 13404 18846 13416
rect 19610 13404 19616 13416
rect 19668 13404 19674 13456
rect 23676 13444 23704 13484
rect 25041 13481 25053 13515
rect 25087 13512 25099 13515
rect 26970 13512 26976 13524
rect 25087 13484 26976 13512
rect 25087 13481 25099 13484
rect 25041 13475 25099 13481
rect 26970 13472 26976 13484
rect 27028 13472 27034 13524
rect 27338 13512 27344 13524
rect 27299 13484 27344 13512
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 27893 13515 27951 13521
rect 27893 13481 27905 13515
rect 27939 13512 27951 13515
rect 28166 13512 28172 13524
rect 27939 13484 28172 13512
rect 27939 13481 27951 13484
rect 27893 13475 27951 13481
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 28534 13512 28540 13524
rect 28495 13484 28540 13512
rect 28534 13472 28540 13484
rect 28592 13472 28598 13524
rect 30006 13512 30012 13524
rect 29967 13484 30012 13512
rect 30006 13472 30012 13484
rect 30064 13472 30070 13524
rect 30650 13472 30656 13524
rect 30708 13512 30714 13524
rect 31113 13515 31171 13521
rect 31113 13512 31125 13515
rect 30708 13484 31125 13512
rect 30708 13472 30714 13484
rect 31113 13481 31125 13484
rect 31159 13481 31171 13515
rect 31113 13475 31171 13481
rect 25225 13447 25283 13453
rect 25225 13444 25237 13447
rect 23676 13416 25237 13444
rect 25225 13413 25237 13416
rect 25271 13413 25283 13447
rect 26421 13447 26479 13453
rect 26421 13444 26433 13447
rect 25225 13407 25283 13413
rect 25332 13416 26433 13444
rect 18414 13376 18420 13388
rect 18375 13348 18420 13376
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 18877 13379 18935 13385
rect 18877 13376 18889 13379
rect 18616 13348 18889 13376
rect 15973 13277 16068 13302
rect 15927 13274 16068 13277
rect 15927 13271 15985 13274
rect 15764 13240 15792 13271
rect 16206 13268 16212 13320
rect 16264 13308 16270 13320
rect 16390 13308 16396 13320
rect 16264 13280 16396 13308
rect 16264 13268 16270 13280
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 17034 13308 17040 13320
rect 16995 13280 17040 13308
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 17696 13317 17730 13324
rect 17681 13311 17739 13317
rect 17681 13277 17693 13311
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13277 17923 13311
rect 18506 13308 18512 13320
rect 18467 13280 18512 13308
rect 17865 13271 17923 13277
rect 16942 13240 16948 13252
rect 15764 13212 16948 13240
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 17880 13240 17908 13271
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 17052 13212 17908 13240
rect 18616 13240 18644 13348
rect 18877 13345 18889 13348
rect 18923 13345 18935 13379
rect 19429 13379 19487 13385
rect 19429 13376 19441 13379
rect 18877 13339 18935 13345
rect 19168 13348 19441 13376
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 19168 13308 19196 13348
rect 19429 13345 19441 13348
rect 19475 13345 19487 13379
rect 21358 13376 21364 13388
rect 19429 13339 19487 13345
rect 19536 13348 21364 13376
rect 18748 13280 19196 13308
rect 18748 13268 18754 13280
rect 19536 13240 19564 13348
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 21637 13379 21695 13385
rect 21637 13345 21649 13379
rect 21683 13376 21695 13379
rect 22002 13376 22008 13388
rect 21683 13348 22008 13376
rect 21683 13345 21695 13348
rect 21637 13339 21695 13345
rect 22002 13336 22008 13348
rect 22060 13336 22066 13388
rect 23385 13379 23443 13385
rect 23385 13345 23397 13379
rect 23431 13376 23443 13379
rect 24210 13376 24216 13388
rect 23431 13348 24216 13376
rect 23431 13345 23443 13348
rect 23385 13339 23443 13345
rect 24210 13336 24216 13348
rect 24268 13336 24274 13388
rect 24854 13336 24860 13388
rect 24912 13376 24918 13388
rect 25332 13376 25360 13416
rect 26421 13413 26433 13416
rect 26467 13444 26479 13447
rect 27706 13444 27712 13456
rect 26467 13416 27712 13444
rect 26467 13413 26479 13416
rect 26421 13407 26479 13413
rect 27706 13404 27712 13416
rect 27764 13404 27770 13456
rect 24912 13348 25360 13376
rect 25757 13379 25815 13385
rect 24912 13336 24918 13348
rect 25757 13345 25769 13379
rect 25803 13376 25815 13379
rect 30653 13379 30711 13385
rect 25803 13348 27200 13376
rect 25803 13345 25815 13348
rect 25757 13339 25815 13345
rect 19794 13268 19800 13320
rect 19852 13268 19858 13320
rect 21177 13311 21235 13317
rect 21177 13277 21189 13311
rect 21223 13277 21235 13311
rect 24026 13308 24032 13320
rect 23987 13280 24032 13308
rect 21177 13271 21235 13277
rect 20901 13243 20959 13249
rect 20901 13240 20913 13243
rect 18616 13212 19564 13240
rect 20824 13212 20913 13240
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 17052 13172 17080 13212
rect 14332 13144 17080 13172
rect 17129 13175 17187 13181
rect 14332 13132 14338 13144
rect 17129 13141 17141 13175
rect 17175 13172 17187 13175
rect 18874 13172 18880 13184
rect 17175 13144 18880 13172
rect 17175 13141 17187 13144
rect 17129 13135 17187 13141
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19610 13132 19616 13184
rect 19668 13172 19674 13184
rect 20824 13172 20852 13212
rect 20901 13209 20913 13212
rect 20947 13209 20959 13243
rect 20901 13203 20959 13209
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 21192 13240 21220 13271
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 25958 13308 25964 13320
rect 24872 13280 25728 13308
rect 25919 13280 25964 13308
rect 21048 13212 21220 13240
rect 21048 13200 21054 13212
rect 21358 13200 21364 13252
rect 21416 13240 21422 13252
rect 21913 13243 21971 13249
rect 21913 13240 21925 13243
rect 21416 13212 21925 13240
rect 21416 13200 21422 13212
rect 21913 13209 21925 13212
rect 21959 13209 21971 13243
rect 21913 13203 21971 13209
rect 22646 13200 22652 13252
rect 22704 13200 22710 13252
rect 24872 13249 24900 13280
rect 24857 13243 24915 13249
rect 24857 13209 24869 13243
rect 24903 13209 24915 13243
rect 24857 13203 24915 13209
rect 25073 13243 25131 13249
rect 25073 13209 25085 13243
rect 25119 13240 25131 13243
rect 25498 13240 25504 13252
rect 25119 13212 25504 13240
rect 25119 13209 25131 13212
rect 25073 13203 25131 13209
rect 25498 13200 25504 13212
rect 25556 13200 25562 13252
rect 25700 13249 25728 13280
rect 25958 13268 25964 13280
rect 26016 13268 26022 13320
rect 27172 13317 27200 13348
rect 30653 13345 30665 13379
rect 30699 13376 30711 13379
rect 30742 13376 30748 13388
rect 30699 13348 30748 13376
rect 30699 13345 30711 13348
rect 30653 13339 30711 13345
rect 30742 13336 30748 13348
rect 30800 13336 30806 13388
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 27341 13311 27399 13317
rect 27341 13277 27353 13311
rect 27387 13308 27399 13311
rect 27430 13308 27436 13320
rect 27387 13280 27436 13308
rect 27387 13277 27399 13280
rect 27341 13271 27399 13277
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 27522 13268 27528 13320
rect 27580 13308 27586 13320
rect 27801 13311 27859 13317
rect 27801 13308 27813 13311
rect 27580 13280 27813 13308
rect 27580 13268 27586 13280
rect 27801 13277 27813 13280
rect 27847 13308 27859 13311
rect 28629 13311 28687 13317
rect 28629 13308 28641 13311
rect 27847 13280 28641 13308
rect 27847 13277 27859 13280
rect 27801 13271 27859 13277
rect 28629 13277 28641 13280
rect 28675 13308 28687 13311
rect 29270 13308 29276 13320
rect 28675 13280 29276 13308
rect 28675 13277 28687 13280
rect 28629 13271 28687 13277
rect 29270 13268 29276 13280
rect 29328 13268 29334 13320
rect 31202 13268 31208 13320
rect 31260 13308 31266 13320
rect 31297 13311 31355 13317
rect 31297 13308 31309 13311
rect 31260 13280 31309 13308
rect 31260 13268 31266 13280
rect 31297 13277 31309 13280
rect 31343 13277 31355 13311
rect 31297 13271 31355 13277
rect 25685 13243 25743 13249
rect 25685 13209 25697 13243
rect 25731 13240 25743 13243
rect 26142 13240 26148 13252
rect 25731 13212 26148 13240
rect 25731 13209 25743 13212
rect 25685 13203 25743 13209
rect 26142 13200 26148 13212
rect 26200 13200 26206 13252
rect 26605 13243 26663 13249
rect 26605 13209 26617 13243
rect 26651 13240 26663 13243
rect 27614 13240 27620 13252
rect 26651 13212 27620 13240
rect 26651 13209 26663 13212
rect 26605 13203 26663 13209
rect 27614 13200 27620 13212
rect 27672 13200 27678 13252
rect 19668 13144 20852 13172
rect 19668 13132 19674 13144
rect 22278 13132 22284 13184
rect 22336 13172 22342 13184
rect 23845 13175 23903 13181
rect 23845 13172 23857 13175
rect 22336 13144 23857 13172
rect 22336 13132 22342 13144
rect 23845 13141 23857 13144
rect 23891 13141 23903 13175
rect 23845 13135 23903 13141
rect 25406 13132 25412 13184
rect 25464 13172 25470 13184
rect 25869 13175 25927 13181
rect 25869 13172 25881 13175
rect 25464 13144 25881 13172
rect 25464 13132 25470 13144
rect 25869 13141 25881 13144
rect 25915 13172 25927 13175
rect 28258 13172 28264 13184
rect 25915 13144 28264 13172
rect 25915 13141 25927 13144
rect 25869 13135 25927 13141
rect 28258 13132 28264 13144
rect 28316 13132 28322 13184
rect 28902 13132 28908 13184
rect 28960 13172 28966 13184
rect 29089 13175 29147 13181
rect 29089 13172 29101 13175
rect 28960 13144 29101 13172
rect 28960 13132 28966 13144
rect 29089 13141 29101 13144
rect 29135 13141 29147 13175
rect 29089 13135 29147 13141
rect 1104 13082 31992 13104
rect 1104 13030 8632 13082
rect 8684 13030 8696 13082
rect 8748 13030 8760 13082
rect 8812 13030 8824 13082
rect 8876 13030 8888 13082
rect 8940 13030 16314 13082
rect 16366 13030 16378 13082
rect 16430 13030 16442 13082
rect 16494 13030 16506 13082
rect 16558 13030 16570 13082
rect 16622 13030 23996 13082
rect 24048 13030 24060 13082
rect 24112 13030 24124 13082
rect 24176 13030 24188 13082
rect 24240 13030 24252 13082
rect 24304 13030 31678 13082
rect 31730 13030 31742 13082
rect 31794 13030 31806 13082
rect 31858 13030 31870 13082
rect 31922 13030 31934 13082
rect 31986 13030 31992 13082
rect 1104 13008 31992 13030
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 15896 12940 22324 12968
rect 15896 12928 15902 12940
rect 16206 12900 16212 12912
rect 16167 12872 16212 12900
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 18138 12900 18144 12912
rect 17604 12872 18144 12900
rect 16224 12832 16252 12860
rect 17604 12841 17632 12872
rect 18138 12860 18144 12872
rect 18196 12900 18202 12912
rect 18196 12872 18368 12900
rect 18196 12860 18202 12872
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16224 12804 16957 12832
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 17770 12832 17776 12844
rect 17731 12804 17776 12832
rect 17589 12795 17647 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18230 12832 18236 12844
rect 18191 12804 18236 12832
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 18340 12832 18368 12872
rect 18414 12860 18420 12912
rect 18472 12900 18478 12912
rect 19045 12903 19103 12909
rect 19045 12900 19057 12903
rect 18472 12872 19057 12900
rect 18472 12860 18478 12872
rect 19045 12869 19057 12872
rect 19091 12900 19103 12903
rect 19150 12900 19156 12912
rect 19091 12872 19156 12900
rect 19091 12869 19103 12872
rect 19045 12863 19103 12869
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 19242 12860 19248 12912
rect 19300 12900 19306 12912
rect 19981 12903 20039 12909
rect 19981 12900 19993 12903
rect 19300 12872 19345 12900
rect 19628 12872 19993 12900
rect 19300 12860 19306 12872
rect 18506 12832 18512 12844
rect 18340 12804 18512 12832
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12764 17095 12767
rect 18782 12764 18788 12776
rect 17083 12736 18788 12764
rect 17083 12733 17095 12736
rect 17037 12727 17095 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 18417 12699 18475 12705
rect 16724 12668 18092 12696
rect 16724 12656 16730 12668
rect 17681 12631 17739 12637
rect 17681 12597 17693 12631
rect 17727 12628 17739 12631
rect 17954 12628 17960 12640
rect 17727 12600 17960 12628
rect 17727 12597 17739 12600
rect 17681 12591 17739 12597
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18064 12628 18092 12668
rect 18417 12665 18429 12699
rect 18463 12696 18475 12699
rect 19518 12696 19524 12708
rect 18463 12668 19524 12696
rect 18463 12665 18475 12668
rect 18417 12659 18475 12665
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 18877 12631 18935 12637
rect 18877 12628 18889 12631
rect 18064 12600 18889 12628
rect 18877 12597 18889 12600
rect 18923 12597 18935 12631
rect 19058 12628 19064 12640
rect 19019 12600 19064 12628
rect 18877 12591 18935 12597
rect 19058 12588 19064 12600
rect 19116 12588 19122 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19628 12628 19656 12872
rect 19981 12869 19993 12872
rect 20027 12869 20039 12903
rect 19981 12863 20039 12869
rect 20990 12860 20996 12912
rect 21048 12860 21054 12912
rect 22296 12909 22324 12940
rect 23842 12928 23848 12980
rect 23900 12968 23906 12980
rect 24305 12971 24363 12977
rect 24305 12968 24317 12971
rect 23900 12940 24317 12968
rect 23900 12928 23906 12940
rect 24305 12937 24317 12940
rect 24351 12968 24363 12971
rect 25682 12968 25688 12980
rect 24351 12940 25688 12968
rect 24351 12937 24363 12940
rect 24305 12931 24363 12937
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 25777 12971 25835 12977
rect 25777 12937 25789 12971
rect 25823 12968 25835 12971
rect 25866 12968 25872 12980
rect 25823 12940 25872 12968
rect 25823 12937 25835 12940
rect 25777 12931 25835 12937
rect 25866 12928 25872 12940
rect 25924 12928 25930 12980
rect 26421 12971 26479 12977
rect 26421 12937 26433 12971
rect 26467 12968 26479 12971
rect 27154 12968 27160 12980
rect 26467 12940 27160 12968
rect 26467 12937 26479 12940
rect 26421 12931 26479 12937
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 27249 12971 27307 12977
rect 27249 12937 27261 12971
rect 27295 12968 27307 12971
rect 27338 12968 27344 12980
rect 27295 12940 27344 12968
rect 27295 12937 27307 12940
rect 27249 12931 27307 12937
rect 27338 12928 27344 12940
rect 27396 12928 27402 12980
rect 22281 12903 22339 12909
rect 22281 12869 22293 12903
rect 22327 12869 22339 12903
rect 29822 12900 29828 12912
rect 23506 12872 29828 12900
rect 22281 12863 22339 12869
rect 29822 12860 29828 12872
rect 29880 12860 29886 12912
rect 22002 12832 22008 12844
rect 21963 12804 22008 12832
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 24210 12832 24216 12844
rect 24171 12804 24216 12832
rect 24210 12792 24216 12804
rect 24268 12792 24274 12844
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 24949 12835 25007 12841
rect 24949 12832 24961 12835
rect 24912 12804 24961 12832
rect 24912 12792 24918 12804
rect 24949 12801 24961 12804
rect 24995 12801 25007 12835
rect 24949 12795 25007 12801
rect 25038 12792 25044 12844
rect 25096 12832 25102 12844
rect 25225 12835 25283 12841
rect 25096 12804 25141 12832
rect 25096 12792 25102 12804
rect 25225 12801 25237 12835
rect 25271 12832 25283 12835
rect 25406 12832 25412 12844
rect 25271 12804 25412 12832
rect 25271 12801 25283 12804
rect 25225 12795 25283 12801
rect 25406 12792 25412 12804
rect 25464 12792 25470 12844
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12832 25927 12835
rect 26234 12832 26240 12844
rect 25915 12804 26240 12832
rect 25915 12801 25927 12804
rect 25869 12795 25927 12801
rect 26234 12792 26240 12804
rect 26292 12792 26298 12844
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12832 26387 12835
rect 26786 12832 26792 12844
rect 26375 12804 26792 12832
rect 26375 12801 26387 12804
rect 26329 12795 26387 12801
rect 26786 12792 26792 12804
rect 26844 12832 26850 12844
rect 26970 12832 26976 12844
rect 26844 12804 26976 12832
rect 26844 12792 26850 12804
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12832 27215 12835
rect 27522 12832 27528 12844
rect 27203 12804 27528 12832
rect 27203 12801 27215 12804
rect 27157 12795 27215 12801
rect 27522 12792 27528 12804
rect 27580 12792 27586 12844
rect 31294 12832 31300 12844
rect 31255 12804 31300 12832
rect 31294 12792 31300 12804
rect 31352 12792 31358 12844
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12764 19763 12767
rect 20622 12764 20628 12776
rect 19751 12736 20628 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 20714 12724 20720 12776
rect 20772 12764 20778 12776
rect 22020 12764 22048 12792
rect 20772 12736 22048 12764
rect 20772 12724 20778 12736
rect 23014 12724 23020 12776
rect 23072 12764 23078 12776
rect 23753 12767 23811 12773
rect 23753 12764 23765 12767
rect 23072 12736 23765 12764
rect 23072 12724 23078 12736
rect 23753 12733 23765 12736
rect 23799 12764 23811 12767
rect 24762 12764 24768 12776
rect 23799 12736 24768 12764
rect 23799 12733 23811 12736
rect 23753 12727 23811 12733
rect 24762 12724 24768 12736
rect 24820 12724 24826 12776
rect 26602 12764 26608 12776
rect 25056 12736 26608 12764
rect 24394 12656 24400 12708
rect 24452 12696 24458 12708
rect 25056 12696 25084 12736
rect 26602 12724 26608 12736
rect 26660 12724 26666 12776
rect 27062 12724 27068 12776
rect 27120 12764 27126 12776
rect 27801 12767 27859 12773
rect 27801 12764 27813 12767
rect 27120 12736 27813 12764
rect 27120 12724 27126 12736
rect 27801 12733 27813 12736
rect 27847 12733 27859 12767
rect 27801 12727 27859 12733
rect 24452 12668 25084 12696
rect 25225 12699 25283 12705
rect 24452 12656 24458 12668
rect 25225 12665 25237 12699
rect 25271 12696 25283 12699
rect 28350 12696 28356 12708
rect 25271 12668 28356 12696
rect 25271 12665 25283 12668
rect 25225 12659 25283 12665
rect 28350 12656 28356 12668
rect 28408 12656 28414 12708
rect 28534 12656 28540 12708
rect 28592 12696 28598 12708
rect 28905 12699 28963 12705
rect 28905 12696 28917 12699
rect 28592 12668 28917 12696
rect 28592 12656 28598 12668
rect 28905 12665 28917 12668
rect 28951 12665 28963 12699
rect 28905 12659 28963 12665
rect 29730 12656 29736 12708
rect 29788 12696 29794 12708
rect 30009 12699 30067 12705
rect 30009 12696 30021 12699
rect 29788 12668 30021 12696
rect 29788 12656 29794 12668
rect 30009 12665 30021 12668
rect 30055 12665 30067 12699
rect 30009 12659 30067 12665
rect 19392 12600 19656 12628
rect 19392 12588 19398 12600
rect 19978 12588 19984 12640
rect 20036 12628 20042 12640
rect 21453 12631 21511 12637
rect 21453 12628 21465 12631
rect 20036 12600 21465 12628
rect 20036 12588 20042 12600
rect 21453 12597 21465 12600
rect 21499 12597 21511 12631
rect 21453 12591 21511 12597
rect 24762 12588 24768 12640
rect 24820 12628 24826 12640
rect 25314 12628 25320 12640
rect 24820 12600 25320 12628
rect 24820 12588 24826 12600
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 28445 12631 28503 12637
rect 28445 12597 28457 12631
rect 28491 12628 28503 12631
rect 28626 12628 28632 12640
rect 28491 12600 28632 12628
rect 28491 12597 28503 12600
rect 28445 12591 28503 12597
rect 28626 12588 28632 12600
rect 28684 12588 28690 12640
rect 29362 12588 29368 12640
rect 29420 12628 29426 12640
rect 29457 12631 29515 12637
rect 29457 12628 29469 12631
rect 29420 12600 29469 12628
rect 29420 12588 29426 12600
rect 29457 12597 29469 12600
rect 29503 12628 29515 12631
rect 30561 12631 30619 12637
rect 30561 12628 30573 12631
rect 29503 12600 30573 12628
rect 29503 12597 29515 12600
rect 29457 12591 29515 12597
rect 30561 12597 30573 12600
rect 30607 12597 30619 12631
rect 30561 12591 30619 12597
rect 1104 12538 31832 12560
rect 1104 12486 4791 12538
rect 4843 12486 4855 12538
rect 4907 12486 4919 12538
rect 4971 12486 4983 12538
rect 5035 12486 5047 12538
rect 5099 12486 12473 12538
rect 12525 12486 12537 12538
rect 12589 12486 12601 12538
rect 12653 12486 12665 12538
rect 12717 12486 12729 12538
rect 12781 12486 20155 12538
rect 20207 12486 20219 12538
rect 20271 12486 20283 12538
rect 20335 12486 20347 12538
rect 20399 12486 20411 12538
rect 20463 12486 27837 12538
rect 27889 12486 27901 12538
rect 27953 12486 27965 12538
rect 28017 12486 28029 12538
rect 28081 12486 28093 12538
rect 28145 12486 31832 12538
rect 1104 12464 31832 12486
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 17034 12424 17040 12436
rect 16264 12396 17040 12424
rect 16264 12384 16270 12396
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 17678 12384 17684 12436
rect 17736 12424 17742 12436
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 17736 12396 18153 12424
rect 17736 12384 17742 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18141 12387 18199 12393
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 19981 12427 20039 12433
rect 19981 12424 19993 12427
rect 19944 12396 19993 12424
rect 19944 12384 19950 12396
rect 19981 12393 19993 12396
rect 20027 12393 20039 12427
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 19981 12387 20039 12393
rect 20088 12396 22845 12424
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 18785 12359 18843 12365
rect 18785 12356 18797 12359
rect 13780 12328 18797 12356
rect 13780 12316 13786 12328
rect 18785 12325 18797 12328
rect 18831 12325 18843 12359
rect 18785 12319 18843 12325
rect 18874 12316 18880 12368
rect 18932 12356 18938 12368
rect 20088 12356 20116 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 22833 12387 22891 12393
rect 23566 12384 23572 12436
rect 23624 12424 23630 12436
rect 24394 12424 24400 12436
rect 23624 12396 24400 12424
rect 23624 12384 23630 12396
rect 24394 12384 24400 12396
rect 24452 12384 24458 12436
rect 24670 12424 24676 12436
rect 24631 12396 24676 12424
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 24912 12396 25084 12424
rect 24912 12384 24918 12396
rect 18932 12328 20116 12356
rect 18932 12316 18938 12328
rect 22278 12316 22284 12368
rect 22336 12356 22342 12368
rect 22738 12356 22744 12368
rect 22336 12328 22744 12356
rect 22336 12316 22342 12328
rect 22738 12316 22744 12328
rect 22796 12316 22802 12368
rect 23661 12359 23719 12365
rect 23661 12325 23673 12359
rect 23707 12356 23719 12359
rect 24946 12356 24952 12368
rect 23707 12328 24952 12356
rect 23707 12325 23719 12328
rect 23661 12319 23719 12325
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 25056 12356 25084 12396
rect 25130 12384 25136 12436
rect 25188 12424 25194 12436
rect 26605 12427 26663 12433
rect 26605 12424 26617 12427
rect 25188 12396 26617 12424
rect 25188 12384 25194 12396
rect 26605 12393 26617 12396
rect 26651 12393 26663 12427
rect 26970 12424 26976 12436
rect 26605 12387 26663 12393
rect 26712 12396 26976 12424
rect 26712 12368 26740 12396
rect 26970 12384 26976 12396
rect 27028 12424 27034 12436
rect 27709 12427 27767 12433
rect 27709 12424 27721 12427
rect 27028 12396 27721 12424
rect 27028 12384 27034 12396
rect 27709 12393 27721 12396
rect 27755 12393 27767 12427
rect 27709 12387 27767 12393
rect 28166 12384 28172 12436
rect 28224 12424 28230 12436
rect 28442 12424 28448 12436
rect 28224 12396 28448 12424
rect 28224 12384 28230 12396
rect 28442 12384 28448 12396
rect 28500 12384 28506 12436
rect 31294 12424 31300 12436
rect 31255 12396 31300 12424
rect 31294 12384 31300 12396
rect 31352 12384 31358 12436
rect 25314 12356 25320 12368
rect 25056 12328 25320 12356
rect 25314 12316 25320 12328
rect 25372 12316 25378 12368
rect 25866 12316 25872 12368
rect 25924 12356 25930 12368
rect 26053 12359 26111 12365
rect 26053 12356 26065 12359
rect 25924 12328 26065 12356
rect 25924 12316 25930 12328
rect 26053 12325 26065 12328
rect 26099 12325 26111 12359
rect 26053 12319 26111 12325
rect 26694 12316 26700 12368
rect 26752 12316 26758 12368
rect 28074 12316 28080 12368
rect 28132 12356 28138 12368
rect 28810 12356 28816 12368
rect 28132 12328 28816 12356
rect 28132 12316 28138 12328
rect 28810 12316 28816 12328
rect 28868 12316 28874 12368
rect 13538 12248 13544 12300
rect 13596 12288 13602 12300
rect 17402 12288 17408 12300
rect 13596 12260 17408 12288
rect 13596 12248 13602 12260
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 18966 12288 18972 12300
rect 17880 12260 18972 12288
rect 17034 12220 17040 12232
rect 16995 12192 17040 12220
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 14918 12112 14924 12164
rect 14976 12152 14982 12164
rect 17880 12152 17908 12260
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12288 20959 12291
rect 27246 12288 27252 12300
rect 20947 12260 23704 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 23676 12232 23704 12260
rect 25424 12260 27252 12288
rect 18046 12220 18052 12232
rect 18007 12192 18052 12220
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 18322 12220 18328 12232
rect 18279 12192 18328 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 18322 12180 18328 12192
rect 18380 12180 18386 12232
rect 18414 12180 18420 12232
rect 18472 12220 18478 12232
rect 18877 12223 18935 12229
rect 18877 12220 18889 12223
rect 18472 12192 18889 12220
rect 18472 12180 18478 12192
rect 18877 12189 18889 12192
rect 18923 12189 18935 12223
rect 19978 12220 19984 12232
rect 19891 12192 19984 12220
rect 18877 12183 18935 12189
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20070 12180 20076 12232
rect 20128 12220 20134 12232
rect 20165 12223 20223 12229
rect 20165 12220 20177 12223
rect 20128 12192 20177 12220
rect 20128 12180 20134 12192
rect 20165 12189 20177 12192
rect 20211 12189 20223 12223
rect 20622 12220 20628 12232
rect 20583 12192 20628 12220
rect 20165 12183 20223 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22796 12192 22845 12220
rect 22796 12180 22802 12192
rect 22833 12189 22845 12192
rect 22879 12220 22891 12223
rect 23014 12220 23020 12232
rect 22879 12192 23020 12220
rect 22879 12189 22891 12192
rect 22833 12183 22891 12189
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 23109 12223 23167 12229
rect 23109 12189 23121 12223
rect 23155 12220 23167 12223
rect 23382 12220 23388 12232
rect 23155 12192 23388 12220
rect 23155 12189 23167 12192
rect 23109 12183 23167 12189
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 14976 12124 17908 12152
rect 18064 12152 18092 12180
rect 19996 12152 20024 12180
rect 22462 12152 22468 12164
rect 18064 12124 20024 12152
rect 22126 12124 22468 12152
rect 14976 12112 14982 12124
rect 22462 12112 22468 12124
rect 22520 12112 22526 12164
rect 23584 12152 23612 12183
rect 23658 12180 23664 12232
rect 23716 12180 23722 12232
rect 24762 12220 24768 12232
rect 24723 12192 24768 12220
rect 24762 12180 24768 12192
rect 24820 12180 24826 12232
rect 24854 12180 24860 12232
rect 24912 12220 24918 12232
rect 25424 12229 25452 12260
rect 27246 12248 27252 12260
rect 27304 12248 27310 12300
rect 28350 12248 28356 12300
rect 28408 12288 28414 12300
rect 29270 12288 29276 12300
rect 28408 12260 29276 12288
rect 28408 12248 28414 12260
rect 29270 12248 29276 12260
rect 29328 12248 29334 12300
rect 25225 12223 25283 12229
rect 25225 12220 25237 12223
rect 24912 12192 25237 12220
rect 24912 12180 24918 12192
rect 25225 12189 25237 12192
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12189 25467 12223
rect 25409 12183 25467 12189
rect 25869 12223 25927 12229
rect 25869 12189 25881 12223
rect 25915 12220 25927 12223
rect 26050 12220 26056 12232
rect 25915 12192 26056 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 26050 12180 26056 12192
rect 26108 12180 26114 12232
rect 26326 12180 26332 12232
rect 26384 12220 26390 12232
rect 26697 12223 26755 12229
rect 26697 12220 26709 12223
rect 26384 12192 26709 12220
rect 26384 12180 26390 12192
rect 26697 12189 26709 12192
rect 26743 12189 26755 12223
rect 26697 12183 26755 12189
rect 26878 12180 26884 12232
rect 26936 12220 26942 12232
rect 28718 12220 28724 12232
rect 26936 12192 28724 12220
rect 26936 12180 26942 12192
rect 28718 12180 28724 12192
rect 28776 12220 28782 12232
rect 30466 12220 30472 12232
rect 28776 12192 30472 12220
rect 28776 12180 28782 12192
rect 30466 12180 30472 12192
rect 30524 12180 30530 12232
rect 24780 12152 24808 12180
rect 25498 12152 25504 12164
rect 23584 12124 24808 12152
rect 25332 12124 25504 12152
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17589 12087 17647 12093
rect 17589 12084 17601 12087
rect 17368 12056 17601 12084
rect 17368 12044 17374 12056
rect 17589 12053 17601 12056
rect 17635 12084 17647 12087
rect 17678 12084 17684 12096
rect 17635 12056 17684 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 19797 12087 19855 12093
rect 19797 12084 19809 12087
rect 18288 12056 19809 12084
rect 18288 12044 18294 12056
rect 19797 12053 19809 12056
rect 19843 12053 19855 12087
rect 19797 12047 19855 12053
rect 19886 12044 19892 12096
rect 19944 12084 19950 12096
rect 21726 12084 21732 12096
rect 19944 12056 21732 12084
rect 19944 12044 19950 12056
rect 21726 12044 21732 12056
rect 21784 12044 21790 12096
rect 22370 12084 22376 12096
rect 22283 12056 22376 12084
rect 22370 12044 22376 12056
rect 22428 12084 22434 12096
rect 23017 12087 23075 12093
rect 23017 12084 23029 12087
rect 22428 12056 23029 12084
rect 22428 12044 22434 12056
rect 23017 12053 23029 12056
rect 23063 12084 23075 12087
rect 24578 12084 24584 12096
rect 23063 12056 24584 12084
rect 23063 12053 23075 12056
rect 23017 12047 23075 12053
rect 24578 12044 24584 12056
rect 24636 12044 24642 12096
rect 24946 12044 24952 12096
rect 25004 12084 25010 12096
rect 25332 12093 25360 12124
rect 25498 12112 25504 12124
rect 25556 12152 25562 12164
rect 29362 12152 29368 12164
rect 25556 12124 29368 12152
rect 25556 12112 25562 12124
rect 29362 12112 29368 12124
rect 29420 12112 29426 12164
rect 25317 12087 25375 12093
rect 25317 12084 25329 12087
rect 25004 12056 25329 12084
rect 25004 12044 25010 12056
rect 25317 12053 25329 12056
rect 25363 12053 25375 12087
rect 27154 12084 27160 12096
rect 27115 12056 27160 12084
rect 25317 12047 25375 12053
rect 27154 12044 27160 12056
rect 27212 12044 27218 12096
rect 27982 12044 27988 12096
rect 28040 12084 28046 12096
rect 28261 12087 28319 12093
rect 28261 12084 28273 12087
rect 28040 12056 28273 12084
rect 28040 12044 28046 12056
rect 28261 12053 28273 12056
rect 28307 12053 28319 12087
rect 28810 12084 28816 12096
rect 28771 12056 28816 12084
rect 28261 12047 28319 12053
rect 28810 12044 28816 12056
rect 28868 12044 28874 12096
rect 29825 12087 29883 12093
rect 29825 12053 29837 12087
rect 29871 12084 29883 12087
rect 30190 12084 30196 12096
rect 29871 12056 30196 12084
rect 29871 12053 29883 12056
rect 29825 12047 29883 12053
rect 30190 12044 30196 12056
rect 30248 12044 30254 12096
rect 30377 12087 30435 12093
rect 30377 12053 30389 12087
rect 30423 12084 30435 12087
rect 30650 12084 30656 12096
rect 30423 12056 30656 12084
rect 30423 12053 30435 12056
rect 30377 12047 30435 12053
rect 30650 12044 30656 12056
rect 30708 12044 30714 12096
rect 1104 11994 31992 12016
rect 1104 11942 8632 11994
rect 8684 11942 8696 11994
rect 8748 11942 8760 11994
rect 8812 11942 8824 11994
rect 8876 11942 8888 11994
rect 8940 11942 16314 11994
rect 16366 11942 16378 11994
rect 16430 11942 16442 11994
rect 16494 11942 16506 11994
rect 16558 11942 16570 11994
rect 16622 11942 23996 11994
rect 24048 11942 24060 11994
rect 24112 11942 24124 11994
rect 24176 11942 24188 11994
rect 24240 11942 24252 11994
rect 24304 11942 31678 11994
rect 31730 11942 31742 11994
rect 31794 11942 31806 11994
rect 31858 11942 31870 11994
rect 31922 11942 31934 11994
rect 31986 11942 31992 11994
rect 1104 11920 31992 11942
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 17770 11880 17776 11892
rect 9640 11852 17776 11880
rect 9640 11840 9646 11852
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 18322 11880 18328 11892
rect 17880 11852 18328 11880
rect 17034 11772 17040 11824
rect 17092 11812 17098 11824
rect 17313 11815 17371 11821
rect 17313 11812 17325 11815
rect 17092 11784 17325 11812
rect 17092 11772 17098 11784
rect 17313 11781 17325 11784
rect 17359 11812 17371 11815
rect 17880 11812 17908 11852
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 19518 11880 19524 11892
rect 19479 11852 19524 11880
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 22002 11880 22008 11892
rect 20272 11852 22008 11880
rect 17359 11784 17908 11812
rect 17359 11781 17371 11784
rect 17313 11775 17371 11781
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 18012 11784 19472 11812
rect 18012 11772 18018 11784
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 18230 11744 18236 11756
rect 15988 11716 18236 11744
rect 15988 11704 15994 11716
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 19444 11753 19472 11784
rect 18969 11747 19027 11753
rect 18969 11744 18981 11747
rect 18380 11716 18981 11744
rect 18380 11704 18386 11716
rect 18969 11713 18981 11716
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 17586 11636 17592 11688
rect 17644 11676 17650 11688
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 17644 11648 18889 11676
rect 17644 11636 17650 11648
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18984 11676 19012 11707
rect 19886 11676 19892 11688
rect 18984 11648 19892 11676
rect 18877 11639 18935 11645
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 16942 11568 16948 11620
rect 17000 11608 17006 11620
rect 20272 11608 20300 11852
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 22173 11883 22231 11889
rect 22173 11849 22185 11883
rect 22219 11880 22231 11883
rect 22738 11880 22744 11892
rect 22219 11852 22744 11880
rect 22219 11849 22231 11852
rect 22173 11843 22231 11849
rect 22738 11840 22744 11852
rect 22796 11840 22802 11892
rect 22922 11880 22928 11892
rect 22883 11852 22928 11880
rect 22922 11840 22928 11852
rect 22980 11840 22986 11892
rect 23566 11880 23572 11892
rect 23527 11852 23572 11880
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 23842 11840 23848 11892
rect 23900 11880 23906 11892
rect 24213 11883 24271 11889
rect 24213 11880 24225 11883
rect 23900 11852 24225 11880
rect 23900 11840 23906 11852
rect 24213 11849 24225 11852
rect 24259 11849 24271 11883
rect 24213 11843 24271 11849
rect 24857 11883 24915 11889
rect 24857 11849 24869 11883
rect 24903 11880 24915 11883
rect 25130 11880 25136 11892
rect 24903 11852 25136 11880
rect 24903 11849 24915 11852
rect 24857 11843 24915 11849
rect 25130 11840 25136 11852
rect 25188 11840 25194 11892
rect 26142 11840 26148 11892
rect 26200 11880 26206 11892
rect 26237 11883 26295 11889
rect 26237 11880 26249 11883
rect 26200 11852 26249 11880
rect 26200 11840 26206 11852
rect 26237 11849 26249 11852
rect 26283 11849 26295 11883
rect 28074 11880 28080 11892
rect 26237 11843 26295 11849
rect 26712 11852 28080 11880
rect 22370 11812 22376 11824
rect 20364 11784 21864 11812
rect 22331 11784 22376 11812
rect 20364 11753 20392 11784
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20956 11716 21005 11744
rect 20956 11704 20962 11716
rect 20993 11713 21005 11716
rect 21039 11713 21051 11747
rect 21266 11744 21272 11756
rect 20993 11707 21051 11713
rect 21100 11716 21272 11744
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 21100 11676 21128 11716
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 20772 11648 21128 11676
rect 20772 11636 20778 11648
rect 21174 11636 21180 11688
rect 21232 11676 21238 11688
rect 21836 11676 21864 11784
rect 22370 11772 22376 11784
rect 22428 11772 22434 11824
rect 26712 11812 26740 11852
rect 28074 11840 28080 11852
rect 28132 11840 28138 11892
rect 28258 11840 28264 11892
rect 28316 11880 28322 11892
rect 28813 11883 28871 11889
rect 28813 11880 28825 11883
rect 28316 11852 28825 11880
rect 28316 11840 28322 11852
rect 28813 11849 28825 11852
rect 28859 11849 28871 11883
rect 28813 11843 28871 11849
rect 27522 11812 27528 11824
rect 23032 11784 24348 11812
rect 21910 11704 21916 11756
rect 21968 11744 21974 11756
rect 23032 11753 23060 11784
rect 23584 11756 23612 11784
rect 23017 11747 23075 11753
rect 21968 11716 22968 11744
rect 21968 11704 21974 11716
rect 22940 11676 22968 11716
rect 23017 11713 23029 11747
rect 23063 11713 23075 11747
rect 23017 11707 23075 11713
rect 23566 11704 23572 11756
rect 23624 11704 23630 11756
rect 23661 11747 23719 11753
rect 23661 11713 23673 11747
rect 23707 11744 23719 11747
rect 23842 11744 23848 11756
rect 23707 11716 23848 11744
rect 23707 11713 23719 11716
rect 23661 11707 23719 11713
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 24320 11753 24348 11784
rect 24872 11784 26740 11812
rect 26804 11784 27528 11812
rect 24872 11756 24900 11784
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11744 24363 11747
rect 24762 11744 24768 11756
rect 24351 11716 24768 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 24762 11704 24768 11716
rect 24820 11704 24826 11756
rect 24854 11704 24860 11756
rect 24912 11704 24918 11756
rect 24949 11747 25007 11753
rect 24949 11713 24961 11747
rect 24995 11744 25007 11747
rect 25038 11744 25044 11756
rect 24995 11716 25044 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11744 25743 11747
rect 25866 11744 25872 11756
rect 25731 11716 25872 11744
rect 25731 11713 25743 11716
rect 25685 11707 25743 11713
rect 25866 11704 25872 11716
rect 25924 11744 25930 11756
rect 26326 11744 26332 11756
rect 25924 11716 26332 11744
rect 25924 11704 25930 11716
rect 26326 11704 26332 11716
rect 26384 11744 26390 11756
rect 26804 11744 26832 11784
rect 27522 11772 27528 11784
rect 27580 11772 27586 11824
rect 27614 11772 27620 11824
rect 27672 11812 27678 11824
rect 29917 11815 29975 11821
rect 29917 11812 29929 11815
rect 27672 11784 29929 11812
rect 27672 11772 27678 11784
rect 29917 11781 29929 11784
rect 29963 11812 29975 11815
rect 30466 11812 30472 11824
rect 29963 11784 30472 11812
rect 29963 11781 29975 11784
rect 29917 11775 29975 11781
rect 30466 11772 30472 11784
rect 30524 11772 30530 11824
rect 31294 11744 31300 11756
rect 26384 11716 26832 11744
rect 31255 11716 31300 11744
rect 26384 11704 26390 11716
rect 31294 11704 31300 11716
rect 31352 11704 31358 11756
rect 25593 11679 25651 11685
rect 25593 11676 25605 11679
rect 21232 11648 21277 11676
rect 21836 11648 22232 11676
rect 22940 11648 25605 11676
rect 21232 11636 21238 11648
rect 17000 11580 20300 11608
rect 20349 11611 20407 11617
rect 17000 11568 17006 11580
rect 20349 11577 20361 11611
rect 20395 11608 20407 11611
rect 22094 11608 22100 11620
rect 20395 11580 22100 11608
rect 20395 11577 20407 11580
rect 20349 11571 20407 11577
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 17310 11540 17316 11552
rect 15160 11512 17316 11540
rect 15160 11500 15166 11512
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 20714 11540 20720 11552
rect 17460 11512 20720 11540
rect 17460 11500 17466 11512
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 20809 11543 20867 11549
rect 20809 11509 20821 11543
rect 20855 11540 20867 11543
rect 21082 11540 21088 11552
rect 20855 11512 21088 11540
rect 20855 11509 20867 11512
rect 20809 11503 20867 11509
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 22204 11549 22232 11648
rect 25593 11645 25605 11648
rect 25639 11645 25651 11679
rect 29454 11676 29460 11688
rect 25593 11639 25651 11645
rect 25700 11648 29460 11676
rect 24578 11568 24584 11620
rect 24636 11608 24642 11620
rect 25700 11608 25728 11648
rect 29454 11636 29460 11648
rect 29512 11636 29518 11688
rect 24636 11580 25728 11608
rect 24636 11568 24642 11580
rect 26786 11568 26792 11620
rect 26844 11608 26850 11620
rect 27157 11611 27215 11617
rect 27157 11608 27169 11611
rect 26844 11580 27169 11608
rect 26844 11568 26850 11580
rect 27157 11577 27169 11580
rect 27203 11608 27215 11611
rect 27982 11608 27988 11620
rect 27203 11580 27988 11608
rect 27203 11577 27215 11580
rect 27157 11571 27215 11577
rect 27982 11568 27988 11580
rect 28040 11608 28046 11620
rect 28261 11611 28319 11617
rect 28261 11608 28273 11611
rect 28040 11580 28273 11608
rect 28040 11568 28046 11580
rect 28261 11577 28273 11580
rect 28307 11577 28319 11611
rect 28261 11571 28319 11577
rect 22189 11543 22247 11549
rect 22189 11509 22201 11543
rect 22235 11540 22247 11543
rect 23382 11540 23388 11552
rect 22235 11512 23388 11540
rect 22235 11509 22247 11512
rect 22189 11503 22247 11509
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 27706 11540 27712 11552
rect 27667 11512 27712 11540
rect 27706 11500 27712 11512
rect 27764 11500 27770 11552
rect 29362 11540 29368 11552
rect 29323 11512 29368 11540
rect 29362 11500 29368 11512
rect 29420 11500 29426 11552
rect 30374 11500 30380 11552
rect 30432 11540 30438 11552
rect 30469 11543 30527 11549
rect 30469 11540 30481 11543
rect 30432 11512 30481 11540
rect 30432 11500 30438 11512
rect 30469 11509 30481 11512
rect 30515 11509 30527 11543
rect 30469 11503 30527 11509
rect 1104 11450 31832 11472
rect 1104 11398 4791 11450
rect 4843 11398 4855 11450
rect 4907 11398 4919 11450
rect 4971 11398 4983 11450
rect 5035 11398 5047 11450
rect 5099 11398 12473 11450
rect 12525 11398 12537 11450
rect 12589 11398 12601 11450
rect 12653 11398 12665 11450
rect 12717 11398 12729 11450
rect 12781 11398 20155 11450
rect 20207 11398 20219 11450
rect 20271 11398 20283 11450
rect 20335 11398 20347 11450
rect 20399 11398 20411 11450
rect 20463 11398 27837 11450
rect 27889 11398 27901 11450
rect 27953 11398 27965 11450
rect 28017 11398 28029 11450
rect 28081 11398 28093 11450
rect 28145 11398 31832 11450
rect 1104 11376 31832 11398
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 20717 11339 20775 11345
rect 20717 11336 20729 11339
rect 16172 11308 20729 11336
rect 16172 11296 16178 11308
rect 20717 11305 20729 11308
rect 20763 11305 20775 11339
rect 21634 11336 21640 11348
rect 21595 11308 21640 11336
rect 20717 11299 20775 11305
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 22186 11336 22192 11348
rect 22147 11308 22192 11336
rect 22186 11296 22192 11308
rect 22244 11296 22250 11348
rect 22833 11339 22891 11345
rect 22833 11305 22845 11339
rect 22879 11336 22891 11339
rect 23290 11336 23296 11348
rect 22879 11308 23296 11336
rect 22879 11305 22891 11308
rect 22833 11299 22891 11305
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 23474 11336 23480 11348
rect 23435 11308 23480 11336
rect 23474 11296 23480 11308
rect 23532 11296 23538 11348
rect 26602 11296 26608 11348
rect 26660 11336 26666 11348
rect 26789 11339 26847 11345
rect 26789 11336 26801 11339
rect 26660 11308 26801 11336
rect 26660 11296 26666 11308
rect 26789 11305 26801 11308
rect 26835 11336 26847 11339
rect 26878 11336 26884 11348
rect 26835 11308 26884 11336
rect 26835 11305 26847 11308
rect 26789 11299 26847 11305
rect 26878 11296 26884 11308
rect 26936 11296 26942 11348
rect 27982 11296 27988 11348
rect 28040 11336 28046 11348
rect 28537 11339 28595 11345
rect 28537 11336 28549 11339
rect 28040 11308 28549 11336
rect 28040 11296 28046 11308
rect 28537 11305 28549 11308
rect 28583 11336 28595 11339
rect 29638 11336 29644 11348
rect 28583 11308 29644 11336
rect 28583 11305 28595 11308
rect 28537 11299 28595 11305
rect 29638 11296 29644 11308
rect 29696 11296 29702 11348
rect 31294 11336 31300 11348
rect 31255 11308 31300 11336
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 19797 11271 19855 11277
rect 19797 11237 19809 11271
rect 19843 11268 19855 11271
rect 21818 11268 21824 11280
rect 19843 11240 21824 11268
rect 19843 11237 19855 11240
rect 19797 11231 19855 11237
rect 21818 11228 21824 11240
rect 21876 11228 21882 11280
rect 22002 11228 22008 11280
rect 22060 11268 22066 11280
rect 28166 11268 28172 11280
rect 22060 11240 28172 11268
rect 22060 11228 22066 11240
rect 28166 11228 28172 11240
rect 28224 11228 28230 11280
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 19242 11200 19248 11212
rect 17368 11172 19248 11200
rect 17368 11160 17374 11172
rect 19242 11160 19248 11172
rect 19300 11200 19306 11212
rect 19300 11172 20208 11200
rect 19300 11160 19306 11172
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11132 19763 11135
rect 19886 11132 19892 11144
rect 19751 11104 19892 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20180 11132 20208 11172
rect 20898 11160 20904 11212
rect 20956 11200 20962 11212
rect 24578 11200 24584 11212
rect 20956 11172 24584 11200
rect 20956 11160 20962 11172
rect 24578 11160 24584 11172
rect 24636 11160 24642 11212
rect 27614 11160 27620 11212
rect 27672 11200 27678 11212
rect 30377 11203 30435 11209
rect 30377 11200 30389 11203
rect 27672 11172 30389 11200
rect 27672 11160 27678 11172
rect 30377 11169 30389 11172
rect 30423 11169 30435 11203
rect 30377 11163 30435 11169
rect 20717 11135 20775 11141
rect 20717 11132 20729 11135
rect 20180 11104 20729 11132
rect 20717 11101 20729 11104
rect 20763 11101 20775 11135
rect 20717 11095 20775 11101
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 21450 11132 21456 11144
rect 20864 11104 20909 11132
rect 21411 11104 21456 11132
rect 20864 11092 20870 11104
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 22002 11092 22008 11144
rect 22060 11132 22066 11144
rect 22097 11135 22155 11141
rect 22097 11132 22109 11135
rect 22060 11104 22109 11132
rect 22060 11092 22066 11104
rect 22097 11101 22109 11104
rect 22143 11132 22155 11135
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 22143 11104 22753 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 22741 11101 22753 11104
rect 22787 11132 22799 11135
rect 23566 11132 23572 11144
rect 22787 11104 23572 11132
rect 22787 11101 22799 11104
rect 22741 11095 22799 11101
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 27433 11135 27491 11141
rect 27433 11101 27445 11135
rect 27479 11132 27491 11135
rect 28258 11132 28264 11144
rect 27479 11104 28264 11132
rect 27479 11101 27491 11104
rect 27433 11095 27491 11101
rect 28258 11092 28264 11104
rect 28316 11092 28322 11144
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 18877 11067 18935 11073
rect 18877 11064 18889 11067
rect 13504 11036 18889 11064
rect 13504 11024 13510 11036
rect 18877 11033 18889 11036
rect 18923 11064 18935 11067
rect 20898 11064 20904 11076
rect 18923 11036 20904 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 20993 11067 21051 11073
rect 20993 11033 21005 11067
rect 21039 11064 21051 11067
rect 22830 11064 22836 11076
rect 21039 11036 22836 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 4154 10956 4160 11008
rect 4212 10996 4218 11008
rect 9490 10996 9496 11008
rect 4212 10968 9496 10996
rect 4212 10956 4218 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 19150 10956 19156 11008
rect 19208 10996 19214 11008
rect 20070 10996 20076 11008
rect 19208 10968 20076 10996
rect 19208 10956 19214 10968
rect 20070 10956 20076 10968
rect 20128 10996 20134 11008
rect 21008 10996 21036 11027
rect 22830 11024 22836 11036
rect 22888 11024 22894 11076
rect 24670 11064 24676 11076
rect 24631 11036 24676 11064
rect 24670 11024 24676 11036
rect 24728 11024 24734 11076
rect 25685 11067 25743 11073
rect 25685 11033 25697 11067
rect 25731 11064 25743 11067
rect 27522 11064 27528 11076
rect 25731 11036 27528 11064
rect 25731 11033 25743 11036
rect 25685 11027 25743 11033
rect 27522 11024 27528 11036
rect 27580 11064 27586 11076
rect 27982 11064 27988 11076
rect 27580 11036 27988 11064
rect 27580 11024 27586 11036
rect 27982 11024 27988 11036
rect 28040 11024 28046 11076
rect 20128 10968 21036 10996
rect 20128 10956 20134 10968
rect 21082 10956 21088 11008
rect 21140 10996 21146 11008
rect 25225 10999 25283 11005
rect 25225 10996 25237 10999
rect 21140 10968 25237 10996
rect 21140 10956 21146 10968
rect 25225 10965 25237 10968
rect 25271 10996 25283 10999
rect 25498 10996 25504 11008
rect 25271 10968 25504 10996
rect 25271 10965 25283 10968
rect 25225 10959 25283 10965
rect 25498 10956 25504 10968
rect 25556 10996 25562 11008
rect 25774 10996 25780 11008
rect 25556 10968 25780 10996
rect 25556 10956 25562 10968
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 26326 10996 26332 11008
rect 26239 10968 26332 10996
rect 26326 10956 26332 10968
rect 26384 10996 26390 11008
rect 27062 10996 27068 11008
rect 26384 10968 27068 10996
rect 26384 10956 26390 10968
rect 27062 10956 27068 10968
rect 27120 10956 27126 11008
rect 27246 10956 27252 11008
rect 27304 10996 27310 11008
rect 27706 10996 27712 11008
rect 27304 10968 27712 10996
rect 27304 10956 27310 10968
rect 27706 10956 27712 10968
rect 27764 10996 27770 11008
rect 27893 10999 27951 11005
rect 27893 10996 27905 10999
rect 27764 10968 27905 10996
rect 27764 10956 27770 10968
rect 27893 10965 27905 10968
rect 27939 10965 27951 10999
rect 27893 10959 27951 10965
rect 28810 10956 28816 11008
rect 28868 10996 28874 11008
rect 28997 10999 29055 11005
rect 28997 10996 29009 10999
rect 28868 10968 29009 10996
rect 28868 10956 28874 10968
rect 28997 10965 29009 10968
rect 29043 10965 29055 10999
rect 29730 10996 29736 11008
rect 29691 10968 29736 10996
rect 28997 10959 29055 10965
rect 29730 10956 29736 10968
rect 29788 10956 29794 11008
rect 1104 10906 31992 10928
rect 1104 10854 8632 10906
rect 8684 10854 8696 10906
rect 8748 10854 8760 10906
rect 8812 10854 8824 10906
rect 8876 10854 8888 10906
rect 8940 10854 16314 10906
rect 16366 10854 16378 10906
rect 16430 10854 16442 10906
rect 16494 10854 16506 10906
rect 16558 10854 16570 10906
rect 16622 10854 23996 10906
rect 24048 10854 24060 10906
rect 24112 10854 24124 10906
rect 24176 10854 24188 10906
rect 24240 10854 24252 10906
rect 24304 10854 31678 10906
rect 31730 10854 31742 10906
rect 31794 10854 31806 10906
rect 31858 10854 31870 10906
rect 31922 10854 31934 10906
rect 31986 10854 31992 10906
rect 1104 10832 31992 10854
rect 19613 10795 19671 10801
rect 19613 10761 19625 10795
rect 19659 10792 19671 10795
rect 19886 10792 19892 10804
rect 19659 10764 19892 10792
rect 19659 10761 19671 10764
rect 19613 10755 19671 10761
rect 19886 10752 19892 10764
rect 19944 10752 19950 10804
rect 20165 10795 20223 10801
rect 20165 10761 20177 10795
rect 20211 10792 20223 10795
rect 20530 10792 20536 10804
rect 20211 10764 20536 10792
rect 20211 10761 20223 10764
rect 20165 10755 20223 10761
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 20898 10792 20904 10804
rect 20859 10764 20904 10792
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 22097 10795 22155 10801
rect 22097 10761 22109 10795
rect 22143 10792 22155 10795
rect 22554 10792 22560 10804
rect 22143 10764 22560 10792
rect 22143 10761 22155 10764
rect 22097 10755 22155 10761
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 22646 10752 22652 10804
rect 22704 10792 22710 10804
rect 22741 10795 22799 10801
rect 22741 10792 22753 10795
rect 22704 10764 22753 10792
rect 22704 10752 22710 10764
rect 22741 10761 22753 10764
rect 22787 10761 22799 10795
rect 22741 10755 22799 10761
rect 23198 10752 23204 10804
rect 23256 10792 23262 10804
rect 23256 10764 24624 10792
rect 23256 10752 23262 10764
rect 11514 10684 11520 10736
rect 11572 10724 11578 10736
rect 11572 10696 22048 10724
rect 11572 10684 11578 10696
rect 22020 10668 22048 10696
rect 22462 10684 22468 10736
rect 22520 10724 22526 10736
rect 23385 10727 23443 10733
rect 23385 10724 23397 10727
rect 22520 10696 23397 10724
rect 22520 10684 22526 10696
rect 23385 10693 23397 10696
rect 23431 10693 23443 10727
rect 24596 10724 24624 10764
rect 24670 10752 24676 10804
rect 24728 10792 24734 10804
rect 29365 10795 29423 10801
rect 29365 10792 29377 10795
rect 24728 10764 29377 10792
rect 24728 10752 24734 10764
rect 29365 10761 29377 10764
rect 29411 10761 29423 10795
rect 31018 10792 31024 10804
rect 30979 10764 31024 10792
rect 29365 10755 29423 10761
rect 31018 10752 31024 10764
rect 31076 10752 31082 10804
rect 28813 10727 28871 10733
rect 28813 10724 28825 10727
rect 24596 10696 28825 10724
rect 23385 10687 23443 10693
rect 28813 10693 28825 10696
rect 28859 10724 28871 10727
rect 30469 10727 30527 10733
rect 30469 10724 30481 10727
rect 28859 10696 30481 10724
rect 28859 10693 28871 10696
rect 28813 10687 28871 10693
rect 30469 10693 30481 10696
rect 30515 10724 30527 10727
rect 32582 10724 32588 10736
rect 30515 10696 32588 10724
rect 30515 10693 30527 10696
rect 30469 10687 30527 10693
rect 32582 10684 32588 10696
rect 32640 10684 32646 10736
rect 20070 10656 20076 10668
rect 20031 10628 20076 10656
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10625 20315 10659
rect 20714 10656 20720 10668
rect 20675 10628 20720 10656
rect 20257 10619 20315 10625
rect 1578 10588 1584 10600
rect 1539 10560 1584 10588
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 20272 10588 20300 10619
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 20898 10656 20904 10668
rect 20859 10628 20904 10656
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 22002 10656 22008 10668
rect 21963 10628 22008 10656
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10656 22707 10659
rect 23477 10659 23535 10665
rect 23477 10656 23489 10659
rect 22695 10628 23489 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 23477 10625 23489 10628
rect 23523 10656 23535 10659
rect 23658 10656 23664 10668
rect 23523 10628 23664 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 23658 10616 23664 10628
rect 23716 10616 23722 10668
rect 24578 10656 24584 10668
rect 24539 10628 24584 10656
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 25130 10616 25136 10668
rect 25188 10656 25194 10668
rect 26326 10656 26332 10668
rect 25188 10628 26332 10656
rect 25188 10616 25194 10628
rect 26326 10616 26332 10628
rect 26384 10616 26390 10668
rect 28994 10588 29000 10600
rect 20272 10560 29000 10588
rect 28994 10548 29000 10560
rect 29052 10548 29058 10600
rect 29914 10588 29920 10600
rect 29875 10560 29920 10588
rect 29914 10548 29920 10560
rect 29972 10548 29978 10600
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 10318 10520 10324 10532
rect 5316 10492 10324 10520
rect 5316 10480 5322 10492
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 22186 10520 22192 10532
rect 20772 10492 22192 10520
rect 20772 10480 20778 10492
rect 22186 10480 22192 10492
rect 22244 10480 22250 10532
rect 22278 10480 22284 10532
rect 22336 10520 22342 10532
rect 23198 10520 23204 10532
rect 22336 10492 23204 10520
rect 22336 10480 22342 10492
rect 23198 10480 23204 10492
rect 23256 10480 23262 10532
rect 26237 10523 26295 10529
rect 26237 10520 26249 10523
rect 23308 10492 26249 10520
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 20806 10452 20812 10464
rect 17736 10424 20812 10452
rect 17736 10412 17742 10424
rect 20806 10412 20812 10424
rect 20864 10452 20870 10464
rect 21082 10452 21088 10464
rect 20864 10424 21088 10452
rect 20864 10412 20870 10424
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 21453 10455 21511 10461
rect 21453 10421 21465 10455
rect 21499 10452 21511 10455
rect 21542 10452 21548 10464
rect 21499 10424 21548 10452
rect 21499 10421 21511 10424
rect 21453 10415 21511 10421
rect 21542 10412 21548 10424
rect 21600 10452 21606 10464
rect 23308 10452 23336 10492
rect 26237 10489 26249 10492
rect 26283 10489 26295 10523
rect 28261 10523 28319 10529
rect 28261 10520 28273 10523
rect 26237 10483 26295 10489
rect 27172 10492 28273 10520
rect 21600 10424 23336 10452
rect 24029 10455 24087 10461
rect 21600 10412 21606 10424
rect 24029 10421 24041 10455
rect 24075 10452 24087 10455
rect 24302 10452 24308 10464
rect 24075 10424 24308 10452
rect 24075 10421 24087 10424
rect 24029 10415 24087 10421
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 25130 10412 25136 10464
rect 25188 10452 25194 10464
rect 25317 10455 25375 10461
rect 25317 10452 25329 10455
rect 25188 10424 25329 10452
rect 25188 10412 25194 10424
rect 25317 10421 25329 10424
rect 25363 10421 25375 10455
rect 25317 10415 25375 10421
rect 26602 10412 26608 10464
rect 26660 10452 26666 10464
rect 27172 10461 27200 10492
rect 28261 10489 28273 10492
rect 28307 10520 28319 10523
rect 28350 10520 28356 10532
rect 28307 10492 28356 10520
rect 28307 10489 28319 10492
rect 28261 10483 28319 10489
rect 28350 10480 28356 10492
rect 28408 10480 28414 10532
rect 31386 10520 31392 10532
rect 28966 10492 31392 10520
rect 27157 10455 27215 10461
rect 27157 10452 27169 10455
rect 26660 10424 27169 10452
rect 26660 10412 26666 10424
rect 27157 10421 27169 10424
rect 27203 10421 27215 10455
rect 27706 10452 27712 10464
rect 27667 10424 27712 10452
rect 27157 10415 27215 10421
rect 27706 10412 27712 10424
rect 27764 10452 27770 10464
rect 28966 10452 28994 10492
rect 31386 10480 31392 10492
rect 31444 10480 31450 10532
rect 27764 10424 28994 10452
rect 27764 10412 27770 10424
rect 1104 10362 31832 10384
rect 1104 10310 4791 10362
rect 4843 10310 4855 10362
rect 4907 10310 4919 10362
rect 4971 10310 4983 10362
rect 5035 10310 5047 10362
rect 5099 10310 12473 10362
rect 12525 10310 12537 10362
rect 12589 10310 12601 10362
rect 12653 10310 12665 10362
rect 12717 10310 12729 10362
rect 12781 10310 20155 10362
rect 20207 10310 20219 10362
rect 20271 10310 20283 10362
rect 20335 10310 20347 10362
rect 20399 10310 20411 10362
rect 20463 10310 27837 10362
rect 27889 10310 27901 10362
rect 27953 10310 27965 10362
rect 28017 10310 28029 10362
rect 28081 10310 28093 10362
rect 28145 10310 31832 10362
rect 1104 10288 31832 10310
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 20714 10248 20720 10260
rect 8168 10220 20720 10248
rect 8168 10208 8174 10220
rect 20714 10208 20720 10220
rect 20772 10208 20778 10260
rect 20990 10248 20996 10260
rect 20951 10220 20996 10248
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22646 10248 22652 10260
rect 22060 10220 22652 10248
rect 22060 10208 22066 10220
rect 22646 10208 22652 10220
rect 22704 10248 22710 10260
rect 22833 10251 22891 10257
rect 22833 10248 22845 10251
rect 22704 10220 22845 10248
rect 22704 10208 22710 10220
rect 22833 10217 22845 10220
rect 22879 10217 22891 10251
rect 23750 10248 23756 10260
rect 23711 10220 23756 10248
rect 22833 10211 22891 10217
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 24394 10208 24400 10260
rect 24452 10248 24458 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 24452 10220 24593 10248
rect 24452 10208 24458 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 25498 10248 25504 10260
rect 25459 10220 25504 10248
rect 24581 10211 24639 10217
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 28258 10208 28264 10260
rect 28316 10248 28322 10260
rect 29733 10251 29791 10257
rect 29733 10248 29745 10251
rect 28316 10220 29745 10248
rect 28316 10208 28322 10220
rect 29733 10217 29745 10220
rect 29779 10217 29791 10251
rect 30282 10248 30288 10260
rect 30243 10220 30288 10248
rect 29733 10211 29791 10217
rect 30282 10208 30288 10220
rect 30340 10208 30346 10260
rect 9306 10140 9312 10192
rect 9364 10180 9370 10192
rect 22186 10180 22192 10192
rect 9364 10152 22192 10180
rect 9364 10140 9370 10152
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 22281 10183 22339 10189
rect 22281 10149 22293 10183
rect 22327 10180 22339 10183
rect 25222 10180 25228 10192
rect 22327 10152 25228 10180
rect 22327 10149 22339 10152
rect 22281 10143 22339 10149
rect 25222 10140 25228 10152
rect 25280 10140 25286 10192
rect 20441 10115 20499 10121
rect 20441 10081 20453 10115
rect 20487 10112 20499 10115
rect 20898 10112 20904 10124
rect 20487 10084 20904 10112
rect 20487 10081 20499 10084
rect 20441 10075 20499 10081
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 21637 10115 21695 10121
rect 21637 10081 21649 10115
rect 21683 10112 21695 10115
rect 23106 10112 23112 10124
rect 21683 10084 23112 10112
rect 21683 10081 21695 10084
rect 21637 10075 21695 10081
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 26786 10112 26792 10124
rect 23256 10084 26792 10112
rect 23256 10072 23262 10084
rect 26786 10072 26792 10084
rect 26844 10072 26850 10124
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 21085 10047 21143 10053
rect 21085 10044 21097 10047
rect 13320 10016 21097 10044
rect 13320 10004 13326 10016
rect 21085 10013 21097 10016
rect 21131 10044 21143 10047
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 21131 10016 21557 10044
rect 21131 10013 21143 10016
rect 21085 10007 21143 10013
rect 21545 10013 21557 10016
rect 21591 10044 21603 10047
rect 22094 10044 22100 10056
rect 21591 10016 22100 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 22094 10004 22100 10016
rect 22152 10044 22158 10056
rect 22189 10047 22247 10053
rect 22189 10044 22201 10047
rect 22152 10016 22201 10044
rect 22152 10004 22158 10016
rect 22189 10013 22201 10016
rect 22235 10044 22247 10047
rect 23658 10044 23664 10056
rect 22235 10016 23664 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 23658 10004 23664 10016
rect 23716 10004 23722 10056
rect 26970 10004 26976 10056
rect 27028 10044 27034 10056
rect 27433 10047 27491 10053
rect 27433 10044 27445 10047
rect 27028 10016 27445 10044
rect 27028 10004 27034 10016
rect 27433 10013 27445 10016
rect 27479 10044 27491 10047
rect 31018 10044 31024 10056
rect 27479 10016 31024 10044
rect 27479 10013 27491 10016
rect 27433 10007 27491 10013
rect 31018 10004 31024 10016
rect 31076 10004 31082 10056
rect 31294 10044 31300 10056
rect 31255 10016 31300 10044
rect 31294 10004 31300 10016
rect 31352 10004 31358 10056
rect 4430 9936 4436 9988
rect 4488 9976 4494 9988
rect 4488 9948 26740 9976
rect 4488 9936 4494 9948
rect 26418 9868 26424 9920
rect 26476 9908 26482 9920
rect 26605 9911 26663 9917
rect 26605 9908 26617 9911
rect 26476 9880 26617 9908
rect 26476 9868 26482 9880
rect 26605 9877 26617 9880
rect 26651 9877 26663 9911
rect 26712 9908 26740 9948
rect 26878 9936 26884 9988
rect 26936 9976 26942 9988
rect 26936 9948 28856 9976
rect 26936 9936 26942 9948
rect 27893 9911 27951 9917
rect 27893 9908 27905 9911
rect 26712 9880 27905 9908
rect 26605 9871 26663 9877
rect 27893 9877 27905 9880
rect 27939 9908 27951 9911
rect 28442 9908 28448 9920
rect 27939 9880 28448 9908
rect 27939 9877 27951 9880
rect 27893 9871 27951 9877
rect 28442 9868 28448 9880
rect 28500 9868 28506 9920
rect 28828 9917 28856 9948
rect 28813 9911 28871 9917
rect 28813 9877 28825 9911
rect 28859 9908 28871 9911
rect 29178 9908 29184 9920
rect 28859 9880 29184 9908
rect 28859 9877 28871 9880
rect 28813 9871 28871 9877
rect 29178 9868 29184 9880
rect 29236 9868 29242 9920
rect 1104 9818 31992 9840
rect 1104 9766 8632 9818
rect 8684 9766 8696 9818
rect 8748 9766 8760 9818
rect 8812 9766 8824 9818
rect 8876 9766 8888 9818
rect 8940 9766 16314 9818
rect 16366 9766 16378 9818
rect 16430 9766 16442 9818
rect 16494 9766 16506 9818
rect 16558 9766 16570 9818
rect 16622 9766 23996 9818
rect 24048 9766 24060 9818
rect 24112 9766 24124 9818
rect 24176 9766 24188 9818
rect 24240 9766 24252 9818
rect 24304 9766 31678 9818
rect 31730 9766 31742 9818
rect 31794 9766 31806 9818
rect 31858 9766 31870 9818
rect 31922 9766 31934 9818
rect 31986 9766 31992 9818
rect 1104 9744 31992 9766
rect 21082 9704 21088 9716
rect 21043 9676 21088 9704
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 21910 9664 21916 9716
rect 21968 9704 21974 9716
rect 22094 9704 22100 9716
rect 21968 9676 22100 9704
rect 21968 9664 21974 9676
rect 22094 9664 22100 9676
rect 22152 9704 22158 9716
rect 22646 9704 22652 9716
rect 22152 9676 22245 9704
rect 22607 9676 22652 9704
rect 22152 9664 22158 9676
rect 22646 9664 22652 9676
rect 22704 9704 22710 9716
rect 23106 9704 23112 9716
rect 22704 9676 23112 9704
rect 22704 9664 22710 9676
rect 23106 9664 23112 9676
rect 23164 9704 23170 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23164 9676 23857 9704
rect 23164 9664 23170 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 24857 9707 24915 9713
rect 24857 9673 24869 9707
rect 24903 9704 24915 9707
rect 25498 9704 25504 9716
rect 24903 9676 25504 9704
rect 24903 9673 24915 9676
rect 24857 9667 24915 9673
rect 25498 9664 25504 9676
rect 25556 9664 25562 9716
rect 29638 9704 29644 9716
rect 29599 9676 29644 9704
rect 29638 9664 29644 9676
rect 29696 9664 29702 9716
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 20622 9636 20628 9648
rect 12400 9608 20628 9636
rect 12400 9596 12406 9608
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 25406 9636 25412 9648
rect 25367 9608 25412 9636
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 28445 9639 28503 9645
rect 28445 9605 28457 9639
rect 28491 9636 28503 9639
rect 28902 9636 28908 9648
rect 28491 9608 28908 9636
rect 28491 9605 28503 9608
rect 28445 9599 28503 9605
rect 28902 9596 28908 9608
rect 28960 9596 28966 9648
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 26602 9568 26608 9580
rect 6972 9540 26608 9568
rect 6972 9528 6978 9540
rect 26602 9528 26608 9540
rect 26660 9568 26666 9580
rect 28810 9568 28816 9580
rect 26660 9540 28816 9568
rect 26660 9528 26666 9540
rect 28810 9528 28816 9540
rect 28868 9528 28874 9580
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 24946 9500 24952 9512
rect 9180 9472 24952 9500
rect 9180 9460 9186 9472
rect 24946 9460 24952 9472
rect 25004 9460 25010 9512
rect 25222 9460 25228 9512
rect 25280 9500 25286 9512
rect 26050 9500 26056 9512
rect 25280 9472 26056 9500
rect 25280 9460 25286 9472
rect 26050 9460 26056 9472
rect 26108 9500 26114 9512
rect 27341 9503 27399 9509
rect 27341 9500 27353 9503
rect 26108 9472 27353 9500
rect 26108 9460 26114 9472
rect 27341 9469 27353 9472
rect 27387 9500 27399 9503
rect 30190 9500 30196 9512
rect 27387 9472 30196 9500
rect 27387 9469 27399 9472
rect 27341 9463 27399 9469
rect 30190 9460 30196 9472
rect 30248 9460 30254 9512
rect 10410 9392 10416 9444
rect 10468 9432 10474 9444
rect 23750 9432 23756 9444
rect 10468 9404 23756 9432
rect 10468 9392 10474 9404
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 25590 9432 25596 9444
rect 23860 9404 25596 9432
rect 7926 9324 7932 9376
rect 7984 9364 7990 9376
rect 23860 9364 23888 9404
rect 25590 9392 25596 9404
rect 25648 9432 25654 9444
rect 25869 9435 25927 9441
rect 25869 9432 25881 9435
rect 25648 9404 25881 9432
rect 25648 9392 25654 9404
rect 25869 9401 25881 9404
rect 25915 9401 25927 9435
rect 32858 9432 32864 9444
rect 25869 9395 25927 9401
rect 30116 9404 32864 9432
rect 30116 9376 30144 9404
rect 32858 9392 32864 9404
rect 32916 9392 32922 9444
rect 26418 9364 26424 9376
rect 7984 9336 23888 9364
rect 26379 9336 26424 9364
rect 7984 9324 7990 9336
rect 26418 9324 26424 9336
rect 26476 9364 26482 9376
rect 28997 9367 29055 9373
rect 28997 9364 29009 9367
rect 26476 9336 29009 9364
rect 26476 9324 26482 9336
rect 28997 9333 29009 9336
rect 29043 9333 29055 9367
rect 30098 9364 30104 9376
rect 30059 9336 30104 9364
rect 28997 9327 29055 9333
rect 30098 9324 30104 9336
rect 30156 9324 30162 9376
rect 31294 9364 31300 9376
rect 31255 9336 31300 9364
rect 31294 9324 31300 9336
rect 31352 9324 31358 9376
rect 1104 9274 31832 9296
rect 1104 9222 4791 9274
rect 4843 9222 4855 9274
rect 4907 9222 4919 9274
rect 4971 9222 4983 9274
rect 5035 9222 5047 9274
rect 5099 9222 12473 9274
rect 12525 9222 12537 9274
rect 12589 9222 12601 9274
rect 12653 9222 12665 9274
rect 12717 9222 12729 9274
rect 12781 9222 20155 9274
rect 20207 9222 20219 9274
rect 20271 9222 20283 9274
rect 20335 9222 20347 9274
rect 20399 9222 20411 9274
rect 20463 9222 27837 9274
rect 27889 9222 27901 9274
rect 27953 9222 27965 9274
rect 28017 9222 28029 9274
rect 28081 9222 28093 9274
rect 28145 9222 31832 9274
rect 1104 9200 31832 9222
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 22922 9160 22928 9172
rect 6880 9132 22928 9160
rect 6880 9120 6886 9132
rect 22922 9120 22928 9132
rect 22980 9120 22986 9172
rect 23106 9160 23112 9172
rect 23067 9132 23112 9160
rect 23106 9120 23112 9132
rect 23164 9120 23170 9172
rect 30190 9160 30196 9172
rect 30151 9132 30196 9160
rect 30190 9120 30196 9132
rect 30248 9120 30254 9172
rect 24857 9095 24915 9101
rect 24857 9061 24869 9095
rect 24903 9092 24915 9095
rect 25314 9092 25320 9104
rect 24903 9064 25320 9092
rect 24903 9061 24915 9064
rect 24857 9055 24915 9061
rect 25314 9052 25320 9064
rect 25372 9092 25378 9104
rect 26053 9095 26111 9101
rect 26053 9092 26065 9095
rect 25372 9064 26065 9092
rect 25372 9052 25378 9064
rect 26053 9061 26065 9064
rect 26099 9092 26111 9095
rect 26142 9092 26148 9104
rect 26099 9064 26148 9092
rect 26099 9061 26111 9064
rect 26053 9055 26111 9061
rect 26142 9052 26148 9064
rect 26200 9052 26206 9104
rect 27430 9052 27436 9104
rect 27488 9092 27494 9104
rect 28077 9095 28135 9101
rect 28077 9092 28089 9095
rect 27488 9064 28089 9092
rect 27488 9052 27494 9064
rect 28077 9061 28089 9064
rect 28123 9092 28135 9095
rect 28166 9092 28172 9104
rect 28123 9064 28172 9092
rect 28123 9061 28135 9064
rect 28077 9055 28135 9061
rect 28166 9052 28172 9064
rect 28224 9052 28230 9104
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 23753 9027 23811 9033
rect 23753 9024 23765 9027
rect 9640 8996 23765 9024
rect 9640 8984 9646 8996
rect 23753 8993 23765 8996
rect 23799 9024 23811 9027
rect 23842 9024 23848 9036
rect 23799 8996 23848 9024
rect 23799 8993 23811 8996
rect 23753 8987 23811 8993
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 27706 9024 27712 9036
rect 24780 8996 27712 9024
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5500 8928 6914 8956
rect 5500 8916 5506 8928
rect 6886 8888 6914 8928
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 24780 8956 24808 8996
rect 27706 8984 27712 8996
rect 27764 8984 27770 9036
rect 28534 9024 28540 9036
rect 28495 8996 28540 9024
rect 28534 8984 28540 8996
rect 28592 9024 28598 9036
rect 30837 9027 30895 9033
rect 30837 9024 30849 9027
rect 28592 8996 30849 9024
rect 28592 8984 28598 8996
rect 30837 8993 30849 8996
rect 30883 8993 30895 9027
rect 30837 8987 30895 8993
rect 20680 8928 24808 8956
rect 26697 8959 26755 8965
rect 20680 8916 20686 8928
rect 26697 8925 26709 8959
rect 26743 8956 26755 8959
rect 28350 8956 28356 8968
rect 26743 8928 28356 8956
rect 26743 8925 26755 8928
rect 26697 8919 26755 8925
rect 28350 8916 28356 8928
rect 28408 8956 28414 8968
rect 29638 8956 29644 8968
rect 28408 8928 29644 8956
rect 28408 8916 28414 8928
rect 29638 8916 29644 8928
rect 29696 8916 29702 8968
rect 27433 8891 27491 8897
rect 27433 8888 27445 8891
rect 6886 8860 27445 8888
rect 27433 8857 27445 8860
rect 27479 8857 27491 8891
rect 27433 8851 27491 8857
rect 21910 8820 21916 8832
rect 21823 8792 21916 8820
rect 21910 8780 21916 8792
rect 21968 8820 21974 8832
rect 22554 8820 22560 8832
rect 21968 8792 22560 8820
rect 21968 8780 21974 8792
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 25222 8780 25228 8832
rect 25280 8820 25286 8832
rect 25317 8823 25375 8829
rect 25317 8820 25329 8823
rect 25280 8792 25329 8820
rect 25280 8780 25286 8792
rect 25317 8789 25329 8792
rect 25363 8789 25375 8823
rect 29086 8820 29092 8832
rect 29047 8792 29092 8820
rect 25317 8783 25375 8789
rect 29086 8780 29092 8792
rect 29144 8780 29150 8832
rect 1104 8730 31992 8752
rect 1104 8678 8632 8730
rect 8684 8678 8696 8730
rect 8748 8678 8760 8730
rect 8812 8678 8824 8730
rect 8876 8678 8888 8730
rect 8940 8678 16314 8730
rect 16366 8678 16378 8730
rect 16430 8678 16442 8730
rect 16494 8678 16506 8730
rect 16558 8678 16570 8730
rect 16622 8678 23996 8730
rect 24048 8678 24060 8730
rect 24112 8678 24124 8730
rect 24176 8678 24188 8730
rect 24240 8678 24252 8730
rect 24304 8678 31678 8730
rect 31730 8678 31742 8730
rect 31794 8678 31806 8730
rect 31858 8678 31870 8730
rect 31922 8678 31934 8730
rect 31986 8678 31992 8730
rect 1104 8656 31992 8678
rect 23106 8576 23112 8628
rect 23164 8616 23170 8628
rect 23661 8619 23719 8625
rect 23661 8616 23673 8619
rect 23164 8588 23673 8616
rect 23164 8576 23170 8588
rect 23661 8585 23673 8588
rect 23707 8616 23719 8619
rect 24305 8619 24363 8625
rect 24305 8616 24317 8619
rect 23707 8588 24317 8616
rect 23707 8585 23719 8588
rect 23661 8579 23719 8585
rect 24305 8585 24317 8588
rect 24351 8616 24363 8619
rect 24857 8619 24915 8625
rect 24857 8616 24869 8619
rect 24351 8588 24869 8616
rect 24351 8585 24363 8588
rect 24305 8579 24363 8585
rect 24857 8585 24869 8588
rect 24903 8585 24915 8619
rect 25498 8616 25504 8628
rect 25459 8588 25504 8616
rect 24857 8579 24915 8585
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 26234 8576 26240 8628
rect 26292 8616 26298 8628
rect 26513 8619 26571 8625
rect 26513 8616 26525 8619
rect 26292 8588 26525 8616
rect 26292 8576 26298 8588
rect 26513 8585 26525 8588
rect 26559 8585 26571 8619
rect 26513 8579 26571 8585
rect 27062 8576 27068 8628
rect 27120 8616 27126 8628
rect 27157 8619 27215 8625
rect 27157 8616 27169 8619
rect 27120 8588 27169 8616
rect 27120 8576 27126 8588
rect 27157 8585 27169 8588
rect 27203 8585 27215 8619
rect 29178 8616 29184 8628
rect 29139 8588 29184 8616
rect 27157 8579 27215 8585
rect 29178 8576 29184 8588
rect 29236 8576 29242 8628
rect 29730 8616 29736 8628
rect 29691 8588 29736 8616
rect 29730 8576 29736 8588
rect 29788 8576 29794 8628
rect 28629 8551 28687 8557
rect 28629 8517 28641 8551
rect 28675 8548 28687 8551
rect 32030 8548 32036 8560
rect 28675 8520 32036 8548
rect 28675 8517 28687 8520
rect 28629 8511 28687 8517
rect 32030 8508 32036 8520
rect 32088 8508 32094 8560
rect 22922 8440 22928 8492
rect 22980 8480 22986 8492
rect 30742 8480 30748 8492
rect 22980 8452 30748 8480
rect 22980 8440 22986 8452
rect 30742 8440 30748 8452
rect 30800 8440 30806 8492
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14332 8384 22508 8412
rect 14332 8372 14338 8384
rect 1578 8344 1584 8356
rect 1539 8316 1584 8344
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 21358 8276 21364 8288
rect 9548 8248 21364 8276
rect 9548 8236 9554 8248
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 22480 8276 22508 8384
rect 22554 8372 22560 8424
rect 22612 8412 22618 8424
rect 23201 8415 23259 8421
rect 23201 8412 23213 8415
rect 22612 8384 23213 8412
rect 22612 8372 22618 8384
rect 23201 8381 23213 8384
rect 23247 8412 23259 8415
rect 28442 8412 28448 8424
rect 23247 8384 28448 8412
rect 23247 8381 23259 8384
rect 23201 8375 23259 8381
rect 28442 8372 28448 8384
rect 28500 8372 28506 8424
rect 26234 8344 26240 8356
rect 26206 8304 26240 8344
rect 26292 8344 26298 8356
rect 27709 8347 27767 8353
rect 27709 8344 27721 8347
rect 26292 8316 27721 8344
rect 26292 8304 26298 8316
rect 27709 8313 27721 8316
rect 27755 8344 27767 8347
rect 28810 8344 28816 8356
rect 27755 8316 28816 8344
rect 27755 8313 27767 8316
rect 27709 8307 27767 8313
rect 28810 8304 28816 8316
rect 28868 8304 28874 8356
rect 30374 8344 30380 8356
rect 30335 8316 30380 8344
rect 30374 8304 30380 8316
rect 30432 8304 30438 8356
rect 31294 8344 31300 8356
rect 31255 8316 31300 8344
rect 31294 8304 31300 8316
rect 31352 8304 31358 8356
rect 26050 8276 26056 8288
rect 22480 8248 26056 8276
rect 26050 8236 26056 8248
rect 26108 8276 26114 8288
rect 26206 8276 26234 8304
rect 26108 8248 26234 8276
rect 26108 8236 26114 8248
rect 1104 8186 31832 8208
rect 1104 8134 4791 8186
rect 4843 8134 4855 8186
rect 4907 8134 4919 8186
rect 4971 8134 4983 8186
rect 5035 8134 5047 8186
rect 5099 8134 12473 8186
rect 12525 8134 12537 8186
rect 12589 8134 12601 8186
rect 12653 8134 12665 8186
rect 12717 8134 12729 8186
rect 12781 8134 20155 8186
rect 20207 8134 20219 8186
rect 20271 8134 20283 8186
rect 20335 8134 20347 8186
rect 20399 8134 20411 8186
rect 20463 8134 27837 8186
rect 27889 8134 27901 8186
rect 27953 8134 27965 8186
rect 28017 8134 28029 8186
rect 28081 8134 28093 8186
rect 28145 8134 31832 8186
rect 1104 8112 31832 8134
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 10376 8044 22094 8072
rect 10376 8032 10382 8044
rect 22066 8004 22094 8044
rect 25222 8032 25228 8084
rect 25280 8072 25286 8084
rect 25866 8072 25872 8084
rect 25280 8044 25872 8072
rect 25280 8032 25286 8044
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 26513 8075 26571 8081
rect 26513 8041 26525 8075
rect 26559 8072 26571 8075
rect 26786 8072 26792 8084
rect 26559 8044 26792 8072
rect 26559 8041 26571 8044
rect 26513 8035 26571 8041
rect 26786 8032 26792 8044
rect 26844 8032 26850 8084
rect 27249 8075 27307 8081
rect 27249 8041 27261 8075
rect 27295 8072 27307 8075
rect 27430 8072 27436 8084
rect 27295 8044 27436 8072
rect 27295 8041 27307 8044
rect 27249 8035 27307 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 28350 8072 28356 8084
rect 28311 8044 28356 8072
rect 28350 8032 28356 8044
rect 28408 8032 28414 8084
rect 28810 8072 28816 8084
rect 28771 8044 28816 8072
rect 28810 8032 28816 8044
rect 28868 8072 28874 8084
rect 29730 8072 29736 8084
rect 28868 8044 29736 8072
rect 28868 8032 28874 8044
rect 29730 8032 29736 8044
rect 29788 8032 29794 8084
rect 30469 8075 30527 8081
rect 30469 8041 30481 8075
rect 30515 8072 30527 8075
rect 30742 8072 30748 8084
rect 30515 8044 30748 8072
rect 30515 8041 30527 8044
rect 30469 8035 30527 8041
rect 30742 8032 30748 8044
rect 30800 8032 30806 8084
rect 31021 8075 31079 8081
rect 31021 8041 31033 8075
rect 31067 8072 31079 8075
rect 31386 8072 31392 8084
rect 31067 8044 31392 8072
rect 31067 8041 31079 8044
rect 31021 8035 31079 8041
rect 31386 8032 31392 8044
rect 31444 8032 31450 8084
rect 32306 8004 32312 8016
rect 22066 7976 32312 8004
rect 32306 7964 32312 7976
rect 32364 7964 32370 8016
rect 21358 7896 21364 7948
rect 21416 7936 21422 7948
rect 21416 7908 27384 7936
rect 21416 7896 21422 7908
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 27246 7868 27252 7880
rect 7708 7840 27252 7868
rect 7708 7828 7714 7840
rect 27246 7828 27252 7840
rect 27304 7828 27310 7880
rect 27356 7868 27384 7908
rect 27614 7896 27620 7948
rect 27672 7936 27678 7948
rect 27801 7939 27859 7945
rect 27801 7936 27813 7939
rect 27672 7908 27813 7936
rect 27672 7896 27678 7908
rect 27801 7905 27813 7908
rect 27847 7936 27859 7939
rect 29178 7936 29184 7948
rect 27847 7908 29184 7936
rect 27847 7905 27859 7908
rect 27801 7899 27859 7905
rect 29178 7896 29184 7908
rect 29236 7936 29242 7948
rect 30190 7936 30196 7948
rect 29236 7908 30196 7936
rect 29236 7896 29242 7908
rect 30190 7896 30196 7908
rect 30248 7896 30254 7948
rect 32766 7868 32772 7880
rect 27356 7840 32772 7868
rect 32766 7828 32772 7840
rect 32824 7828 32830 7880
rect 22066 7772 25452 7800
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 22066 7732 22094 7772
rect 24854 7732 24860 7744
rect 9272 7704 22094 7732
rect 24815 7704 24860 7732
rect 9272 7692 9278 7704
rect 24854 7692 24860 7704
rect 24912 7692 24918 7744
rect 25424 7741 25452 7772
rect 28350 7760 28356 7812
rect 28408 7800 28414 7812
rect 29086 7800 29092 7812
rect 28408 7772 29092 7800
rect 28408 7760 28414 7772
rect 29086 7760 29092 7772
rect 29144 7760 29150 7812
rect 25409 7735 25467 7741
rect 25409 7701 25421 7735
rect 25455 7732 25467 7735
rect 26326 7732 26332 7744
rect 25455 7704 26332 7732
rect 25455 7701 25467 7704
rect 25409 7695 25467 7701
rect 26326 7692 26332 7704
rect 26384 7732 26390 7744
rect 26694 7732 26700 7744
rect 26384 7704 26700 7732
rect 26384 7692 26390 7704
rect 26694 7692 26700 7704
rect 26752 7692 26758 7744
rect 1104 7642 31992 7664
rect 1104 7590 8632 7642
rect 8684 7590 8696 7642
rect 8748 7590 8760 7642
rect 8812 7590 8824 7642
rect 8876 7590 8888 7642
rect 8940 7590 16314 7642
rect 16366 7590 16378 7642
rect 16430 7590 16442 7642
rect 16494 7590 16506 7642
rect 16558 7590 16570 7642
rect 16622 7590 23996 7642
rect 24048 7590 24060 7642
rect 24112 7590 24124 7642
rect 24176 7590 24188 7642
rect 24240 7590 24252 7642
rect 24304 7590 31678 7642
rect 31730 7590 31742 7642
rect 31794 7590 31806 7642
rect 31858 7590 31870 7642
rect 31922 7590 31934 7642
rect 31986 7590 31992 7642
rect 1104 7568 31992 7590
rect 25682 7488 25688 7540
rect 25740 7528 25746 7540
rect 28261 7531 28319 7537
rect 28261 7528 28273 7531
rect 25740 7500 28273 7528
rect 25740 7488 25746 7500
rect 28261 7497 28273 7500
rect 28307 7497 28319 7531
rect 28261 7491 28319 7497
rect 28905 7531 28963 7537
rect 28905 7497 28917 7531
rect 28951 7528 28963 7531
rect 32122 7528 32128 7540
rect 28951 7500 32128 7528
rect 28951 7497 28963 7500
rect 28905 7491 28963 7497
rect 32122 7488 32128 7500
rect 32180 7488 32186 7540
rect 26050 7460 26056 7472
rect 26011 7432 26056 7460
rect 26050 7420 26056 7432
rect 26108 7420 26114 7472
rect 26602 7460 26608 7472
rect 26563 7432 26608 7460
rect 26602 7420 26608 7432
rect 26660 7420 26666 7472
rect 27522 7420 27528 7472
rect 27580 7460 27586 7472
rect 27617 7463 27675 7469
rect 27617 7460 27629 7463
rect 27580 7432 27629 7460
rect 27580 7420 27586 7432
rect 27617 7429 27629 7432
rect 27663 7429 27675 7463
rect 27617 7423 27675 7429
rect 28534 7420 28540 7472
rect 28592 7460 28598 7472
rect 29365 7463 29423 7469
rect 29365 7460 29377 7463
rect 28592 7432 29377 7460
rect 28592 7420 28598 7432
rect 29365 7429 29377 7432
rect 29411 7429 29423 7463
rect 30466 7460 30472 7472
rect 30427 7432 30472 7460
rect 29365 7423 29423 7429
rect 30466 7420 30472 7432
rect 30524 7420 30530 7472
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 26786 7392 26792 7404
rect 24912 7364 26792 7392
rect 24912 7352 24918 7364
rect 26786 7352 26792 7364
rect 26844 7352 26850 7404
rect 29914 7324 29920 7336
rect 29875 7296 29920 7324
rect 29914 7284 29920 7296
rect 29972 7324 29978 7336
rect 30282 7324 30288 7336
rect 29972 7296 30288 7324
rect 29972 7284 29978 7296
rect 30282 7284 30288 7296
rect 30340 7284 30346 7336
rect 31294 7256 31300 7268
rect 31255 7228 31300 7256
rect 31294 7216 31300 7228
rect 31352 7216 31358 7268
rect 24946 7188 24952 7200
rect 24859 7160 24952 7188
rect 24946 7148 24952 7160
rect 25004 7188 25010 7200
rect 25501 7191 25559 7197
rect 25501 7188 25513 7191
rect 25004 7160 25513 7188
rect 25004 7148 25010 7160
rect 25501 7157 25513 7160
rect 25547 7188 25559 7191
rect 25682 7188 25688 7200
rect 25547 7160 25688 7188
rect 25547 7157 25559 7160
rect 25501 7151 25559 7157
rect 25682 7148 25688 7160
rect 25740 7148 25746 7200
rect 1104 7098 31832 7120
rect 1104 7046 4791 7098
rect 4843 7046 4855 7098
rect 4907 7046 4919 7098
rect 4971 7046 4983 7098
rect 5035 7046 5047 7098
rect 5099 7046 12473 7098
rect 12525 7046 12537 7098
rect 12589 7046 12601 7098
rect 12653 7046 12665 7098
rect 12717 7046 12729 7098
rect 12781 7046 20155 7098
rect 20207 7046 20219 7098
rect 20271 7046 20283 7098
rect 20335 7046 20347 7098
rect 20399 7046 20411 7098
rect 20463 7046 27837 7098
rect 27889 7046 27901 7098
rect 27953 7046 27965 7098
rect 28017 7046 28029 7098
rect 28081 7046 28093 7098
rect 28145 7046 31832 7098
rect 1104 7024 31832 7046
rect 25866 6876 25872 6928
rect 25924 6916 25930 6928
rect 25924 6888 27384 6916
rect 25924 6876 25930 6888
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 27356 6848 27384 6888
rect 28169 6851 28227 6857
rect 28169 6848 28181 6851
rect 4304 6820 6914 6848
rect 27356 6820 28181 6848
rect 4304 6808 4310 6820
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 6886 6780 6914 6820
rect 28169 6817 28181 6820
rect 28215 6817 28227 6851
rect 28169 6811 28227 6817
rect 29089 6851 29147 6857
rect 29089 6817 29101 6851
rect 29135 6848 29147 6851
rect 29454 6848 29460 6860
rect 29135 6820 29460 6848
rect 29135 6817 29147 6820
rect 29089 6811 29147 6817
rect 29454 6808 29460 6820
rect 29512 6808 29518 6860
rect 30009 6851 30067 6857
rect 30009 6817 30021 6851
rect 30055 6848 30067 6851
rect 31110 6848 31116 6860
rect 30055 6820 31116 6848
rect 30055 6817 30067 6820
rect 30009 6811 30067 6817
rect 31110 6808 31116 6820
rect 31168 6808 31174 6860
rect 26418 6780 26424 6792
rect 6886 6752 26424 6780
rect 26418 6740 26424 6752
rect 26476 6780 26482 6792
rect 29362 6780 29368 6792
rect 26476 6752 29368 6780
rect 26476 6740 26482 6752
rect 29362 6740 29368 6752
rect 29420 6740 29426 6792
rect 31018 6780 31024 6792
rect 30979 6752 31024 6780
rect 31018 6740 31024 6752
rect 31076 6740 31082 6792
rect 27341 6715 27399 6721
rect 27341 6681 27353 6715
rect 27387 6712 27399 6715
rect 27614 6712 27620 6724
rect 27387 6684 27620 6712
rect 27387 6681 27399 6684
rect 27341 6675 27399 6681
rect 27614 6672 27620 6684
rect 27672 6672 27678 6724
rect 30466 6712 30472 6724
rect 30427 6684 30472 6712
rect 30466 6672 30472 6684
rect 30524 6672 30530 6724
rect 25682 6644 25688 6656
rect 25643 6616 25688 6644
rect 25682 6604 25688 6616
rect 25740 6604 25746 6656
rect 26234 6644 26240 6656
rect 26195 6616 26240 6644
rect 26234 6604 26240 6616
rect 26292 6604 26298 6656
rect 26786 6644 26792 6656
rect 26747 6616 26792 6644
rect 26786 6604 26792 6616
rect 26844 6604 26850 6656
rect 1104 6554 31992 6576
rect 1104 6502 8632 6554
rect 8684 6502 8696 6554
rect 8748 6502 8760 6554
rect 8812 6502 8824 6554
rect 8876 6502 8888 6554
rect 8940 6502 16314 6554
rect 16366 6502 16378 6554
rect 16430 6502 16442 6554
rect 16494 6502 16506 6554
rect 16558 6502 16570 6554
rect 16622 6502 23996 6554
rect 24048 6502 24060 6554
rect 24112 6502 24124 6554
rect 24176 6502 24188 6554
rect 24240 6502 24252 6554
rect 24304 6502 31678 6554
rect 31730 6502 31742 6554
rect 31794 6502 31806 6554
rect 31858 6502 31870 6554
rect 31922 6502 31934 6554
rect 31986 6502 31992 6554
rect 1104 6480 31992 6502
rect 29730 6440 29736 6452
rect 29691 6412 29736 6440
rect 29730 6400 29736 6412
rect 29788 6400 29794 6452
rect 25682 6196 25688 6248
rect 25740 6236 25746 6248
rect 26605 6239 26663 6245
rect 26605 6236 26617 6239
rect 25740 6208 26617 6236
rect 25740 6196 25746 6208
rect 26605 6205 26617 6208
rect 26651 6236 26663 6239
rect 27614 6236 27620 6248
rect 26651 6208 27620 6236
rect 26651 6205 26663 6208
rect 26605 6199 26663 6205
rect 27614 6196 27620 6208
rect 27672 6196 27678 6248
rect 28718 6236 28724 6248
rect 28679 6208 28724 6236
rect 28718 6196 28724 6208
rect 28776 6236 28782 6248
rect 30377 6239 30435 6245
rect 30377 6236 30389 6239
rect 28776 6208 30389 6236
rect 28776 6196 28782 6208
rect 30377 6205 30389 6208
rect 30423 6205 30435 6239
rect 30377 6199 30435 6205
rect 28169 6171 28227 6177
rect 28169 6168 28181 6171
rect 22066 6140 28181 6168
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 22066 6100 22094 6140
rect 28169 6137 28181 6140
rect 28215 6168 28227 6171
rect 29086 6168 29092 6180
rect 28215 6140 29092 6168
rect 28215 6137 28227 6140
rect 28169 6131 28227 6137
rect 29086 6128 29092 6140
rect 29144 6128 29150 6180
rect 27706 6100 27712 6112
rect 4580 6072 22094 6100
rect 27667 6072 27712 6100
rect 4580 6060 4586 6072
rect 27706 6060 27712 6072
rect 27764 6060 27770 6112
rect 31294 6100 31300 6112
rect 31255 6072 31300 6100
rect 31294 6060 31300 6072
rect 31352 6060 31358 6112
rect 1104 6010 31832 6032
rect 1104 5958 4791 6010
rect 4843 5958 4855 6010
rect 4907 5958 4919 6010
rect 4971 5958 4983 6010
rect 5035 5958 5047 6010
rect 5099 5958 12473 6010
rect 12525 5958 12537 6010
rect 12589 5958 12601 6010
rect 12653 5958 12665 6010
rect 12717 5958 12729 6010
rect 12781 5958 20155 6010
rect 20207 5958 20219 6010
rect 20271 5958 20283 6010
rect 20335 5958 20347 6010
rect 20399 5958 20411 6010
rect 20463 5958 27837 6010
rect 27889 5958 27901 6010
rect 27953 5958 27965 6010
rect 28017 5958 28029 6010
rect 28081 5958 28093 6010
rect 28145 5958 31832 6010
rect 1104 5936 31832 5958
rect 28629 5899 28687 5905
rect 28629 5896 28641 5899
rect 22066 5868 28641 5896
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 22066 5692 22094 5868
rect 28629 5865 28641 5868
rect 28675 5896 28687 5899
rect 28994 5896 29000 5908
rect 28675 5868 29000 5896
rect 28675 5865 28687 5868
rect 28629 5859 28687 5865
rect 28994 5856 29000 5868
rect 29052 5856 29058 5908
rect 29178 5896 29184 5908
rect 29139 5868 29184 5896
rect 29178 5856 29184 5868
rect 29236 5856 29242 5908
rect 27706 5788 27712 5840
rect 27764 5828 27770 5840
rect 28258 5828 28264 5840
rect 27764 5800 28264 5828
rect 27764 5788 27770 5800
rect 28258 5788 28264 5800
rect 28316 5828 28322 5840
rect 29733 5831 29791 5837
rect 29733 5828 29745 5831
rect 28316 5800 29745 5828
rect 28316 5788 28322 5800
rect 29733 5797 29745 5800
rect 29779 5797 29791 5831
rect 29733 5791 29791 5797
rect 26602 5720 26608 5772
rect 26660 5760 26666 5772
rect 30285 5763 30343 5769
rect 30285 5760 30297 5763
rect 26660 5732 30297 5760
rect 26660 5720 26666 5732
rect 30285 5729 30297 5732
rect 30331 5729 30343 5763
rect 30285 5723 30343 5729
rect 31294 5692 31300 5704
rect 8536 5664 22094 5692
rect 31255 5664 31300 5692
rect 8536 5652 8542 5664
rect 31294 5652 31300 5664
rect 31352 5652 31358 5704
rect 27525 5559 27583 5565
rect 27525 5525 27537 5559
rect 27571 5556 27583 5559
rect 27614 5556 27620 5568
rect 27571 5528 27620 5556
rect 27571 5525 27583 5528
rect 27525 5519 27583 5525
rect 27614 5516 27620 5528
rect 27672 5556 27678 5568
rect 28077 5559 28135 5565
rect 28077 5556 28089 5559
rect 27672 5528 28089 5556
rect 27672 5516 27678 5528
rect 28077 5525 28089 5528
rect 28123 5556 28135 5559
rect 28350 5556 28356 5568
rect 28123 5528 28356 5556
rect 28123 5525 28135 5528
rect 28077 5519 28135 5525
rect 28350 5516 28356 5528
rect 28408 5516 28414 5568
rect 1104 5466 31992 5488
rect 1104 5414 8632 5466
rect 8684 5414 8696 5466
rect 8748 5414 8760 5466
rect 8812 5414 8824 5466
rect 8876 5414 8888 5466
rect 8940 5414 16314 5466
rect 16366 5414 16378 5466
rect 16430 5414 16442 5466
rect 16494 5414 16506 5466
rect 16558 5414 16570 5466
rect 16622 5414 23996 5466
rect 24048 5414 24060 5466
rect 24112 5414 24124 5466
rect 24176 5414 24188 5466
rect 24240 5414 24252 5466
rect 24304 5414 31678 5466
rect 31730 5414 31742 5466
rect 31794 5414 31806 5466
rect 31858 5414 31870 5466
rect 31922 5414 31934 5466
rect 31986 5414 31992 5466
rect 1104 5392 31992 5414
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 27801 5355 27859 5361
rect 8260 5324 27292 5352
rect 8260 5312 8266 5324
rect 12158 5244 12164 5296
rect 12216 5284 12222 5296
rect 27154 5284 27160 5296
rect 12216 5256 27160 5284
rect 12216 5244 12222 5256
rect 27154 5244 27160 5256
rect 27212 5244 27218 5296
rect 27264 5284 27292 5324
rect 27801 5321 27813 5355
rect 27847 5352 27859 5355
rect 31202 5352 31208 5364
rect 27847 5324 31208 5352
rect 27847 5321 27859 5324
rect 27801 5315 27859 5321
rect 31202 5312 31208 5324
rect 31260 5312 31266 5364
rect 30650 5284 30656 5296
rect 27264 5256 30656 5284
rect 30650 5244 30656 5256
rect 30708 5244 30714 5296
rect 24394 5176 24400 5228
rect 24452 5216 24458 5228
rect 30929 5219 30987 5225
rect 30929 5216 30941 5219
rect 24452 5188 30941 5216
rect 24452 5176 24458 5188
rect 30929 5185 30941 5188
rect 30975 5185 30987 5219
rect 30929 5179 30987 5185
rect 26234 5108 26240 5160
rect 26292 5148 26298 5160
rect 29362 5148 29368 5160
rect 26292 5120 29040 5148
rect 29323 5120 29368 5148
rect 26292 5108 26298 5120
rect 29012 5080 29040 5120
rect 29362 5108 29368 5120
rect 29420 5108 29426 5160
rect 30377 5083 30435 5089
rect 30377 5080 30389 5083
rect 29012 5052 30389 5080
rect 30377 5049 30389 5052
rect 30423 5049 30435 5083
rect 30377 5043 30435 5049
rect 28350 5012 28356 5024
rect 28311 4984 28356 5012
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 28442 4972 28448 5024
rect 28500 5012 28506 5024
rect 28902 5012 28908 5024
rect 28500 4984 28908 5012
rect 28500 4972 28506 4984
rect 28902 4972 28908 4984
rect 28960 4972 28966 5024
rect 1104 4922 31832 4944
rect 1104 4870 4791 4922
rect 4843 4870 4855 4922
rect 4907 4870 4919 4922
rect 4971 4870 4983 4922
rect 5035 4870 5047 4922
rect 5099 4870 12473 4922
rect 12525 4870 12537 4922
rect 12589 4870 12601 4922
rect 12653 4870 12665 4922
rect 12717 4870 12729 4922
rect 12781 4870 20155 4922
rect 20207 4870 20219 4922
rect 20271 4870 20283 4922
rect 20335 4870 20347 4922
rect 20399 4870 20411 4922
rect 20463 4870 27837 4922
rect 27889 4870 27901 4922
rect 27953 4870 27965 4922
rect 28017 4870 28029 4922
rect 28081 4870 28093 4922
rect 28145 4870 31832 4922
rect 1104 4848 31832 4870
rect 28902 4768 28908 4820
rect 28960 4808 28966 4820
rect 29089 4811 29147 4817
rect 29089 4808 29101 4811
rect 28960 4780 29101 4808
rect 28960 4768 28966 4780
rect 29089 4777 29101 4780
rect 29135 4777 29147 4811
rect 29089 4771 29147 4777
rect 26142 4700 26148 4752
rect 26200 4740 26206 4752
rect 29917 4743 29975 4749
rect 29917 4740 29929 4743
rect 26200 4712 29929 4740
rect 26200 4700 26206 4712
rect 29917 4709 29929 4712
rect 29963 4709 29975 4743
rect 29917 4703 29975 4709
rect 27246 4632 27252 4684
rect 27304 4672 27310 4684
rect 30469 4675 30527 4681
rect 30469 4672 30481 4675
rect 27304 4644 30481 4672
rect 27304 4632 27310 4644
rect 30469 4641 30481 4644
rect 30515 4641 30527 4675
rect 30469 4635 30527 4641
rect 26786 4564 26792 4616
rect 26844 4604 26850 4616
rect 31021 4607 31079 4613
rect 31021 4604 31033 4607
rect 26844 4576 31033 4604
rect 26844 4564 26850 4576
rect 31021 4573 31033 4576
rect 31067 4573 31079 4607
rect 31021 4567 31079 4573
rect 1104 4378 31992 4400
rect 1104 4326 8632 4378
rect 8684 4326 8696 4378
rect 8748 4326 8760 4378
rect 8812 4326 8824 4378
rect 8876 4326 8888 4378
rect 8940 4326 16314 4378
rect 16366 4326 16378 4378
rect 16430 4326 16442 4378
rect 16494 4326 16506 4378
rect 16558 4326 16570 4378
rect 16622 4326 23996 4378
rect 24048 4326 24060 4378
rect 24112 4326 24124 4378
rect 24176 4326 24188 4378
rect 24240 4326 24252 4378
rect 24304 4326 31678 4378
rect 31730 4326 31742 4378
rect 31794 4326 31806 4378
rect 31858 4326 31870 4378
rect 31922 4326 31934 4378
rect 31986 4326 31992 4378
rect 1104 4304 31992 4326
rect 29917 4131 29975 4137
rect 29917 4097 29929 4131
rect 29963 4128 29975 4131
rect 30558 4128 30564 4140
rect 29963 4100 30564 4128
rect 29963 4097 29975 4100
rect 29917 4091 29975 4097
rect 30558 4088 30564 4100
rect 30616 4088 30622 4140
rect 1578 4060 1584 4072
rect 1539 4032 1584 4060
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 28350 3884 28356 3936
rect 28408 3924 28414 3936
rect 30466 3924 30472 3936
rect 28408 3896 30472 3924
rect 28408 3884 28414 3896
rect 30466 3884 30472 3896
rect 30524 3884 30530 3936
rect 31294 3924 31300 3936
rect 31255 3896 31300 3924
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 1104 3834 31832 3856
rect 1104 3782 4791 3834
rect 4843 3782 4855 3834
rect 4907 3782 4919 3834
rect 4971 3782 4983 3834
rect 5035 3782 5047 3834
rect 5099 3782 12473 3834
rect 12525 3782 12537 3834
rect 12589 3782 12601 3834
rect 12653 3782 12665 3834
rect 12717 3782 12729 3834
rect 12781 3782 20155 3834
rect 20207 3782 20219 3834
rect 20271 3782 20283 3834
rect 20335 3782 20347 3834
rect 20399 3782 20411 3834
rect 20463 3782 27837 3834
rect 27889 3782 27901 3834
rect 27953 3782 27965 3834
rect 28017 3782 28029 3834
rect 28081 3782 28093 3834
rect 28145 3782 31832 3834
rect 1104 3760 31832 3782
rect 30466 3680 30472 3732
rect 30524 3720 30530 3732
rect 30561 3723 30619 3729
rect 30561 3720 30573 3723
rect 30524 3692 30573 3720
rect 30524 3680 30530 3692
rect 30561 3689 30573 3692
rect 30607 3689 30619 3723
rect 30561 3683 30619 3689
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 31294 3516 31300 3528
rect 31255 3488 31300 3516
rect 31294 3476 31300 3488
rect 31352 3476 31358 3528
rect 1104 3290 31992 3312
rect 1104 3238 8632 3290
rect 8684 3238 8696 3290
rect 8748 3238 8760 3290
rect 8812 3238 8824 3290
rect 8876 3238 8888 3290
rect 8940 3238 16314 3290
rect 16366 3238 16378 3290
rect 16430 3238 16442 3290
rect 16494 3238 16506 3290
rect 16558 3238 16570 3290
rect 16622 3238 23996 3290
rect 24048 3238 24060 3290
rect 24112 3238 24124 3290
rect 24176 3238 24188 3290
rect 24240 3238 24252 3290
rect 24304 3238 31678 3290
rect 31730 3238 31742 3290
rect 31794 3238 31806 3290
rect 31858 3238 31870 3290
rect 31922 3238 31934 3290
rect 31986 3238 31992 3290
rect 1104 3216 31992 3238
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 1104 2746 31832 2768
rect 1104 2694 4791 2746
rect 4843 2694 4855 2746
rect 4907 2694 4919 2746
rect 4971 2694 4983 2746
rect 5035 2694 5047 2746
rect 5099 2694 12473 2746
rect 12525 2694 12537 2746
rect 12589 2694 12601 2746
rect 12653 2694 12665 2746
rect 12717 2694 12729 2746
rect 12781 2694 20155 2746
rect 20207 2694 20219 2746
rect 20271 2694 20283 2746
rect 20335 2694 20347 2746
rect 20399 2694 20411 2746
rect 20463 2694 27837 2746
rect 27889 2694 27901 2746
rect 27953 2694 27965 2746
rect 28017 2694 28029 2746
rect 28081 2694 28093 2746
rect 28145 2694 31832 2746
rect 1104 2672 31832 2694
rect 1394 2388 1400 2440
rect 1452 2428 1458 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1452 2400 1593 2428
rect 1452 2388 1458 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1104 2202 31992 2224
rect 1104 2150 8632 2202
rect 8684 2150 8696 2202
rect 8748 2150 8760 2202
rect 8812 2150 8824 2202
rect 8876 2150 8888 2202
rect 8940 2150 16314 2202
rect 16366 2150 16378 2202
rect 16430 2150 16442 2202
rect 16494 2150 16506 2202
rect 16558 2150 16570 2202
rect 16622 2150 23996 2202
rect 24048 2150 24060 2202
rect 24112 2150 24124 2202
rect 24176 2150 24188 2202
rect 24240 2150 24252 2202
rect 24304 2150 31678 2202
rect 31730 2150 31742 2202
rect 31794 2150 31806 2202
rect 31858 2150 31870 2202
rect 31922 2150 31934 2202
rect 31986 2150 31992 2202
rect 1104 2128 31992 2150
<< via1 >>
rect 9128 33464 9180 33516
rect 27528 33464 27580 33516
rect 10140 33328 10192 33380
rect 24584 33328 24636 33380
rect 12900 33260 12952 33312
rect 27620 33260 27672 33312
rect 13176 33192 13228 33244
rect 25412 33192 25464 33244
rect 12808 33124 12860 33176
rect 25688 33124 25740 33176
rect 10508 32920 10560 32972
rect 22100 32920 22152 32972
rect 13636 32784 13688 32836
rect 18236 32784 18288 32836
rect 19892 32784 19944 32836
rect 25228 32784 25280 32836
rect 9588 32716 9640 32768
rect 21640 32716 21692 32768
rect 8632 32614 8684 32666
rect 8696 32614 8748 32666
rect 8760 32614 8812 32666
rect 8824 32614 8876 32666
rect 8888 32614 8940 32666
rect 16314 32614 16366 32666
rect 16378 32614 16430 32666
rect 16442 32614 16494 32666
rect 16506 32614 16558 32666
rect 16570 32614 16622 32666
rect 23996 32614 24048 32666
rect 24060 32614 24112 32666
rect 24124 32614 24176 32666
rect 24188 32614 24240 32666
rect 24252 32614 24304 32666
rect 31678 32614 31730 32666
rect 31742 32614 31794 32666
rect 31806 32614 31858 32666
rect 31870 32614 31922 32666
rect 31934 32614 31986 32666
rect 18236 32555 18288 32564
rect 18236 32521 18245 32555
rect 18245 32521 18279 32555
rect 18279 32521 18288 32555
rect 18236 32512 18288 32521
rect 21272 32512 21324 32564
rect 24584 32555 24636 32564
rect 24584 32521 24593 32555
rect 24593 32521 24627 32555
rect 24627 32521 24636 32555
rect 24584 32512 24636 32521
rect 21456 32487 21508 32496
rect 21456 32453 21465 32487
rect 21465 32453 21499 32487
rect 21499 32453 21508 32487
rect 21456 32444 21508 32453
rect 24860 32444 24912 32496
rect 25136 32444 25188 32496
rect 28172 32444 28224 32496
rect 940 32376 992 32428
rect 2228 32419 2280 32428
rect 2228 32385 2237 32419
rect 2237 32385 2271 32419
rect 2271 32385 2280 32419
rect 2228 32376 2280 32385
rect 2872 32419 2924 32428
rect 2872 32385 2881 32419
rect 2881 32385 2915 32419
rect 2915 32385 2924 32419
rect 2872 32376 2924 32385
rect 4620 32419 4672 32428
rect 4620 32385 4629 32419
rect 4629 32385 4663 32419
rect 4663 32385 4672 32419
rect 4620 32376 4672 32385
rect 5816 32419 5868 32428
rect 5816 32385 5825 32419
rect 5825 32385 5859 32419
rect 5859 32385 5868 32419
rect 5816 32376 5868 32385
rect 8208 32419 8260 32428
rect 8208 32385 8217 32419
rect 8217 32385 8251 32419
rect 8251 32385 8260 32419
rect 8208 32376 8260 32385
rect 9404 32419 9456 32428
rect 9404 32385 9413 32419
rect 9413 32385 9447 32419
rect 9447 32385 9456 32419
rect 9404 32376 9456 32385
rect 11796 32419 11848 32428
rect 11796 32385 11805 32419
rect 11805 32385 11839 32419
rect 11839 32385 11848 32419
rect 11796 32376 11848 32385
rect 12992 32419 13044 32428
rect 12992 32385 13001 32419
rect 13001 32385 13035 32419
rect 13035 32385 13044 32419
rect 12992 32376 13044 32385
rect 15384 32419 15436 32428
rect 15384 32385 15393 32419
rect 15393 32385 15427 32419
rect 15427 32385 15436 32419
rect 15384 32376 15436 32385
rect 16672 32376 16724 32428
rect 18880 32376 18932 32428
rect 20076 32376 20128 32428
rect 22468 32376 22520 32428
rect 23664 32376 23716 32428
rect 23848 32376 23900 32428
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 26056 32376 26108 32428
rect 27252 32376 27304 32428
rect 29644 32376 29696 32428
rect 30932 32419 30984 32428
rect 30932 32385 30941 32419
rect 30941 32385 30975 32419
rect 30975 32385 30984 32419
rect 30932 32376 30984 32385
rect 13544 32308 13596 32360
rect 20628 32308 20680 32360
rect 21180 32308 21232 32360
rect 26516 32308 26568 32360
rect 27528 32308 27580 32360
rect 32220 32308 32272 32360
rect 11612 32240 11664 32292
rect 14832 32240 14884 32292
rect 14924 32283 14976 32292
rect 14924 32249 14933 32283
rect 14933 32249 14967 32283
rect 14967 32249 14976 32283
rect 14924 32240 14976 32249
rect 16948 32240 17000 32292
rect 19064 32240 19116 32292
rect 21548 32240 21600 32292
rect 23112 32240 23164 32292
rect 26884 32240 26936 32292
rect 28356 32283 28408 32292
rect 28356 32249 28365 32283
rect 28365 32249 28399 32283
rect 28399 32249 28408 32283
rect 28356 32240 28408 32249
rect 12348 32172 12400 32224
rect 13084 32172 13136 32224
rect 15108 32172 15160 32224
rect 16028 32172 16080 32224
rect 17776 32215 17828 32224
rect 17776 32181 17785 32215
rect 17785 32181 17819 32215
rect 17819 32181 17828 32215
rect 17776 32172 17828 32181
rect 18788 32172 18840 32224
rect 21088 32172 21140 32224
rect 22376 32172 22428 32224
rect 23296 32215 23348 32224
rect 23296 32181 23305 32215
rect 23305 32181 23339 32215
rect 23339 32181 23348 32215
rect 23296 32172 23348 32181
rect 23572 32172 23624 32224
rect 25044 32172 25096 32224
rect 25228 32172 25280 32224
rect 30288 32172 30340 32224
rect 30840 32172 30892 32224
rect 4791 32070 4843 32122
rect 4855 32070 4907 32122
rect 4919 32070 4971 32122
rect 4983 32070 5035 32122
rect 5047 32070 5099 32122
rect 12473 32070 12525 32122
rect 12537 32070 12589 32122
rect 12601 32070 12653 32122
rect 12665 32070 12717 32122
rect 12729 32070 12781 32122
rect 20155 32070 20207 32122
rect 20219 32070 20271 32122
rect 20283 32070 20335 32122
rect 20347 32070 20399 32122
rect 20411 32070 20463 32122
rect 27837 32070 27889 32122
rect 27901 32070 27953 32122
rect 27965 32070 28017 32122
rect 28029 32070 28081 32122
rect 28093 32070 28145 32122
rect 1584 32011 1636 32020
rect 1584 31977 1593 32011
rect 1593 31977 1627 32011
rect 1627 31977 1636 32011
rect 1584 31968 1636 31977
rect 14832 31968 14884 32020
rect 18236 31968 18288 32020
rect 18788 32011 18840 32020
rect 18788 31977 18797 32011
rect 18797 31977 18831 32011
rect 18831 31977 18840 32011
rect 18788 31968 18840 31977
rect 19892 32011 19944 32020
rect 19892 31977 19901 32011
rect 19901 31977 19935 32011
rect 19935 31977 19944 32011
rect 19892 31968 19944 31977
rect 19984 31968 20036 32020
rect 21180 32011 21232 32020
rect 11888 31900 11940 31952
rect 20076 31900 20128 31952
rect 21180 31977 21189 32011
rect 21189 31977 21223 32011
rect 21223 31977 21232 32011
rect 21180 31968 21232 31977
rect 22744 31968 22796 32020
rect 23112 32011 23164 32020
rect 23112 31977 23121 32011
rect 23121 31977 23155 32011
rect 23155 31977 23164 32011
rect 23112 31968 23164 31977
rect 23848 32011 23900 32020
rect 23848 31977 23857 32011
rect 23857 31977 23891 32011
rect 23891 31977 23900 32011
rect 23848 31968 23900 31977
rect 24492 31968 24544 32020
rect 25228 32011 25280 32020
rect 25228 31977 25237 32011
rect 25237 31977 25271 32011
rect 25271 31977 25280 32011
rect 25228 31968 25280 31977
rect 24584 31900 24636 31952
rect 24768 31900 24820 31952
rect 26332 31968 26384 32020
rect 26516 32011 26568 32020
rect 26516 31977 26525 32011
rect 26525 31977 26559 32011
rect 26559 31977 26568 32011
rect 26516 31968 26568 31977
rect 27528 31968 27580 32020
rect 30564 32011 30616 32020
rect 30564 31977 30573 32011
rect 30573 31977 30607 32011
rect 30607 31977 30616 32011
rect 30564 31968 30616 31977
rect 29276 31900 29328 31952
rect 31208 31943 31260 31952
rect 31208 31909 31217 31943
rect 31217 31909 31251 31943
rect 31251 31909 31260 31943
rect 31208 31900 31260 31909
rect 15936 31832 15988 31884
rect 24400 31832 24452 31884
rect 14740 31764 14792 31816
rect 15844 31764 15896 31816
rect 16672 31807 16724 31816
rect 16672 31773 16681 31807
rect 16681 31773 16715 31807
rect 16715 31773 16724 31807
rect 16672 31764 16724 31773
rect 20812 31764 20864 31816
rect 21180 31764 21232 31816
rect 10324 31696 10376 31748
rect 14464 31739 14516 31748
rect 14464 31705 14473 31739
rect 14473 31705 14507 31739
rect 14507 31705 14516 31739
rect 14464 31696 14516 31705
rect 15660 31696 15712 31748
rect 18328 31696 18380 31748
rect 24676 31764 24728 31816
rect 24768 31807 24820 31816
rect 24768 31773 24777 31807
rect 24777 31773 24811 31807
rect 24811 31773 24820 31807
rect 27712 31832 27764 31884
rect 32496 31832 32548 31884
rect 24768 31764 24820 31773
rect 11520 31671 11572 31680
rect 11520 31637 11529 31671
rect 11529 31637 11563 31671
rect 11563 31637 11572 31671
rect 11520 31628 11572 31637
rect 12348 31628 12400 31680
rect 14648 31628 14700 31680
rect 16212 31628 16264 31680
rect 17408 31628 17460 31680
rect 19892 31628 19944 31680
rect 21824 31628 21876 31680
rect 23112 31628 23164 31680
rect 23848 31628 23900 31680
rect 25780 31764 25832 31816
rect 26148 31764 26200 31816
rect 29736 31807 29788 31816
rect 29736 31773 29745 31807
rect 29745 31773 29779 31807
rect 29779 31773 29788 31807
rect 29736 31764 29788 31773
rect 29828 31764 29880 31816
rect 26976 31696 27028 31748
rect 27712 31696 27764 31748
rect 28724 31739 28776 31748
rect 28724 31705 28733 31739
rect 28733 31705 28767 31739
rect 28767 31705 28776 31739
rect 28724 31696 28776 31705
rect 28816 31628 28868 31680
rect 8632 31526 8684 31578
rect 8696 31526 8748 31578
rect 8760 31526 8812 31578
rect 8824 31526 8876 31578
rect 8888 31526 8940 31578
rect 16314 31526 16366 31578
rect 16378 31526 16430 31578
rect 16442 31526 16494 31578
rect 16506 31526 16558 31578
rect 16570 31526 16622 31578
rect 23996 31526 24048 31578
rect 24060 31526 24112 31578
rect 24124 31526 24176 31578
rect 24188 31526 24240 31578
rect 24252 31526 24304 31578
rect 31678 31526 31730 31578
rect 31742 31526 31794 31578
rect 31806 31526 31858 31578
rect 31870 31526 31922 31578
rect 31934 31526 31986 31578
rect 16764 31424 16816 31476
rect 16948 31424 17000 31476
rect 19156 31424 19208 31476
rect 21456 31424 21508 31476
rect 22744 31424 22796 31476
rect 23756 31424 23808 31476
rect 23848 31424 23900 31476
rect 24492 31424 24544 31476
rect 24584 31424 24636 31476
rect 28264 31467 28316 31476
rect 28264 31433 28273 31467
rect 28273 31433 28307 31467
rect 28307 31433 28316 31467
rect 28264 31424 28316 31433
rect 14740 31356 14792 31408
rect 17040 31356 17092 31408
rect 21180 31399 21232 31408
rect 21180 31365 21189 31399
rect 21189 31365 21223 31399
rect 21223 31365 21232 31399
rect 21180 31356 21232 31365
rect 22100 31399 22152 31408
rect 22100 31365 22109 31399
rect 22109 31365 22143 31399
rect 22143 31365 22152 31399
rect 22100 31356 22152 31365
rect 13544 31331 13596 31340
rect 13544 31297 13553 31331
rect 13553 31297 13587 31331
rect 13587 31297 13596 31331
rect 13544 31288 13596 31297
rect 14832 31288 14884 31340
rect 18420 31288 18472 31340
rect 20536 31288 20588 31340
rect 22100 31220 22152 31272
rect 22192 31220 22244 31272
rect 23572 31288 23624 31340
rect 23756 31288 23808 31340
rect 24492 31288 24544 31340
rect 23664 31220 23716 31272
rect 23848 31220 23900 31272
rect 12348 31152 12400 31204
rect 16212 31152 16264 31204
rect 18052 31152 18104 31204
rect 18144 31152 18196 31204
rect 22376 31152 22428 31204
rect 22468 31152 22520 31204
rect 25872 31288 25924 31340
rect 26148 31288 26200 31340
rect 27160 31288 27212 31340
rect 30748 31288 30800 31340
rect 26700 31220 26752 31272
rect 25044 31152 25096 31204
rect 26608 31152 26660 31204
rect 1584 31127 1636 31136
rect 1584 31093 1593 31127
rect 1593 31093 1627 31127
rect 1627 31093 1636 31127
rect 1584 31084 1636 31093
rect 10508 31127 10560 31136
rect 10508 31093 10517 31127
rect 10517 31093 10551 31127
rect 10551 31093 10560 31127
rect 10508 31084 10560 31093
rect 11796 31084 11848 31136
rect 12164 31084 12216 31136
rect 12808 31084 12860 31136
rect 14004 31127 14056 31136
rect 14004 31093 14013 31127
rect 14013 31093 14047 31127
rect 14047 31093 14056 31127
rect 14004 31084 14056 31093
rect 14740 31084 14792 31136
rect 15568 31084 15620 31136
rect 17224 31084 17276 31136
rect 17776 31084 17828 31136
rect 18972 31084 19024 31136
rect 19800 31084 19852 31136
rect 22008 31084 22060 31136
rect 23756 31084 23808 31136
rect 23848 31084 23900 31136
rect 24308 31127 24360 31136
rect 24308 31093 24317 31127
rect 24317 31093 24351 31127
rect 24351 31093 24360 31127
rect 24308 31084 24360 31093
rect 24584 31084 24636 31136
rect 24768 31084 24820 31136
rect 24860 31084 24912 31136
rect 25504 31084 25556 31136
rect 32128 31220 32180 31272
rect 26884 31152 26936 31204
rect 27252 31127 27304 31136
rect 27252 31093 27261 31127
rect 27261 31093 27295 31127
rect 27295 31093 27304 31127
rect 27252 31084 27304 31093
rect 27344 31084 27396 31136
rect 29368 31084 29420 31136
rect 30012 31127 30064 31136
rect 30012 31093 30021 31127
rect 30021 31093 30055 31127
rect 30055 31093 30064 31127
rect 30012 31084 30064 31093
rect 30656 31127 30708 31136
rect 30656 31093 30665 31127
rect 30665 31093 30699 31127
rect 30699 31093 30708 31127
rect 30656 31084 30708 31093
rect 32036 31084 32088 31136
rect 4791 30982 4843 31034
rect 4855 30982 4907 31034
rect 4919 30982 4971 31034
rect 4983 30982 5035 31034
rect 5047 30982 5099 31034
rect 12473 30982 12525 31034
rect 12537 30982 12589 31034
rect 12601 30982 12653 31034
rect 12665 30982 12717 31034
rect 12729 30982 12781 31034
rect 20155 30982 20207 31034
rect 20219 30982 20271 31034
rect 20283 30982 20335 31034
rect 20347 30982 20399 31034
rect 20411 30982 20463 31034
rect 27837 30982 27889 31034
rect 27901 30982 27953 31034
rect 27965 30982 28017 31034
rect 28029 30982 28081 31034
rect 28093 30982 28145 31034
rect 9036 30880 9088 30932
rect 10324 30923 10376 30932
rect 10324 30889 10333 30923
rect 10333 30889 10367 30923
rect 10367 30889 10376 30923
rect 10324 30880 10376 30889
rect 4068 30812 4120 30864
rect 14004 30880 14056 30932
rect 16120 30923 16172 30932
rect 16120 30889 16129 30923
rect 16129 30889 16163 30923
rect 16163 30889 16172 30923
rect 16120 30880 16172 30889
rect 17224 30880 17276 30932
rect 17684 30923 17736 30932
rect 17684 30889 17693 30923
rect 17693 30889 17727 30923
rect 17727 30889 17736 30923
rect 17684 30880 17736 30889
rect 18328 30923 18380 30932
rect 18328 30889 18337 30923
rect 18337 30889 18371 30923
rect 18371 30889 18380 30923
rect 18328 30880 18380 30889
rect 18696 30880 18748 30932
rect 19340 30880 19392 30932
rect 23020 30880 23072 30932
rect 24584 30880 24636 30932
rect 24768 30923 24820 30932
rect 24768 30889 24777 30923
rect 24777 30889 24811 30923
rect 24811 30889 24820 30923
rect 24768 30880 24820 30889
rect 24952 30923 25004 30932
rect 24952 30889 24961 30923
rect 24961 30889 24995 30923
rect 24995 30889 25004 30923
rect 24952 30880 25004 30889
rect 25228 30880 25280 30932
rect 11888 30812 11940 30864
rect 21364 30812 21416 30864
rect 21456 30812 21508 30864
rect 11428 30787 11480 30796
rect 11428 30753 11437 30787
rect 11437 30753 11471 30787
rect 11471 30753 11480 30787
rect 11428 30744 11480 30753
rect 11796 30744 11848 30796
rect 13084 30744 13136 30796
rect 11060 30676 11112 30728
rect 11520 30676 11572 30728
rect 12072 30676 12124 30728
rect 12256 30676 12308 30728
rect 15568 30676 15620 30728
rect 13360 30608 13412 30660
rect 17132 30651 17184 30660
rect 17132 30617 17141 30651
rect 17141 30617 17175 30651
rect 17175 30617 17184 30651
rect 17132 30608 17184 30617
rect 17500 30744 17552 30796
rect 17868 30676 17920 30728
rect 22376 30676 22428 30728
rect 22836 30676 22888 30728
rect 23204 30812 23256 30864
rect 26240 30812 26292 30864
rect 28724 30880 28776 30932
rect 28816 30923 28868 30932
rect 28816 30889 28825 30923
rect 28825 30889 28859 30923
rect 28859 30889 28868 30923
rect 28816 30880 28868 30889
rect 29736 30812 29788 30864
rect 23388 30744 23440 30796
rect 23296 30719 23348 30728
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 23572 30676 23624 30728
rect 18052 30608 18104 30660
rect 11244 30540 11296 30592
rect 12348 30540 12400 30592
rect 14648 30540 14700 30592
rect 15660 30540 15712 30592
rect 15752 30540 15804 30592
rect 17684 30540 17736 30592
rect 18972 30540 19024 30592
rect 19524 30583 19576 30592
rect 19524 30549 19533 30583
rect 19533 30549 19567 30583
rect 19567 30549 19576 30583
rect 19524 30540 19576 30549
rect 20352 30583 20404 30592
rect 20352 30549 20361 30583
rect 20361 30549 20395 30583
rect 20395 30549 20404 30583
rect 20352 30540 20404 30549
rect 20904 30583 20956 30592
rect 20904 30549 20913 30583
rect 20913 30549 20947 30583
rect 20947 30549 20956 30583
rect 20904 30540 20956 30549
rect 21732 30608 21784 30660
rect 22928 30608 22980 30660
rect 24492 30608 24544 30660
rect 24676 30608 24728 30660
rect 28448 30744 28500 30796
rect 23020 30540 23072 30592
rect 23848 30540 23900 30592
rect 25228 30540 25280 30592
rect 25504 30540 25556 30592
rect 26608 30676 26660 30728
rect 26424 30608 26476 30660
rect 25964 30540 26016 30592
rect 27436 30676 27488 30728
rect 28172 30676 28224 30728
rect 28356 30719 28408 30728
rect 28356 30685 28365 30719
rect 28365 30685 28399 30719
rect 28399 30685 28408 30719
rect 28356 30676 28408 30685
rect 30472 30676 30524 30728
rect 31576 30676 31628 30728
rect 28908 30608 28960 30660
rect 29000 30540 29052 30592
rect 30104 30583 30156 30592
rect 30104 30549 30113 30583
rect 30113 30549 30147 30583
rect 30147 30549 30156 30583
rect 30104 30540 30156 30549
rect 30564 30583 30616 30592
rect 30564 30549 30573 30583
rect 30573 30549 30607 30583
rect 30607 30549 30616 30583
rect 30564 30540 30616 30549
rect 8632 30438 8684 30490
rect 8696 30438 8748 30490
rect 8760 30438 8812 30490
rect 8824 30438 8876 30490
rect 8888 30438 8940 30490
rect 16314 30438 16366 30490
rect 16378 30438 16430 30490
rect 16442 30438 16494 30490
rect 16506 30438 16558 30490
rect 16570 30438 16622 30490
rect 23996 30438 24048 30490
rect 24060 30438 24112 30490
rect 24124 30438 24176 30490
rect 24188 30438 24240 30490
rect 24252 30438 24304 30490
rect 31678 30438 31730 30490
rect 31742 30438 31794 30490
rect 31806 30438 31858 30490
rect 31870 30438 31922 30490
rect 31934 30438 31986 30490
rect 2688 30336 2740 30388
rect 9036 30268 9088 30320
rect 10048 30336 10100 30388
rect 11152 30336 11204 30388
rect 14648 30336 14700 30388
rect 14924 30336 14976 30388
rect 19248 30336 19300 30388
rect 19432 30336 19484 30388
rect 9864 30200 9916 30252
rect 12348 30268 12400 30320
rect 13636 30268 13688 30320
rect 16120 30268 16172 30320
rect 19340 30268 19392 30320
rect 19800 30268 19852 30320
rect 20444 30311 20496 30320
rect 20444 30277 20453 30311
rect 20453 30277 20487 30311
rect 20487 30277 20496 30311
rect 20444 30268 20496 30277
rect 20628 30268 20680 30320
rect 21364 30336 21416 30388
rect 23112 30336 23164 30388
rect 12072 30200 12124 30252
rect 18328 30200 18380 30252
rect 18604 30200 18656 30252
rect 22376 30200 22428 30252
rect 22652 30268 22704 30320
rect 23204 30311 23256 30320
rect 23204 30277 23213 30311
rect 23213 30277 23247 30311
rect 23247 30277 23256 30311
rect 23204 30268 23256 30277
rect 22928 30243 22980 30252
rect 22928 30209 22937 30243
rect 22937 30209 22971 30243
rect 22971 30209 22980 30243
rect 22928 30200 22980 30209
rect 23756 30224 23808 30276
rect 24216 30268 24268 30320
rect 24952 30336 25004 30388
rect 25044 30336 25096 30388
rect 25320 30336 25372 30388
rect 25504 30336 25556 30388
rect 25872 30336 25924 30388
rect 26240 30336 26292 30388
rect 26884 30336 26936 30388
rect 1584 30175 1636 30184
rect 1584 30141 1593 30175
rect 1593 30141 1627 30175
rect 1627 30141 1636 30175
rect 1584 30132 1636 30141
rect 14096 30132 14148 30184
rect 14188 30132 14240 30184
rect 15108 30175 15160 30184
rect 15108 30141 15117 30175
rect 15117 30141 15151 30175
rect 15151 30141 15160 30175
rect 15108 30132 15160 30141
rect 15476 30132 15528 30184
rect 17408 30132 17460 30184
rect 20076 30132 20128 30184
rect 21180 30132 21232 30184
rect 23020 30132 23072 30184
rect 23112 30132 23164 30184
rect 23756 30132 23808 30184
rect 24676 30200 24728 30252
rect 24952 30200 25004 30252
rect 25504 30243 25556 30252
rect 25504 30209 25513 30243
rect 25513 30209 25547 30243
rect 25547 30209 25556 30243
rect 25504 30200 25556 30209
rect 25228 30132 25280 30184
rect 25412 30132 25464 30184
rect 9496 30039 9548 30048
rect 9496 30005 9505 30039
rect 9505 30005 9539 30039
rect 9539 30005 9548 30039
rect 9496 29996 9548 30005
rect 10416 29996 10468 30048
rect 18144 30064 18196 30116
rect 12808 29996 12860 30048
rect 12992 30039 13044 30048
rect 12992 30005 13001 30039
rect 13001 30005 13035 30039
rect 13035 30005 13044 30039
rect 12992 29996 13044 30005
rect 13268 29996 13320 30048
rect 14372 29996 14424 30048
rect 14464 29996 14516 30048
rect 16028 29996 16080 30048
rect 17408 29996 17460 30048
rect 17960 29996 18012 30048
rect 18604 29996 18656 30048
rect 18880 30039 18932 30048
rect 18880 30005 18889 30039
rect 18889 30005 18923 30039
rect 18923 30005 18932 30039
rect 18880 29996 18932 30005
rect 19248 30064 19300 30116
rect 21548 30064 21600 30116
rect 21916 30064 21968 30116
rect 22928 30064 22980 30116
rect 23572 30064 23624 30116
rect 22192 29996 22244 30048
rect 22652 29996 22704 30048
rect 23112 30039 23164 30048
rect 23112 30005 23121 30039
rect 23121 30005 23155 30039
rect 23155 30005 23164 30039
rect 23112 29996 23164 30005
rect 23204 29996 23256 30048
rect 24124 30064 24176 30116
rect 24768 30064 24820 30116
rect 26792 30268 26844 30320
rect 27988 30336 28040 30388
rect 27068 30200 27120 30252
rect 26056 30132 26108 30184
rect 30012 30268 30064 30320
rect 30104 30268 30156 30320
rect 26240 30064 26292 30116
rect 26792 30064 26844 30116
rect 27988 30243 28040 30252
rect 27988 30209 27997 30243
rect 27997 30209 28031 30243
rect 28031 30209 28040 30243
rect 27988 30200 28040 30209
rect 28540 30200 28592 30252
rect 28908 30200 28960 30252
rect 29736 30243 29788 30252
rect 29736 30209 29745 30243
rect 29745 30209 29779 30243
rect 29779 30209 29788 30243
rect 29736 30200 29788 30209
rect 30196 30200 30248 30252
rect 27436 30132 27488 30184
rect 27896 30132 27948 30184
rect 29552 30132 29604 30184
rect 24676 30039 24728 30048
rect 24676 30005 24685 30039
rect 24685 30005 24719 30039
rect 24719 30005 24728 30039
rect 24676 29996 24728 30005
rect 27068 29996 27120 30048
rect 27344 29996 27396 30048
rect 28080 29996 28132 30048
rect 28632 30039 28684 30048
rect 28632 30005 28641 30039
rect 28641 30005 28675 30039
rect 28675 30005 28684 30039
rect 28632 29996 28684 30005
rect 29828 30064 29880 30116
rect 29460 29996 29512 30048
rect 30380 29996 30432 30048
rect 30564 30039 30616 30048
rect 30564 30005 30573 30039
rect 30573 30005 30607 30039
rect 30607 30005 30616 30039
rect 30564 29996 30616 30005
rect 31208 30039 31260 30048
rect 31208 30005 31217 30039
rect 31217 30005 31251 30039
rect 31251 30005 31260 30039
rect 31208 29996 31260 30005
rect 4791 29894 4843 29946
rect 4855 29894 4907 29946
rect 4919 29894 4971 29946
rect 4983 29894 5035 29946
rect 5047 29894 5099 29946
rect 12473 29894 12525 29946
rect 12537 29894 12589 29946
rect 12601 29894 12653 29946
rect 12665 29894 12717 29946
rect 12729 29894 12781 29946
rect 20155 29894 20207 29946
rect 20219 29894 20271 29946
rect 20283 29894 20335 29946
rect 20347 29894 20399 29946
rect 20411 29894 20463 29946
rect 27837 29894 27889 29946
rect 27901 29894 27953 29946
rect 27965 29894 28017 29946
rect 28029 29894 28081 29946
rect 28093 29894 28145 29946
rect 11244 29792 11296 29844
rect 13360 29792 13412 29844
rect 14372 29792 14424 29844
rect 16856 29792 16908 29844
rect 16948 29792 17000 29844
rect 17776 29792 17828 29844
rect 18236 29792 18288 29844
rect 19432 29792 19484 29844
rect 19984 29792 20036 29844
rect 20352 29792 20404 29844
rect 20720 29792 20772 29844
rect 21364 29792 21416 29844
rect 22100 29792 22152 29844
rect 24124 29792 24176 29844
rect 24216 29792 24268 29844
rect 24860 29792 24912 29844
rect 25228 29792 25280 29844
rect 25872 29835 25924 29844
rect 25872 29801 25881 29835
rect 25881 29801 25915 29835
rect 25915 29801 25924 29835
rect 25872 29792 25924 29801
rect 26148 29792 26200 29844
rect 26332 29792 26384 29844
rect 26608 29835 26660 29844
rect 26608 29801 26617 29835
rect 26617 29801 26651 29835
rect 26651 29801 26660 29835
rect 26608 29792 26660 29801
rect 26976 29792 27028 29844
rect 29184 29792 29236 29844
rect 9956 29724 10008 29776
rect 10508 29724 10560 29776
rect 14188 29724 14240 29776
rect 9404 29588 9456 29640
rect 9588 29520 9640 29572
rect 11152 29656 11204 29708
rect 11244 29656 11296 29708
rect 13084 29656 13136 29708
rect 16212 29724 16264 29776
rect 18788 29724 18840 29776
rect 20260 29724 20312 29776
rect 14648 29656 14700 29708
rect 19248 29656 19300 29708
rect 19616 29656 19668 29708
rect 19892 29656 19944 29708
rect 20628 29656 20680 29708
rect 21180 29724 21232 29776
rect 17132 29588 17184 29640
rect 19524 29588 19576 29640
rect 19984 29588 20036 29640
rect 20720 29588 20772 29640
rect 21272 29656 21324 29708
rect 21916 29724 21968 29776
rect 22836 29724 22888 29776
rect 23940 29724 23992 29776
rect 26056 29724 26108 29776
rect 28356 29724 28408 29776
rect 30104 29724 30156 29776
rect 12348 29520 12400 29572
rect 14832 29520 14884 29572
rect 7840 29452 7892 29504
rect 10508 29452 10560 29504
rect 12072 29495 12124 29504
rect 12072 29461 12081 29495
rect 12081 29461 12115 29495
rect 12115 29461 12124 29495
rect 12072 29452 12124 29461
rect 14188 29452 14240 29504
rect 15016 29452 15068 29504
rect 17040 29520 17092 29572
rect 17684 29520 17736 29572
rect 16028 29452 16080 29504
rect 16856 29452 16908 29504
rect 17224 29452 17276 29504
rect 17592 29495 17644 29504
rect 17592 29461 17601 29495
rect 17601 29461 17635 29495
rect 17635 29461 17644 29495
rect 17592 29452 17644 29461
rect 18328 29452 18380 29504
rect 19064 29520 19116 29572
rect 20168 29520 20220 29572
rect 20352 29520 20404 29572
rect 20444 29520 20496 29572
rect 21180 29588 21232 29640
rect 21456 29631 21508 29640
rect 21456 29597 21465 29631
rect 21465 29597 21499 29631
rect 21499 29597 21508 29631
rect 21456 29588 21508 29597
rect 21916 29588 21968 29640
rect 22284 29656 22336 29708
rect 22560 29588 22612 29640
rect 23572 29656 23624 29708
rect 23756 29656 23808 29708
rect 26332 29656 26384 29708
rect 27436 29656 27488 29708
rect 27528 29656 27580 29708
rect 27712 29656 27764 29708
rect 20996 29520 21048 29572
rect 22192 29520 22244 29572
rect 23296 29588 23348 29640
rect 23664 29631 23716 29640
rect 23664 29597 23673 29631
rect 23673 29597 23707 29631
rect 23707 29597 23716 29631
rect 23664 29588 23716 29597
rect 24676 29588 24728 29640
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 25596 29588 25648 29640
rect 26516 29631 26568 29640
rect 22836 29452 22888 29504
rect 23572 29520 23624 29572
rect 24216 29452 24268 29504
rect 25872 29495 25924 29504
rect 25872 29461 25899 29495
rect 25899 29461 25924 29495
rect 25872 29452 25924 29461
rect 26240 29520 26292 29572
rect 26516 29597 26525 29631
rect 26525 29597 26559 29631
rect 26559 29597 26568 29631
rect 26516 29588 26568 29597
rect 27896 29588 27948 29640
rect 28080 29631 28132 29640
rect 28080 29597 28089 29631
rect 28089 29597 28123 29631
rect 28123 29597 28132 29631
rect 28080 29588 28132 29597
rect 27344 29452 27396 29504
rect 28632 29656 28684 29708
rect 28816 29631 28868 29640
rect 28816 29597 28825 29631
rect 28825 29597 28859 29631
rect 28859 29597 28868 29631
rect 28816 29588 28868 29597
rect 28356 29520 28408 29572
rect 28632 29520 28684 29572
rect 29000 29588 29052 29640
rect 29920 29631 29972 29640
rect 29920 29597 29929 29631
rect 29929 29597 29963 29631
rect 29963 29597 29972 29631
rect 29920 29588 29972 29597
rect 31116 29588 31168 29640
rect 29000 29452 29052 29504
rect 31024 29452 31076 29504
rect 31300 29452 31352 29504
rect 8632 29350 8684 29402
rect 8696 29350 8748 29402
rect 8760 29350 8812 29402
rect 8824 29350 8876 29402
rect 8888 29350 8940 29402
rect 16314 29350 16366 29402
rect 16378 29350 16430 29402
rect 16442 29350 16494 29402
rect 16506 29350 16558 29402
rect 16570 29350 16622 29402
rect 23996 29350 24048 29402
rect 24060 29350 24112 29402
rect 24124 29350 24176 29402
rect 24188 29350 24240 29402
rect 24252 29350 24304 29402
rect 31678 29350 31730 29402
rect 31742 29350 31794 29402
rect 31806 29350 31858 29402
rect 31870 29350 31922 29402
rect 31934 29350 31986 29402
rect 10416 29248 10468 29300
rect 9036 29180 9088 29232
rect 12256 29248 12308 29300
rect 12808 29248 12860 29300
rect 13636 29248 13688 29300
rect 12072 29180 12124 29232
rect 11152 29112 11204 29164
rect 11888 29112 11940 29164
rect 13728 29180 13780 29232
rect 15476 29248 15528 29300
rect 16028 29248 16080 29300
rect 17408 29248 17460 29300
rect 18696 29248 18748 29300
rect 20444 29248 20496 29300
rect 20628 29291 20680 29300
rect 20628 29257 20637 29291
rect 20637 29257 20671 29291
rect 20671 29257 20680 29291
rect 20628 29248 20680 29257
rect 15568 29180 15620 29232
rect 22284 29248 22336 29300
rect 22376 29248 22428 29300
rect 21456 29180 21508 29232
rect 22560 29248 22612 29300
rect 15844 29112 15896 29164
rect 17776 29112 17828 29164
rect 18052 29155 18104 29164
rect 18052 29121 18061 29155
rect 18061 29121 18095 29155
rect 18095 29121 18104 29155
rect 18052 29112 18104 29121
rect 18236 29112 18288 29164
rect 19248 29112 19300 29164
rect 19892 29155 19944 29164
rect 19892 29121 19901 29155
rect 19901 29121 19935 29155
rect 19935 29121 19944 29155
rect 19892 29112 19944 29121
rect 14372 29044 14424 29096
rect 16764 29044 16816 29096
rect 17040 29044 17092 29096
rect 20076 29155 20128 29164
rect 20076 29121 20085 29155
rect 20085 29121 20119 29155
rect 20119 29121 20128 29155
rect 20076 29112 20128 29121
rect 20444 29112 20496 29164
rect 20720 29112 20772 29164
rect 9956 29019 10008 29028
rect 9956 28985 9965 29019
rect 9965 28985 9999 29019
rect 9999 28985 10008 29019
rect 9956 28976 10008 28985
rect 11336 28976 11388 29028
rect 14740 28976 14792 29028
rect 15568 28976 15620 29028
rect 16212 29019 16264 29028
rect 13636 28908 13688 28960
rect 14188 28908 14240 28960
rect 15752 28951 15804 28960
rect 15752 28917 15761 28951
rect 15761 28917 15795 28951
rect 15795 28917 15804 28951
rect 15752 28908 15804 28917
rect 16212 28985 16221 29019
rect 16221 28985 16255 29019
rect 16255 28985 16264 29019
rect 16212 28976 16264 28985
rect 17224 28976 17276 29028
rect 18788 28976 18840 29028
rect 20260 28976 20312 29028
rect 22744 29112 22796 29164
rect 23296 29155 23348 29164
rect 23296 29121 23305 29155
rect 23305 29121 23339 29155
rect 23339 29121 23348 29155
rect 23296 29112 23348 29121
rect 23664 29155 23716 29164
rect 23664 29121 23673 29155
rect 23673 29121 23707 29155
rect 23707 29121 23716 29155
rect 23664 29112 23716 29121
rect 21088 28976 21140 29028
rect 22192 28976 22244 29028
rect 22284 28976 22336 29028
rect 23296 29019 23348 29028
rect 23296 28985 23305 29019
rect 23305 28985 23339 29019
rect 23339 28985 23348 29019
rect 23296 28976 23348 28985
rect 24032 29112 24084 29164
rect 24308 29112 24360 29164
rect 24676 29155 24728 29164
rect 24676 29121 24685 29155
rect 24685 29121 24719 29155
rect 24719 29121 24728 29155
rect 25228 29180 25280 29232
rect 26332 29248 26384 29300
rect 27988 29248 28040 29300
rect 28264 29248 28316 29300
rect 28448 29248 28500 29300
rect 28632 29248 28684 29300
rect 30196 29291 30248 29300
rect 25872 29180 25924 29232
rect 24676 29112 24728 29121
rect 24952 29155 25004 29164
rect 24952 29121 24961 29155
rect 24961 29121 24995 29155
rect 24995 29121 25004 29155
rect 24952 29112 25004 29121
rect 25136 29112 25188 29164
rect 23572 28976 23624 29028
rect 23664 28976 23716 29028
rect 24032 28976 24084 29028
rect 24400 29044 24452 29096
rect 25228 29044 25280 29096
rect 25688 29112 25740 29164
rect 26516 29112 26568 29164
rect 26332 29044 26384 29096
rect 26976 29112 27028 29164
rect 27528 29180 27580 29232
rect 30196 29257 30205 29291
rect 30205 29257 30239 29291
rect 30239 29257 30248 29291
rect 30196 29248 30248 29257
rect 26792 29044 26844 29096
rect 24308 28976 24360 29028
rect 26148 28976 26200 29028
rect 26424 28976 26476 29028
rect 26700 28976 26752 29028
rect 27068 28976 27120 29028
rect 27620 29044 27672 29096
rect 27712 29044 27764 29096
rect 27436 28976 27488 29028
rect 24400 28908 24452 28960
rect 25320 28908 25372 28960
rect 26516 28908 26568 28960
rect 26792 28908 26844 28960
rect 26976 28908 27028 28960
rect 27252 28908 27304 28960
rect 27620 28908 27672 28960
rect 28356 29112 28408 29164
rect 28448 29112 28500 29164
rect 32404 29180 32456 29232
rect 28632 29044 28684 29096
rect 29460 29112 29512 29164
rect 29828 29112 29880 29164
rect 30012 29155 30064 29164
rect 30012 29121 30021 29155
rect 30021 29121 30055 29155
rect 30055 29121 30064 29155
rect 30012 29112 30064 29121
rect 30380 29112 30432 29164
rect 32864 29044 32916 29096
rect 28908 28976 28960 29028
rect 29368 28976 29420 29028
rect 29736 28976 29788 29028
rect 31208 29019 31260 29028
rect 31208 28985 31217 29019
rect 31217 28985 31251 29019
rect 31251 28985 31260 29019
rect 31208 28976 31260 28985
rect 28816 28908 28868 28960
rect 29184 28908 29236 28960
rect 30196 28908 30248 28960
rect 4791 28806 4843 28858
rect 4855 28806 4907 28858
rect 4919 28806 4971 28858
rect 4983 28806 5035 28858
rect 5047 28806 5099 28858
rect 12473 28806 12525 28858
rect 12537 28806 12589 28858
rect 12601 28806 12653 28858
rect 12665 28806 12717 28858
rect 12729 28806 12781 28858
rect 20155 28806 20207 28858
rect 20219 28806 20271 28858
rect 20283 28806 20335 28858
rect 20347 28806 20399 28858
rect 20411 28806 20463 28858
rect 27837 28806 27889 28858
rect 27901 28806 27953 28858
rect 27965 28806 28017 28858
rect 28029 28806 28081 28858
rect 28093 28806 28145 28858
rect 9864 28747 9916 28756
rect 9864 28713 9873 28747
rect 9873 28713 9907 28747
rect 9907 28713 9916 28747
rect 9864 28704 9916 28713
rect 11796 28704 11848 28756
rect 12072 28704 12124 28756
rect 6368 28636 6420 28688
rect 12440 28636 12492 28688
rect 13820 28704 13872 28756
rect 16028 28704 16080 28756
rect 17132 28747 17184 28756
rect 17132 28713 17141 28747
rect 17141 28713 17175 28747
rect 17175 28713 17184 28747
rect 17132 28704 17184 28713
rect 17408 28704 17460 28756
rect 18052 28704 18104 28756
rect 18512 28704 18564 28756
rect 20260 28704 20312 28756
rect 20536 28704 20588 28756
rect 21548 28704 21600 28756
rect 22008 28704 22060 28756
rect 17592 28679 17644 28688
rect 17592 28645 17601 28679
rect 17601 28645 17635 28679
rect 17635 28645 17644 28679
rect 17592 28636 17644 28645
rect 17776 28636 17828 28688
rect 21824 28636 21876 28688
rect 23112 28704 23164 28756
rect 23204 28704 23256 28756
rect 23388 28704 23440 28756
rect 23480 28704 23532 28756
rect 22928 28636 22980 28688
rect 23572 28636 23624 28688
rect 19708 28568 19760 28620
rect 1584 28543 1636 28552
rect 1584 28509 1593 28543
rect 1593 28509 1627 28543
rect 1627 28509 1636 28543
rect 1584 28500 1636 28509
rect 9036 28500 9088 28552
rect 4160 28364 4212 28416
rect 11060 28500 11112 28552
rect 13176 28543 13228 28552
rect 13176 28509 13185 28543
rect 13185 28509 13219 28543
rect 13219 28509 13228 28543
rect 13176 28500 13228 28509
rect 14188 28432 14240 28484
rect 15752 28432 15804 28484
rect 9404 28364 9456 28416
rect 10416 28407 10468 28416
rect 10416 28373 10425 28407
rect 10425 28373 10459 28407
rect 10459 28373 10468 28407
rect 10416 28364 10468 28373
rect 10876 28364 10928 28416
rect 11520 28407 11572 28416
rect 11520 28373 11529 28407
rect 11529 28373 11563 28407
rect 11563 28373 11572 28407
rect 11520 28364 11572 28373
rect 15200 28407 15252 28416
rect 15200 28373 15209 28407
rect 15209 28373 15243 28407
rect 15243 28373 15252 28407
rect 15200 28364 15252 28373
rect 15292 28364 15344 28416
rect 16856 28432 16908 28484
rect 18236 28500 18288 28552
rect 18696 28543 18748 28552
rect 18696 28509 18705 28543
rect 18705 28509 18739 28543
rect 18739 28509 18748 28543
rect 18696 28500 18748 28509
rect 20444 28568 20496 28620
rect 19340 28432 19392 28484
rect 19984 28500 20036 28552
rect 20720 28568 20772 28620
rect 20812 28568 20864 28620
rect 23756 28704 23808 28756
rect 25596 28704 25648 28756
rect 25780 28747 25832 28756
rect 25780 28713 25789 28747
rect 25789 28713 25823 28747
rect 25823 28713 25832 28747
rect 25780 28704 25832 28713
rect 25872 28704 25924 28756
rect 26516 28704 26568 28756
rect 26884 28704 26936 28756
rect 26976 28747 27028 28756
rect 26976 28713 26985 28747
rect 26985 28713 27019 28747
rect 27019 28713 27028 28747
rect 26976 28704 27028 28713
rect 24584 28636 24636 28688
rect 24952 28636 25004 28688
rect 25044 28636 25096 28688
rect 21916 28500 21968 28552
rect 22192 28543 22244 28552
rect 22192 28509 22201 28543
rect 22201 28509 22235 28543
rect 22235 28509 22244 28543
rect 22192 28500 22244 28509
rect 20352 28475 20404 28484
rect 20352 28441 20361 28475
rect 20361 28441 20395 28475
rect 20395 28441 20404 28475
rect 20352 28432 20404 28441
rect 20444 28432 20496 28484
rect 21180 28432 21232 28484
rect 21456 28432 21508 28484
rect 22560 28500 22612 28552
rect 24124 28568 24176 28620
rect 24216 28568 24268 28620
rect 25320 28568 25372 28620
rect 25596 28568 25648 28620
rect 25780 28568 25832 28620
rect 26792 28636 26844 28688
rect 31392 28704 31444 28756
rect 30012 28636 30064 28688
rect 16672 28364 16724 28416
rect 17960 28364 18012 28416
rect 19616 28364 19668 28416
rect 20720 28364 20772 28416
rect 20812 28364 20864 28416
rect 21364 28364 21416 28416
rect 21548 28364 21600 28416
rect 22100 28364 22152 28416
rect 22284 28364 22336 28416
rect 22744 28432 22796 28484
rect 24584 28500 24636 28552
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 25412 28500 25464 28552
rect 23940 28432 23992 28484
rect 24124 28432 24176 28484
rect 25780 28432 25832 28484
rect 23039 28407 23091 28416
rect 23039 28373 23063 28407
rect 23063 28373 23091 28407
rect 23039 28364 23091 28373
rect 23572 28407 23624 28416
rect 23572 28373 23581 28407
rect 23581 28373 23615 28407
rect 23615 28373 23624 28407
rect 23572 28364 23624 28373
rect 23756 28364 23808 28416
rect 25688 28364 25740 28416
rect 25872 28364 25924 28416
rect 26240 28500 26292 28552
rect 26792 28543 26844 28552
rect 26792 28509 26801 28543
rect 26801 28509 26835 28543
rect 26835 28509 26844 28543
rect 26792 28500 26844 28509
rect 27804 28500 27856 28552
rect 28264 28500 28316 28552
rect 29092 28568 29144 28620
rect 29460 28500 29512 28552
rect 30012 28500 30064 28552
rect 27712 28475 27764 28484
rect 27712 28441 27721 28475
rect 27721 28441 27755 28475
rect 27755 28441 27764 28475
rect 27712 28432 27764 28441
rect 27896 28475 27948 28484
rect 27896 28441 27905 28475
rect 27905 28441 27939 28475
rect 27939 28441 27948 28475
rect 27896 28432 27948 28441
rect 26884 28364 26936 28416
rect 27068 28364 27120 28416
rect 27620 28364 27672 28416
rect 28264 28364 28316 28416
rect 29184 28432 29236 28484
rect 30564 28500 30616 28552
rect 31300 28500 31352 28552
rect 32404 28432 32456 28484
rect 28540 28364 28592 28416
rect 29000 28364 29052 28416
rect 29092 28364 29144 28416
rect 29460 28364 29512 28416
rect 29828 28407 29880 28416
rect 29828 28373 29837 28407
rect 29837 28373 29871 28407
rect 29871 28373 29880 28407
rect 29828 28364 29880 28373
rect 30380 28364 30432 28416
rect 31300 28364 31352 28416
rect 8632 28262 8684 28314
rect 8696 28262 8748 28314
rect 8760 28262 8812 28314
rect 8824 28262 8876 28314
rect 8888 28262 8940 28314
rect 16314 28262 16366 28314
rect 16378 28262 16430 28314
rect 16442 28262 16494 28314
rect 16506 28262 16558 28314
rect 16570 28262 16622 28314
rect 23996 28262 24048 28314
rect 24060 28262 24112 28314
rect 24124 28262 24176 28314
rect 24188 28262 24240 28314
rect 24252 28262 24304 28314
rect 31678 28262 31730 28314
rect 31742 28262 31794 28314
rect 31806 28262 31858 28314
rect 31870 28262 31922 28314
rect 31934 28262 31986 28314
rect 9588 28160 9640 28212
rect 14556 28160 14608 28212
rect 14740 28203 14792 28212
rect 14740 28169 14749 28203
rect 14749 28169 14783 28203
rect 14783 28169 14792 28203
rect 14740 28160 14792 28169
rect 15384 28160 15436 28212
rect 15936 28160 15988 28212
rect 18604 28160 18656 28212
rect 18696 28160 18748 28212
rect 19156 28160 19208 28212
rect 19340 28160 19392 28212
rect 19616 28160 19668 28212
rect 21180 28160 21232 28212
rect 21824 28160 21876 28212
rect 11428 28092 11480 28144
rect 11980 28092 12032 28144
rect 12808 28135 12860 28144
rect 12808 28101 12817 28135
rect 12817 28101 12851 28135
rect 12851 28101 12860 28135
rect 12808 28092 12860 28101
rect 13268 28135 13320 28144
rect 13268 28101 13277 28135
rect 13277 28101 13311 28135
rect 13311 28101 13320 28135
rect 13268 28092 13320 28101
rect 14924 28092 14976 28144
rect 16580 28092 16632 28144
rect 17224 28135 17276 28144
rect 17224 28101 17233 28135
rect 17233 28101 17267 28135
rect 17267 28101 17276 28135
rect 17224 28092 17276 28101
rect 13360 28024 13412 28076
rect 10508 27956 10560 28008
rect 13912 27956 13964 28008
rect 14372 27956 14424 28008
rect 14556 27956 14608 28008
rect 18788 28024 18840 28076
rect 18978 28067 19030 28076
rect 18978 28033 18981 28067
rect 18981 28033 19015 28067
rect 19015 28033 19030 28067
rect 18978 28024 19030 28033
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 19156 28024 19208 28033
rect 19340 28024 19392 28076
rect 20260 28024 20312 28076
rect 20536 28024 20588 28076
rect 8300 27888 8352 27940
rect 11336 27888 11388 27940
rect 11796 27888 11848 27940
rect 11980 27888 12032 27940
rect 15292 27888 15344 27940
rect 15752 27888 15804 27940
rect 19616 27956 19668 28008
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 8116 27820 8168 27872
rect 8392 27863 8444 27872
rect 8392 27829 8401 27863
rect 8401 27829 8435 27863
rect 8435 27829 8444 27863
rect 8392 27820 8444 27829
rect 9680 27820 9732 27872
rect 11244 27820 11296 27872
rect 12072 27820 12124 27872
rect 12808 27820 12860 27872
rect 15108 27820 15160 27872
rect 15660 27820 15712 27872
rect 19800 27888 19852 27940
rect 20076 27956 20128 28008
rect 22192 28135 22244 28144
rect 22192 28101 22201 28135
rect 22201 28101 22235 28135
rect 22235 28101 22244 28135
rect 22192 28092 22244 28101
rect 22284 28092 22336 28144
rect 23480 28160 23532 28212
rect 23664 28160 23716 28212
rect 24216 28160 24268 28212
rect 20812 28024 20864 28076
rect 20904 27956 20956 28008
rect 21640 28024 21692 28076
rect 22744 28024 22796 28076
rect 23572 28092 23624 28144
rect 23940 28092 23992 28144
rect 27988 28160 28040 28212
rect 28172 28203 28224 28212
rect 28172 28169 28181 28203
rect 28181 28169 28215 28203
rect 28215 28169 28224 28203
rect 28172 28160 28224 28169
rect 21824 27956 21876 28008
rect 23020 28067 23072 28076
rect 23020 28033 23048 28067
rect 23048 28033 23072 28067
rect 23204 28067 23256 28076
rect 23020 28024 23072 28033
rect 23204 28033 23213 28067
rect 23213 28033 23247 28067
rect 23247 28033 23256 28067
rect 23204 28024 23256 28033
rect 24400 28135 24452 28144
rect 24400 28101 24409 28135
rect 24409 28101 24443 28135
rect 24443 28101 24452 28135
rect 24400 28092 24452 28101
rect 25412 28092 25464 28144
rect 24124 28024 24176 28076
rect 24952 28024 25004 28076
rect 25228 28067 25280 28076
rect 25228 28033 25237 28067
rect 25237 28033 25271 28067
rect 25271 28033 25280 28067
rect 25228 28024 25280 28033
rect 26608 28092 26660 28144
rect 26700 28092 26752 28144
rect 26052 28067 26104 28076
rect 21272 27888 21324 27940
rect 22560 27888 22612 27940
rect 24400 27956 24452 28008
rect 24584 27956 24636 28008
rect 26052 28033 26061 28067
rect 26061 28033 26095 28067
rect 26095 28033 26104 28067
rect 26052 28024 26104 28033
rect 26148 28067 26200 28076
rect 26148 28033 26157 28067
rect 26157 28033 26191 28067
rect 26191 28033 26200 28067
rect 26148 28024 26200 28033
rect 26792 28024 26844 28076
rect 26976 28024 27028 28076
rect 27620 28024 27672 28076
rect 28080 28024 28132 28076
rect 28356 28067 28408 28076
rect 28356 28033 28365 28067
rect 28365 28033 28399 28067
rect 28399 28033 28408 28067
rect 28356 28024 28408 28033
rect 28816 28092 28868 28144
rect 29276 28135 29328 28144
rect 29276 28101 29285 28135
rect 29285 28101 29319 28135
rect 29319 28101 29328 28135
rect 29276 28092 29328 28101
rect 29460 28135 29512 28144
rect 29460 28101 29469 28135
rect 29469 28101 29503 28135
rect 29503 28101 29512 28135
rect 29460 28092 29512 28101
rect 30748 28092 30800 28144
rect 25412 27956 25464 28008
rect 19064 27820 19116 27872
rect 22192 27820 22244 27872
rect 24216 27888 24268 27940
rect 24860 27820 24912 27872
rect 25228 27863 25280 27872
rect 25228 27829 25237 27863
rect 25237 27829 25271 27863
rect 25271 27829 25280 27863
rect 25228 27820 25280 27829
rect 25596 27820 25648 27872
rect 25780 27888 25832 27940
rect 26608 27956 26660 28008
rect 27804 27956 27856 28008
rect 26884 27888 26936 27940
rect 26700 27820 26752 27872
rect 26792 27820 26844 27872
rect 27436 27820 27488 27872
rect 28448 27863 28500 27872
rect 28448 27829 28457 27863
rect 28457 27829 28491 27863
rect 28491 27829 28500 27863
rect 28448 27820 28500 27829
rect 29552 28024 29604 28076
rect 30012 28024 30064 28076
rect 30104 28024 30156 28076
rect 28816 27956 28868 28008
rect 30288 27956 30340 28008
rect 29828 27888 29880 27940
rect 30196 27888 30248 27940
rect 31024 28067 31076 28076
rect 31024 28033 31033 28067
rect 31033 28033 31067 28067
rect 31067 28033 31076 28067
rect 31024 28024 31076 28033
rect 31024 27888 31076 27940
rect 29460 27820 29512 27872
rect 30288 27820 30340 27872
rect 4791 27718 4843 27770
rect 4855 27718 4907 27770
rect 4919 27718 4971 27770
rect 4983 27718 5035 27770
rect 5047 27718 5099 27770
rect 12473 27718 12525 27770
rect 12537 27718 12589 27770
rect 12601 27718 12653 27770
rect 12665 27718 12717 27770
rect 12729 27718 12781 27770
rect 20155 27718 20207 27770
rect 20219 27718 20271 27770
rect 20283 27718 20335 27770
rect 20347 27718 20399 27770
rect 20411 27718 20463 27770
rect 27837 27718 27889 27770
rect 27901 27718 27953 27770
rect 27965 27718 28017 27770
rect 28029 27718 28081 27770
rect 28093 27718 28145 27770
rect 8392 27616 8444 27668
rect 12992 27616 13044 27668
rect 14372 27616 14424 27668
rect 15384 27616 15436 27668
rect 15752 27616 15804 27668
rect 16580 27616 16632 27668
rect 16948 27616 17000 27668
rect 17408 27616 17460 27668
rect 17500 27659 17552 27668
rect 17500 27625 17509 27659
rect 17509 27625 17543 27659
rect 17543 27625 17552 27659
rect 17500 27616 17552 27625
rect 17868 27616 17920 27668
rect 9036 27548 9088 27600
rect 10048 27548 10100 27600
rect 11796 27548 11848 27600
rect 10140 27480 10192 27532
rect 10324 27523 10376 27532
rect 10324 27489 10333 27523
rect 10333 27489 10367 27523
rect 10367 27489 10376 27523
rect 10324 27480 10376 27489
rect 10416 27480 10468 27532
rect 12900 27548 12952 27600
rect 13636 27548 13688 27600
rect 17960 27548 18012 27600
rect 18328 27548 18380 27600
rect 18420 27548 18472 27600
rect 20260 27616 20312 27668
rect 20812 27616 20864 27668
rect 21272 27616 21324 27668
rect 21548 27616 21600 27668
rect 21640 27616 21692 27668
rect 19340 27548 19392 27600
rect 20076 27548 20128 27600
rect 11244 27412 11296 27464
rect 12164 27412 12216 27464
rect 13544 27480 13596 27532
rect 17040 27480 17092 27532
rect 17592 27480 17644 27532
rect 14188 27412 14240 27464
rect 16120 27412 16172 27464
rect 17132 27412 17184 27464
rect 3884 27344 3936 27396
rect 7380 27387 7432 27396
rect 7380 27353 7389 27387
rect 7389 27353 7423 27387
rect 7423 27353 7432 27387
rect 7380 27344 7432 27353
rect 8024 27387 8076 27396
rect 8024 27353 8033 27387
rect 8033 27353 8067 27387
rect 8067 27353 8076 27387
rect 8024 27344 8076 27353
rect 10324 27344 10376 27396
rect 12072 27387 12124 27396
rect 12072 27353 12081 27387
rect 12081 27353 12115 27387
rect 12115 27353 12124 27387
rect 12072 27344 12124 27353
rect 14004 27344 14056 27396
rect 14832 27344 14884 27396
rect 15660 27344 15712 27396
rect 18236 27412 18288 27464
rect 18420 27412 18472 27464
rect 18696 27455 18748 27464
rect 18696 27421 18705 27455
rect 18705 27421 18739 27455
rect 18739 27421 18748 27455
rect 18696 27412 18748 27421
rect 17592 27344 17644 27396
rect 19340 27412 19392 27464
rect 19892 27455 19944 27464
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 20260 27412 20312 27464
rect 20720 27523 20772 27532
rect 20720 27489 20729 27523
rect 20729 27489 20763 27523
rect 20763 27489 20772 27523
rect 20720 27480 20772 27489
rect 21272 27523 21324 27532
rect 21272 27489 21281 27523
rect 21281 27489 21315 27523
rect 21315 27489 21324 27523
rect 21272 27480 21324 27489
rect 20168 27344 20220 27396
rect 6368 27319 6420 27328
rect 6368 27285 6377 27319
rect 6377 27285 6411 27319
rect 6411 27285 6420 27319
rect 6368 27276 6420 27285
rect 7288 27276 7340 27328
rect 9036 27276 9088 27328
rect 9404 27276 9456 27328
rect 11612 27276 11664 27328
rect 11888 27276 11940 27328
rect 16764 27276 16816 27328
rect 16856 27276 16908 27328
rect 20720 27276 20772 27328
rect 20904 27276 20956 27328
rect 21088 27412 21140 27464
rect 23296 27548 23348 27600
rect 23572 27616 23624 27668
rect 24860 27616 24912 27668
rect 25596 27616 25648 27668
rect 26148 27616 26200 27668
rect 22744 27480 22796 27532
rect 24584 27480 24636 27532
rect 23204 27412 23256 27464
rect 21272 27344 21324 27396
rect 21640 27276 21692 27328
rect 22192 27344 22244 27396
rect 22284 27344 22336 27396
rect 22836 27344 22888 27396
rect 22928 27276 22980 27328
rect 23572 27276 23624 27328
rect 24216 27412 24268 27464
rect 26240 27591 26292 27600
rect 26240 27557 26249 27591
rect 26249 27557 26283 27591
rect 26283 27557 26292 27591
rect 26240 27548 26292 27557
rect 26884 27548 26936 27600
rect 26976 27548 27028 27600
rect 29092 27616 29144 27668
rect 29644 27616 29696 27668
rect 30564 27616 30616 27668
rect 25228 27455 25280 27464
rect 23940 27344 23992 27396
rect 25228 27421 25237 27455
rect 25237 27421 25271 27455
rect 25271 27421 25280 27455
rect 25228 27412 25280 27421
rect 25504 27412 25556 27464
rect 25964 27412 26016 27464
rect 26148 27412 26200 27464
rect 27620 27480 27672 27532
rect 26332 27344 26384 27396
rect 24032 27276 24084 27328
rect 24860 27276 24912 27328
rect 25320 27276 25372 27328
rect 25688 27276 25740 27328
rect 26608 27344 26660 27396
rect 27528 27412 27580 27464
rect 28724 27480 28776 27532
rect 28816 27480 28868 27532
rect 29000 27480 29052 27532
rect 27620 27344 27672 27396
rect 27804 27344 27856 27396
rect 28172 27455 28224 27464
rect 28172 27421 28193 27455
rect 28193 27421 28224 27455
rect 28172 27412 28224 27421
rect 29092 27387 29144 27396
rect 26976 27276 27028 27328
rect 27068 27319 27120 27328
rect 27068 27285 27077 27319
rect 27077 27285 27111 27319
rect 27111 27285 27120 27319
rect 29092 27353 29101 27387
rect 29101 27353 29135 27387
rect 29135 27353 29144 27387
rect 29092 27344 29144 27353
rect 28724 27319 28776 27328
rect 27068 27276 27120 27285
rect 28724 27285 28733 27319
rect 28733 27285 28767 27319
rect 28767 27285 28776 27319
rect 28724 27276 28776 27285
rect 28908 27319 28960 27328
rect 28908 27285 28935 27319
rect 28935 27285 28960 27319
rect 28908 27276 28960 27285
rect 29552 27480 29604 27532
rect 30564 27523 30616 27532
rect 29828 27344 29880 27396
rect 30564 27489 30573 27523
rect 30573 27489 30607 27523
rect 30607 27489 30616 27523
rect 30564 27480 30616 27489
rect 30196 27412 30248 27464
rect 8632 27174 8684 27226
rect 8696 27174 8748 27226
rect 8760 27174 8812 27226
rect 8824 27174 8876 27226
rect 8888 27174 8940 27226
rect 16314 27174 16366 27226
rect 16378 27174 16430 27226
rect 16442 27174 16494 27226
rect 16506 27174 16558 27226
rect 16570 27174 16622 27226
rect 23996 27174 24048 27226
rect 24060 27174 24112 27226
rect 24124 27174 24176 27226
rect 24188 27174 24240 27226
rect 24252 27174 24304 27226
rect 31678 27174 31730 27226
rect 31742 27174 31794 27226
rect 31806 27174 31858 27226
rect 31870 27174 31922 27226
rect 31934 27174 31986 27226
rect 8484 27072 8536 27124
rect 9588 27072 9640 27124
rect 10048 27115 10100 27124
rect 10048 27081 10057 27115
rect 10057 27081 10091 27115
rect 10091 27081 10100 27115
rect 10048 27072 10100 27081
rect 11060 27072 11112 27124
rect 13268 27072 13320 27124
rect 15292 27072 15344 27124
rect 15660 27115 15712 27124
rect 15660 27081 15669 27115
rect 15669 27081 15703 27115
rect 15703 27081 15712 27115
rect 15660 27072 15712 27081
rect 6276 27004 6328 27056
rect 10324 27004 10376 27056
rect 11796 27004 11848 27056
rect 16028 27004 16080 27056
rect 16488 27004 16540 27056
rect 16764 27004 16816 27056
rect 17132 27004 17184 27056
rect 9128 26936 9180 26988
rect 17040 26936 17092 26988
rect 17316 26936 17368 26988
rect 18236 27004 18288 27056
rect 19892 27072 19944 27124
rect 18052 26936 18104 26988
rect 19064 26936 19116 26988
rect 19156 26936 19208 26988
rect 19616 26936 19668 26988
rect 20168 27004 20220 27056
rect 21364 27072 21416 27124
rect 22928 27072 22980 27124
rect 23376 27072 23428 27124
rect 23480 27072 23532 27124
rect 24032 27115 24084 27124
rect 24032 27081 24041 27115
rect 24041 27081 24075 27115
rect 24075 27081 24084 27115
rect 24032 27072 24084 27081
rect 9496 26868 9548 26920
rect 14188 26868 14240 26920
rect 17500 26868 17552 26920
rect 18236 26868 18288 26920
rect 18604 26911 18656 26920
rect 18604 26877 18613 26911
rect 18613 26877 18647 26911
rect 18647 26877 18656 26911
rect 18604 26868 18656 26877
rect 18972 26868 19024 26920
rect 11612 26800 11664 26852
rect 11980 26800 12032 26852
rect 15384 26800 15436 26852
rect 7288 26775 7340 26784
rect 7288 26741 7297 26775
rect 7297 26741 7331 26775
rect 7331 26741 7340 26775
rect 7288 26732 7340 26741
rect 9588 26732 9640 26784
rect 10508 26775 10560 26784
rect 10508 26741 10517 26775
rect 10517 26741 10551 26775
rect 10551 26741 10560 26775
rect 10508 26732 10560 26741
rect 10876 26732 10928 26784
rect 12992 26775 13044 26784
rect 12992 26741 13001 26775
rect 13001 26741 13035 26775
rect 13035 26741 13044 26775
rect 12992 26732 13044 26741
rect 13452 26775 13504 26784
rect 13452 26741 13461 26775
rect 13461 26741 13495 26775
rect 13495 26741 13504 26775
rect 13452 26732 13504 26741
rect 13636 26732 13688 26784
rect 15108 26732 15160 26784
rect 15292 26732 15344 26784
rect 16212 26800 16264 26852
rect 17040 26800 17092 26852
rect 17316 26800 17368 26852
rect 16580 26732 16632 26784
rect 17132 26732 17184 26784
rect 17960 26732 18012 26784
rect 18328 26800 18380 26852
rect 18785 26775 18837 26784
rect 18785 26741 18797 26775
rect 18797 26741 18831 26775
rect 18831 26741 18837 26775
rect 19432 26775 19484 26784
rect 18785 26732 18837 26741
rect 19432 26741 19441 26775
rect 19441 26741 19475 26775
rect 19475 26741 19484 26775
rect 19432 26732 19484 26741
rect 19616 26732 19668 26784
rect 19892 26732 19944 26784
rect 20076 26732 20128 26784
rect 20536 26800 20588 26852
rect 21364 26936 21416 26988
rect 21456 26936 21508 26988
rect 22192 26936 22244 26988
rect 22560 26979 22612 26988
rect 22560 26945 22569 26979
rect 22569 26945 22603 26979
rect 22603 26945 22612 26979
rect 22560 26936 22612 26945
rect 21548 26868 21600 26920
rect 22100 26800 22152 26852
rect 22284 26868 22336 26920
rect 23664 27004 23716 27056
rect 23940 27004 23992 27056
rect 26148 27072 26200 27124
rect 27896 27072 27948 27124
rect 27988 27072 28040 27124
rect 28356 27115 28408 27124
rect 28356 27081 28365 27115
rect 28365 27081 28399 27115
rect 28399 27081 28408 27115
rect 28356 27072 28408 27081
rect 22928 26979 22980 26988
rect 22928 26945 22937 26979
rect 22937 26945 22971 26979
rect 22971 26945 22980 26979
rect 22928 26936 22980 26945
rect 23204 26936 23256 26988
rect 23480 26936 23532 26988
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 24400 26936 24452 26988
rect 23296 26868 23348 26920
rect 23388 26868 23440 26920
rect 23848 26911 23900 26920
rect 23848 26877 23857 26911
rect 23857 26877 23891 26911
rect 23891 26877 23900 26911
rect 24124 26911 24176 26920
rect 23848 26868 23900 26877
rect 24124 26877 24133 26911
rect 24133 26877 24167 26911
rect 24167 26877 24176 26911
rect 24124 26868 24176 26877
rect 24308 26868 24360 26920
rect 25320 26979 25372 26988
rect 25320 26945 25362 26979
rect 25362 26945 25372 26979
rect 25320 26936 25372 26945
rect 25504 26979 25556 26988
rect 25504 26945 25513 26979
rect 25513 26945 25547 26979
rect 25547 26945 25556 26979
rect 25504 26936 25556 26945
rect 26332 26979 26384 26988
rect 26332 26945 26341 26979
rect 26341 26945 26375 26979
rect 26375 26945 26384 26979
rect 26332 26936 26384 26945
rect 26424 26979 26476 26988
rect 26424 26945 26433 26979
rect 26433 26945 26467 26979
rect 26467 26945 26476 26979
rect 26424 26936 26476 26945
rect 26884 26936 26936 26988
rect 23020 26800 23072 26852
rect 23204 26800 23256 26852
rect 20444 26732 20496 26784
rect 22560 26732 22612 26784
rect 23388 26732 23440 26784
rect 23572 26800 23624 26852
rect 24400 26800 24452 26852
rect 25872 26800 25924 26852
rect 26792 26868 26844 26920
rect 28816 27004 28868 27056
rect 29276 27004 29328 27056
rect 27252 26936 27304 26988
rect 27528 26979 27580 26988
rect 27528 26945 27537 26979
rect 27537 26945 27571 26979
rect 27571 26945 27580 26979
rect 27528 26936 27580 26945
rect 27712 26979 27764 26988
rect 27712 26945 27721 26979
rect 27721 26945 27755 26979
rect 27755 26945 27764 26979
rect 27712 26936 27764 26945
rect 27896 26936 27948 26988
rect 28540 26936 28592 26988
rect 28908 26936 28960 26988
rect 29368 26936 29420 26988
rect 29552 26979 29604 26988
rect 29552 26945 29561 26979
rect 29561 26945 29595 26979
rect 29595 26945 29604 26979
rect 29552 26936 29604 26945
rect 29828 27072 29880 27124
rect 30196 27072 30248 27124
rect 30472 27115 30524 27124
rect 30472 27081 30481 27115
rect 30481 27081 30515 27115
rect 30515 27081 30524 27115
rect 30472 27072 30524 27081
rect 31484 27072 31536 27124
rect 30104 27047 30156 27056
rect 30104 27013 30113 27047
rect 30113 27013 30147 27047
rect 30147 27013 30156 27047
rect 30104 27004 30156 27013
rect 31024 27004 31076 27056
rect 31668 27004 31720 27056
rect 30196 26936 30248 26988
rect 31208 26936 31260 26988
rect 29368 26843 29420 26852
rect 29368 26809 29377 26843
rect 29377 26809 29411 26843
rect 29411 26809 29420 26843
rect 29368 26800 29420 26809
rect 31760 26868 31812 26920
rect 30932 26800 30984 26852
rect 25596 26732 25648 26784
rect 26240 26732 26292 26784
rect 26792 26732 26844 26784
rect 26884 26732 26936 26784
rect 27068 26732 27120 26784
rect 27528 26732 27580 26784
rect 27896 26732 27948 26784
rect 28080 26732 28132 26784
rect 28173 26732 28225 26784
rect 28724 26732 28776 26784
rect 29276 26732 29328 26784
rect 29828 26732 29880 26784
rect 4791 26630 4843 26682
rect 4855 26630 4907 26682
rect 4919 26630 4971 26682
rect 4983 26630 5035 26682
rect 5047 26630 5099 26682
rect 12473 26630 12525 26682
rect 12537 26630 12589 26682
rect 12601 26630 12653 26682
rect 12665 26630 12717 26682
rect 12729 26630 12781 26682
rect 20155 26630 20207 26682
rect 20219 26630 20271 26682
rect 20283 26630 20335 26682
rect 20347 26630 20399 26682
rect 20411 26630 20463 26682
rect 27837 26630 27889 26682
rect 27901 26630 27953 26682
rect 27965 26630 28017 26682
rect 28029 26630 28081 26682
rect 28093 26630 28145 26682
rect 10968 26528 11020 26580
rect 12256 26528 12308 26580
rect 12348 26528 12400 26580
rect 13084 26571 13136 26580
rect 10600 26460 10652 26512
rect 11612 26460 11664 26512
rect 13084 26537 13093 26571
rect 13093 26537 13127 26571
rect 13127 26537 13136 26571
rect 13084 26528 13136 26537
rect 13268 26528 13320 26580
rect 13636 26528 13688 26580
rect 14648 26571 14700 26580
rect 14648 26537 14657 26571
rect 14657 26537 14691 26571
rect 14691 26537 14700 26571
rect 14648 26528 14700 26537
rect 5172 26392 5224 26444
rect 11796 26392 11848 26444
rect 12256 26392 12308 26444
rect 16212 26528 16264 26580
rect 16856 26528 16908 26580
rect 17040 26528 17092 26580
rect 17592 26528 17644 26580
rect 17868 26528 17920 26580
rect 20536 26528 20588 26580
rect 15292 26460 15344 26512
rect 16580 26460 16632 26512
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 9312 26367 9364 26376
rect 9312 26333 9321 26367
rect 9321 26333 9355 26367
rect 9355 26333 9364 26367
rect 9312 26324 9364 26333
rect 9404 26324 9456 26376
rect 12900 26324 12952 26376
rect 15936 26367 15988 26376
rect 6828 26256 6880 26308
rect 7932 26299 7984 26308
rect 7472 26231 7524 26240
rect 7472 26197 7481 26231
rect 7481 26197 7515 26231
rect 7515 26197 7524 26231
rect 7472 26188 7524 26197
rect 7932 26265 7941 26299
rect 7941 26265 7975 26299
rect 7975 26265 7984 26299
rect 7932 26256 7984 26265
rect 9772 26299 9824 26308
rect 9772 26265 9781 26299
rect 9781 26265 9815 26299
rect 9815 26265 9824 26299
rect 9772 26256 9824 26265
rect 12072 26299 12124 26308
rect 12072 26265 12081 26299
rect 12081 26265 12115 26299
rect 12115 26265 12124 26299
rect 12072 26256 12124 26265
rect 14464 26256 14516 26308
rect 15108 26256 15160 26308
rect 15660 26256 15712 26308
rect 15936 26333 15945 26367
rect 15945 26333 15979 26367
rect 15979 26333 15988 26367
rect 15936 26324 15988 26333
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 16580 26367 16632 26376
rect 16580 26333 16589 26367
rect 16589 26333 16623 26367
rect 16623 26333 16632 26367
rect 16580 26324 16632 26333
rect 16672 26324 16724 26376
rect 17408 26392 17460 26444
rect 17592 26392 17644 26444
rect 17868 26392 17920 26444
rect 18236 26460 18288 26512
rect 19616 26460 19668 26512
rect 15844 26256 15896 26308
rect 16488 26256 16540 26308
rect 17040 26367 17092 26376
rect 17040 26333 17050 26367
rect 17050 26333 17084 26367
rect 17084 26333 17092 26367
rect 17040 26324 17092 26333
rect 18236 26324 18288 26376
rect 18420 26324 18472 26376
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 19156 26324 19208 26376
rect 19708 26324 19760 26376
rect 19984 26324 20036 26376
rect 20076 26367 20128 26376
rect 20076 26333 20085 26367
rect 20085 26333 20119 26367
rect 20119 26333 20128 26367
rect 20628 26460 20680 26512
rect 20352 26392 20404 26444
rect 22008 26528 22060 26580
rect 21180 26460 21232 26512
rect 25044 26528 25096 26580
rect 25596 26528 25648 26580
rect 20076 26324 20128 26333
rect 21180 26324 21232 26376
rect 23112 26460 23164 26512
rect 22192 26392 22244 26444
rect 22560 26392 22612 26444
rect 17408 26256 17460 26308
rect 19892 26256 19944 26308
rect 22560 26256 22612 26308
rect 23480 26460 23532 26512
rect 23388 26392 23440 26444
rect 23572 26367 23624 26376
rect 23572 26333 23581 26367
rect 23581 26333 23615 26367
rect 23615 26333 23624 26367
rect 23572 26324 23624 26333
rect 12348 26188 12400 26240
rect 12716 26188 12768 26240
rect 13636 26231 13688 26240
rect 13636 26197 13645 26231
rect 13645 26197 13679 26231
rect 13679 26197 13688 26231
rect 13636 26188 13688 26197
rect 17040 26188 17092 26240
rect 17132 26188 17184 26240
rect 18144 26188 18196 26240
rect 18604 26188 18656 26240
rect 19064 26188 19116 26240
rect 21364 26188 21416 26240
rect 21916 26188 21968 26240
rect 22376 26188 22428 26240
rect 23480 26299 23532 26308
rect 23480 26265 23489 26299
rect 23489 26265 23523 26299
rect 23523 26265 23532 26299
rect 23480 26256 23532 26265
rect 22744 26188 22796 26240
rect 25688 26460 25740 26512
rect 26424 26460 26476 26512
rect 26700 26460 26752 26512
rect 25872 26392 25924 26444
rect 23848 26324 23900 26376
rect 23940 26324 23992 26376
rect 25136 26324 25188 26376
rect 24584 26299 24636 26308
rect 24584 26265 24593 26299
rect 24593 26265 24627 26299
rect 24627 26265 24636 26299
rect 24584 26256 24636 26265
rect 24676 26188 24728 26240
rect 25688 26324 25740 26376
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 26424 26367 26476 26376
rect 26424 26333 26433 26367
rect 26433 26333 26467 26367
rect 26467 26333 26476 26367
rect 26424 26324 26476 26333
rect 26608 26324 26660 26376
rect 27068 26367 27120 26376
rect 27068 26333 27077 26367
rect 27077 26333 27111 26367
rect 27111 26333 27120 26367
rect 27068 26324 27120 26333
rect 27160 26367 27212 26376
rect 27160 26333 27172 26367
rect 27172 26333 27206 26367
rect 27206 26333 27212 26367
rect 27528 26435 27580 26444
rect 27528 26401 27537 26435
rect 27537 26401 27571 26435
rect 27571 26401 27580 26435
rect 27528 26392 27580 26401
rect 27712 26392 27764 26444
rect 28908 26528 28960 26580
rect 29368 26528 29420 26580
rect 30932 26571 30984 26580
rect 30932 26537 30941 26571
rect 30941 26537 30975 26571
rect 30975 26537 30984 26571
rect 30932 26528 30984 26537
rect 28264 26460 28316 26512
rect 29000 26460 29052 26512
rect 29552 26460 29604 26512
rect 29828 26460 29880 26512
rect 30104 26460 30156 26512
rect 30840 26460 30892 26512
rect 28080 26392 28132 26444
rect 27160 26324 27212 26333
rect 27896 26324 27948 26376
rect 28172 26367 28224 26376
rect 28172 26333 28181 26367
rect 28181 26333 28215 26367
rect 28215 26333 28224 26367
rect 28172 26324 28224 26333
rect 28724 26324 28776 26376
rect 29000 26367 29052 26376
rect 29000 26333 29009 26367
rect 29009 26333 29043 26367
rect 29043 26333 29052 26367
rect 29000 26324 29052 26333
rect 29092 26367 29144 26376
rect 29092 26333 29101 26367
rect 29101 26333 29135 26367
rect 29135 26333 29144 26367
rect 29092 26324 29144 26333
rect 29368 26324 29420 26376
rect 31208 26392 31260 26444
rect 30840 26367 30892 26376
rect 27988 26256 28040 26308
rect 29828 26256 29880 26308
rect 30840 26333 30849 26367
rect 30849 26333 30883 26367
rect 30883 26333 30892 26367
rect 30840 26324 30892 26333
rect 31484 26324 31536 26376
rect 31852 26256 31904 26308
rect 25780 26188 25832 26240
rect 29092 26188 29144 26240
rect 30840 26188 30892 26240
rect 30932 26188 30984 26240
rect 31668 26188 31720 26240
rect 31760 26188 31812 26240
rect 8632 26086 8684 26138
rect 8696 26086 8748 26138
rect 8760 26086 8812 26138
rect 8824 26086 8876 26138
rect 8888 26086 8940 26138
rect 16314 26086 16366 26138
rect 16378 26086 16430 26138
rect 16442 26086 16494 26138
rect 16506 26086 16558 26138
rect 16570 26086 16622 26138
rect 23996 26086 24048 26138
rect 24060 26086 24112 26138
rect 24124 26086 24176 26138
rect 24188 26086 24240 26138
rect 24252 26086 24304 26138
rect 31678 26086 31730 26138
rect 31742 26086 31794 26138
rect 31806 26086 31858 26138
rect 31870 26086 31922 26138
rect 31934 26086 31986 26138
rect 32128 26120 32180 26172
rect 7932 25984 7984 26036
rect 11888 25984 11940 26036
rect 11152 25959 11204 25968
rect 11152 25925 11161 25959
rect 11161 25925 11195 25959
rect 11195 25925 11204 25959
rect 11152 25916 11204 25925
rect 11428 25916 11480 25968
rect 13544 25848 13596 25900
rect 8576 25780 8628 25832
rect 10600 25780 10652 25832
rect 12164 25780 12216 25832
rect 13084 25780 13136 25832
rect 13728 25984 13780 26036
rect 13912 25984 13964 26036
rect 16488 25984 16540 26036
rect 18696 25984 18748 26036
rect 13728 25848 13780 25900
rect 14832 25891 14884 25900
rect 14832 25857 14841 25891
rect 14841 25857 14875 25891
rect 14875 25857 14884 25891
rect 14832 25848 14884 25857
rect 15016 25891 15068 25900
rect 15016 25857 15025 25891
rect 15025 25857 15059 25891
rect 15059 25857 15068 25891
rect 15016 25848 15068 25857
rect 15292 25848 15344 25900
rect 16212 25848 16264 25900
rect 16396 25848 16448 25900
rect 16856 25848 16908 25900
rect 13912 25780 13964 25832
rect 16672 25780 16724 25832
rect 16764 25780 16816 25832
rect 16948 25780 17000 25832
rect 7656 25712 7708 25764
rect 9312 25712 9364 25764
rect 11796 25712 11848 25764
rect 14372 25712 14424 25764
rect 17224 25712 17276 25764
rect 18236 25916 18288 25968
rect 17592 25848 17644 25900
rect 18420 25848 18472 25900
rect 18236 25780 18288 25832
rect 18880 25848 18932 25900
rect 19255 25858 19307 25910
rect 19064 25780 19116 25832
rect 19616 25848 19668 25900
rect 20076 25891 20128 25900
rect 7472 25644 7524 25696
rect 8116 25644 8168 25696
rect 12164 25644 12216 25696
rect 13452 25644 13504 25696
rect 14280 25687 14332 25696
rect 14280 25653 14289 25687
rect 14289 25653 14323 25687
rect 14323 25653 14332 25687
rect 14280 25644 14332 25653
rect 14648 25644 14700 25696
rect 16396 25644 16448 25696
rect 17408 25644 17460 25696
rect 17684 25687 17736 25696
rect 17684 25653 17693 25687
rect 17693 25653 17727 25687
rect 17727 25653 17736 25687
rect 17684 25644 17736 25653
rect 17868 25644 17920 25696
rect 18236 25644 18288 25696
rect 18604 25712 18656 25764
rect 19248 25712 19300 25764
rect 19708 25780 19760 25832
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 21364 25916 21416 25968
rect 21732 25916 21784 25968
rect 22744 25984 22796 26036
rect 25044 25984 25096 26036
rect 25596 25984 25648 26036
rect 28908 25984 28960 26036
rect 29184 25984 29236 26036
rect 20260 25891 20312 25900
rect 20260 25857 20269 25891
rect 20269 25857 20303 25891
rect 20303 25857 20312 25891
rect 20260 25848 20312 25857
rect 20444 25848 20496 25900
rect 19432 25644 19484 25696
rect 19524 25644 19576 25696
rect 20444 25712 20496 25764
rect 20628 25712 20680 25764
rect 20812 25712 20864 25764
rect 19800 25644 19852 25696
rect 21272 25780 21324 25832
rect 21732 25780 21784 25832
rect 22192 25848 22244 25900
rect 24492 25916 24544 25968
rect 25688 25916 25740 25968
rect 26516 25916 26568 25968
rect 23112 25848 23164 25900
rect 26056 25848 26108 25900
rect 27068 25848 27120 25900
rect 27712 25916 27764 25968
rect 30380 25984 30432 26036
rect 30748 26027 30800 26036
rect 30748 25993 30757 26027
rect 30757 25993 30791 26027
rect 30791 25993 30800 26027
rect 30748 25984 30800 25993
rect 29644 25916 29696 25968
rect 22376 25712 22428 25764
rect 21732 25644 21784 25696
rect 21916 25644 21968 25696
rect 22192 25644 22244 25696
rect 22560 25780 22612 25832
rect 24032 25780 24084 25832
rect 24768 25780 24820 25832
rect 25964 25780 26016 25832
rect 26148 25780 26200 25832
rect 26516 25780 26568 25832
rect 27528 25891 27580 25900
rect 27528 25857 27537 25891
rect 27537 25857 27571 25891
rect 27571 25857 27580 25891
rect 27528 25848 27580 25857
rect 28816 25848 28868 25900
rect 29828 25891 29880 25900
rect 27620 25780 27672 25832
rect 27712 25780 27764 25832
rect 29184 25780 29236 25832
rect 25872 25712 25924 25764
rect 27160 25712 27212 25764
rect 27436 25712 27488 25764
rect 27804 25712 27856 25764
rect 24676 25644 24728 25696
rect 25412 25644 25464 25696
rect 25964 25644 26016 25696
rect 26148 25644 26200 25696
rect 28356 25712 28408 25764
rect 29276 25712 29328 25764
rect 29828 25857 29837 25891
rect 29837 25857 29871 25891
rect 29871 25857 29880 25891
rect 29828 25848 29880 25857
rect 30380 25891 30432 25900
rect 30380 25857 30389 25891
rect 30389 25857 30423 25891
rect 30423 25857 30432 25891
rect 30380 25848 30432 25857
rect 30932 25848 30984 25900
rect 29736 25823 29788 25832
rect 29736 25789 29745 25823
rect 29745 25789 29779 25823
rect 29779 25789 29788 25823
rect 29736 25780 29788 25789
rect 29644 25712 29696 25764
rect 31208 25780 31260 25832
rect 30932 25712 30984 25764
rect 30472 25644 30524 25696
rect 30748 25644 30800 25696
rect 31208 25687 31260 25696
rect 31208 25653 31217 25687
rect 31217 25653 31251 25687
rect 31251 25653 31260 25687
rect 31208 25644 31260 25653
rect 4791 25542 4843 25594
rect 4855 25542 4907 25594
rect 4919 25542 4971 25594
rect 4983 25542 5035 25594
rect 5047 25542 5099 25594
rect 12473 25542 12525 25594
rect 12537 25542 12589 25594
rect 12601 25542 12653 25594
rect 12665 25542 12717 25594
rect 12729 25542 12781 25594
rect 20155 25542 20207 25594
rect 20219 25542 20271 25594
rect 20283 25542 20335 25594
rect 20347 25542 20399 25594
rect 20411 25542 20463 25594
rect 27837 25542 27889 25594
rect 27901 25542 27953 25594
rect 27965 25542 28017 25594
rect 28029 25542 28081 25594
rect 28093 25542 28145 25594
rect 6276 25483 6328 25492
rect 6276 25449 6285 25483
rect 6285 25449 6319 25483
rect 6319 25449 6328 25483
rect 6276 25440 6328 25449
rect 6368 25440 6420 25492
rect 8484 25440 8536 25492
rect 11244 25440 11296 25492
rect 11612 25440 11664 25492
rect 11888 25483 11940 25492
rect 11888 25449 11897 25483
rect 11897 25449 11931 25483
rect 11931 25449 11940 25483
rect 11888 25440 11940 25449
rect 13636 25483 13688 25492
rect 13636 25449 13645 25483
rect 13645 25449 13679 25483
rect 13679 25449 13688 25483
rect 13636 25440 13688 25449
rect 6828 25372 6880 25424
rect 7472 25372 7524 25424
rect 12808 25372 12860 25424
rect 9036 25304 9088 25356
rect 11612 25304 11664 25356
rect 14464 25440 14516 25492
rect 13912 25372 13964 25424
rect 14280 25372 14332 25424
rect 15200 25440 15252 25492
rect 16764 25483 16816 25492
rect 16764 25449 16773 25483
rect 16773 25449 16807 25483
rect 16807 25449 16816 25483
rect 16764 25440 16816 25449
rect 17132 25483 17184 25492
rect 17132 25449 17141 25483
rect 17141 25449 17175 25483
rect 17175 25449 17184 25483
rect 17132 25440 17184 25449
rect 17224 25440 17276 25492
rect 17500 25440 17552 25492
rect 17776 25440 17828 25492
rect 18420 25440 18472 25492
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 11796 25236 11848 25288
rect 13176 25236 13228 25288
rect 14740 25304 14792 25356
rect 13636 25236 13688 25288
rect 14464 25236 14516 25288
rect 10600 25168 10652 25220
rect 12900 25168 12952 25220
rect 5816 25143 5868 25152
rect 5816 25109 5825 25143
rect 5825 25109 5859 25143
rect 5859 25109 5868 25143
rect 5816 25100 5868 25109
rect 9864 25100 9916 25152
rect 11428 25143 11480 25152
rect 11428 25109 11437 25143
rect 11437 25109 11471 25143
rect 11471 25109 11480 25143
rect 11428 25100 11480 25109
rect 11796 25100 11848 25152
rect 13176 25100 13228 25152
rect 15568 25236 15620 25288
rect 15936 25372 15988 25424
rect 16488 25372 16540 25424
rect 16580 25372 16632 25424
rect 17316 25372 17368 25424
rect 16212 25304 16264 25356
rect 20168 25440 20220 25492
rect 21180 25483 21232 25492
rect 21180 25449 21189 25483
rect 21189 25449 21223 25483
rect 21223 25449 21232 25483
rect 21180 25440 21232 25449
rect 13636 25100 13688 25152
rect 15200 25100 15252 25152
rect 15660 25100 15712 25152
rect 17316 25236 17368 25288
rect 17500 25236 17552 25288
rect 17868 25168 17920 25220
rect 19156 25304 19208 25356
rect 18328 25236 18380 25288
rect 18512 25279 18564 25288
rect 18512 25245 18547 25279
rect 18547 25245 18564 25279
rect 18512 25236 18564 25245
rect 18788 25236 18840 25288
rect 19340 25304 19392 25356
rect 19984 25372 20036 25424
rect 20444 25372 20496 25424
rect 20536 25372 20588 25424
rect 21364 25372 21416 25424
rect 21548 25440 21600 25492
rect 23664 25440 23716 25492
rect 23940 25440 23992 25492
rect 24124 25440 24176 25492
rect 24860 25440 24912 25492
rect 24952 25440 25004 25492
rect 21272 25304 21324 25356
rect 22008 25372 22060 25424
rect 22284 25372 22336 25424
rect 23756 25372 23808 25424
rect 24584 25372 24636 25424
rect 25964 25372 26016 25424
rect 26424 25440 26476 25492
rect 27988 25440 28040 25492
rect 29644 25440 29696 25492
rect 29736 25440 29788 25492
rect 30932 25483 30984 25492
rect 22652 25304 22704 25356
rect 23112 25304 23164 25356
rect 23204 25304 23256 25356
rect 25228 25304 25280 25356
rect 27068 25372 27120 25424
rect 27252 25372 27304 25424
rect 19432 25279 19484 25288
rect 19432 25245 19441 25279
rect 19441 25245 19475 25279
rect 19475 25245 19484 25279
rect 19432 25236 19484 25245
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 20352 25279 20404 25288
rect 19524 25236 19576 25245
rect 20352 25245 20361 25279
rect 20361 25245 20395 25279
rect 20395 25245 20404 25279
rect 20352 25236 20404 25245
rect 18236 25168 18288 25220
rect 16764 25100 16816 25152
rect 17408 25100 17460 25152
rect 18052 25100 18104 25152
rect 18604 25100 18656 25152
rect 18788 25100 18840 25152
rect 19340 25168 19392 25220
rect 19616 25168 19668 25220
rect 19892 25168 19944 25220
rect 20536 25168 20588 25220
rect 20720 25100 20772 25152
rect 20904 25236 20956 25288
rect 20996 25168 21048 25220
rect 22284 25279 22336 25288
rect 22284 25245 22293 25279
rect 22293 25245 22327 25279
rect 22327 25245 22336 25279
rect 22284 25236 22336 25245
rect 24308 25236 24360 25288
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 22652 25168 22704 25220
rect 21364 25100 21416 25152
rect 21548 25100 21600 25152
rect 22008 25100 22060 25152
rect 23204 25100 23256 25152
rect 23572 25100 23624 25152
rect 24216 25100 24268 25152
rect 24860 25100 24912 25152
rect 25136 25100 25188 25152
rect 26424 25100 26476 25152
rect 26976 25236 27028 25288
rect 27160 25279 27212 25288
rect 27160 25245 27169 25279
rect 27169 25245 27203 25279
rect 27203 25245 27212 25279
rect 27160 25236 27212 25245
rect 27252 25279 27304 25288
rect 27252 25245 27261 25279
rect 27261 25245 27295 25279
rect 27295 25245 27304 25279
rect 27804 25304 27856 25356
rect 30564 25372 30616 25424
rect 30380 25304 30432 25356
rect 27252 25236 27304 25245
rect 27712 25236 27764 25288
rect 28172 25236 28224 25288
rect 26700 25168 26752 25220
rect 28264 25168 28316 25220
rect 28816 25236 28868 25288
rect 29828 25236 29880 25288
rect 30104 25236 30156 25288
rect 30564 25236 30616 25288
rect 30932 25449 30941 25483
rect 30941 25449 30975 25483
rect 30975 25449 30984 25483
rect 30932 25440 30984 25449
rect 30840 25372 30892 25424
rect 29184 25211 29236 25220
rect 29184 25177 29193 25211
rect 29193 25177 29227 25211
rect 29227 25177 29236 25211
rect 29184 25168 29236 25177
rect 29736 25143 29788 25152
rect 29736 25109 29745 25143
rect 29745 25109 29779 25143
rect 29779 25109 29788 25143
rect 29736 25100 29788 25109
rect 30840 25100 30892 25152
rect 8632 24998 8684 25050
rect 8696 24998 8748 25050
rect 8760 24998 8812 25050
rect 8824 24998 8876 25050
rect 8888 24998 8940 25050
rect 16314 24998 16366 25050
rect 16378 24998 16430 25050
rect 16442 24998 16494 25050
rect 16506 24998 16558 25050
rect 16570 24998 16622 25050
rect 23996 24998 24048 25050
rect 24060 24998 24112 25050
rect 24124 24998 24176 25050
rect 24188 24998 24240 25050
rect 24252 24998 24304 25050
rect 31678 24998 31730 25050
rect 31742 24998 31794 25050
rect 31806 24998 31858 25050
rect 31870 24998 31922 25050
rect 31934 24998 31986 25050
rect 11428 24896 11480 24948
rect 12164 24896 12216 24948
rect 13360 24896 13412 24948
rect 14740 24896 14792 24948
rect 4252 24828 4304 24880
rect 5172 24760 5224 24812
rect 8392 24760 8444 24812
rect 9312 24760 9364 24812
rect 9588 24760 9640 24812
rect 12900 24828 12952 24880
rect 14832 24828 14884 24880
rect 4344 24692 4396 24744
rect 10232 24692 10284 24744
rect 12716 24760 12768 24812
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 14280 24760 14332 24812
rect 15384 24828 15436 24880
rect 15660 24896 15712 24948
rect 20168 24896 20220 24948
rect 20536 24896 20588 24948
rect 20996 24896 21048 24948
rect 15936 24871 15988 24880
rect 12900 24692 12952 24744
rect 12992 24692 13044 24744
rect 13360 24692 13412 24744
rect 15568 24760 15620 24812
rect 15384 24692 15436 24744
rect 15936 24837 15945 24871
rect 15945 24837 15979 24871
rect 15979 24837 15988 24871
rect 15936 24828 15988 24837
rect 16120 24871 16172 24880
rect 16120 24837 16161 24871
rect 16161 24837 16172 24871
rect 16120 24828 16172 24837
rect 16580 24828 16632 24880
rect 17776 24828 17828 24880
rect 16764 24760 16816 24812
rect 17224 24760 17276 24812
rect 18788 24828 18840 24880
rect 18052 24760 18104 24812
rect 18144 24760 18196 24812
rect 18604 24760 18656 24812
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 19248 24828 19300 24880
rect 18972 24760 19024 24769
rect 19800 24760 19852 24812
rect 20076 24828 20128 24880
rect 21916 24896 21968 24948
rect 22284 24896 22336 24948
rect 24584 24896 24636 24948
rect 24952 24896 25004 24948
rect 26516 24896 26568 24948
rect 26700 24896 26752 24948
rect 23572 24828 23624 24880
rect 23848 24828 23900 24880
rect 25044 24828 25096 24880
rect 6000 24667 6052 24676
rect 6000 24633 6009 24667
rect 6009 24633 6043 24667
rect 6043 24633 6052 24667
rect 6000 24624 6052 24633
rect 7748 24599 7800 24608
rect 7748 24565 7757 24599
rect 7757 24565 7791 24599
rect 7791 24565 7800 24599
rect 7748 24556 7800 24565
rect 9772 24624 9824 24676
rect 14740 24624 14792 24676
rect 15936 24624 15988 24676
rect 16488 24624 16540 24676
rect 17408 24624 17460 24676
rect 18880 24735 18932 24744
rect 18052 24624 18104 24676
rect 18880 24701 18889 24735
rect 18889 24701 18923 24735
rect 18923 24701 18932 24735
rect 18880 24692 18932 24701
rect 19708 24692 19760 24744
rect 8484 24556 8536 24608
rect 8944 24599 8996 24608
rect 8944 24565 8953 24599
rect 8953 24565 8987 24599
rect 8987 24565 8996 24599
rect 8944 24556 8996 24565
rect 9680 24556 9732 24608
rect 10232 24556 10284 24608
rect 11060 24556 11112 24608
rect 11888 24556 11940 24608
rect 12256 24556 12308 24608
rect 14464 24556 14516 24608
rect 16028 24556 16080 24608
rect 16856 24556 16908 24608
rect 17592 24556 17644 24608
rect 17960 24556 18012 24608
rect 19248 24624 19300 24676
rect 22100 24760 22152 24812
rect 25596 24803 25648 24812
rect 20168 24692 20220 24744
rect 21088 24735 21140 24744
rect 21088 24701 21097 24735
rect 21097 24701 21131 24735
rect 21131 24701 21140 24735
rect 21088 24692 21140 24701
rect 19156 24556 19208 24608
rect 19708 24556 19760 24608
rect 19800 24556 19852 24608
rect 21272 24624 21324 24676
rect 21548 24692 21600 24744
rect 21824 24692 21876 24744
rect 25596 24769 25605 24803
rect 25605 24769 25639 24803
rect 25639 24769 25648 24803
rect 25596 24760 25648 24769
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 23020 24692 23072 24744
rect 23112 24692 23164 24744
rect 21824 24556 21876 24608
rect 22468 24556 22520 24608
rect 22652 24599 22704 24608
rect 22652 24565 22661 24599
rect 22661 24565 22695 24599
rect 22695 24565 22704 24599
rect 22652 24556 22704 24565
rect 22928 24624 22980 24676
rect 25044 24692 25096 24744
rect 26792 24828 26844 24880
rect 26516 24760 26568 24812
rect 26976 24828 27028 24880
rect 27228 24828 27280 24880
rect 27620 24896 27672 24948
rect 28816 24896 28868 24948
rect 29092 24896 29144 24948
rect 30840 24896 30892 24948
rect 31116 24828 31168 24880
rect 31484 24828 31536 24880
rect 27068 24760 27120 24812
rect 27712 24760 27764 24812
rect 28172 24760 28224 24812
rect 28448 24760 28500 24812
rect 24676 24624 24728 24676
rect 27988 24692 28040 24744
rect 28724 24803 28776 24812
rect 28724 24769 28733 24803
rect 28733 24769 28767 24803
rect 28767 24769 28776 24803
rect 28724 24760 28776 24769
rect 29276 24760 29328 24812
rect 29736 24760 29788 24812
rect 29828 24803 29880 24812
rect 29828 24769 29862 24803
rect 29862 24769 29880 24803
rect 29828 24760 29880 24769
rect 30380 24760 30432 24812
rect 30012 24692 30064 24744
rect 30748 24803 30800 24812
rect 30748 24769 30757 24803
rect 30757 24769 30791 24803
rect 30791 24769 30800 24803
rect 30748 24760 30800 24769
rect 30932 24803 30984 24812
rect 30932 24769 30941 24803
rect 30941 24769 30975 24803
rect 30975 24769 30984 24803
rect 30932 24760 30984 24769
rect 32220 24760 32272 24812
rect 24308 24556 24360 24608
rect 25044 24599 25096 24608
rect 25044 24565 25053 24599
rect 25053 24565 25087 24599
rect 25087 24565 25096 24599
rect 25044 24556 25096 24565
rect 25780 24556 25832 24608
rect 27252 24556 27304 24608
rect 27528 24556 27580 24608
rect 27712 24599 27764 24608
rect 27712 24565 27721 24599
rect 27721 24565 27755 24599
rect 27755 24565 27764 24599
rect 27712 24556 27764 24565
rect 29736 24624 29788 24676
rect 32496 24692 32548 24744
rect 30840 24667 30892 24676
rect 30840 24633 30849 24667
rect 30849 24633 30883 24667
rect 30883 24633 30892 24667
rect 30840 24624 30892 24633
rect 28448 24556 28500 24608
rect 29276 24556 29328 24608
rect 32588 24556 32640 24608
rect 4791 24454 4843 24506
rect 4855 24454 4907 24506
rect 4919 24454 4971 24506
rect 4983 24454 5035 24506
rect 5047 24454 5099 24506
rect 12473 24454 12525 24506
rect 12537 24454 12589 24506
rect 12601 24454 12653 24506
rect 12665 24454 12717 24506
rect 12729 24454 12781 24506
rect 20155 24454 20207 24506
rect 20219 24454 20271 24506
rect 20283 24454 20335 24506
rect 20347 24454 20399 24506
rect 20411 24454 20463 24506
rect 27837 24454 27889 24506
rect 27901 24454 27953 24506
rect 27965 24454 28017 24506
rect 28029 24454 28081 24506
rect 28093 24454 28145 24506
rect 4160 24395 4212 24404
rect 4160 24361 4169 24395
rect 4169 24361 4203 24395
rect 4203 24361 4212 24395
rect 4160 24352 4212 24361
rect 6920 24352 6972 24404
rect 8484 24352 8536 24404
rect 10232 24352 10284 24404
rect 11796 24352 11848 24404
rect 5816 24327 5868 24336
rect 5816 24293 5825 24327
rect 5825 24293 5859 24327
rect 5859 24293 5868 24327
rect 5816 24284 5868 24293
rect 8944 24216 8996 24268
rect 9588 24216 9640 24268
rect 9680 24216 9732 24268
rect 10232 24216 10284 24268
rect 11888 24216 11940 24268
rect 13544 24284 13596 24336
rect 13912 24284 13964 24336
rect 14740 24395 14792 24404
rect 14740 24361 14749 24395
rect 14749 24361 14783 24395
rect 14783 24361 14792 24395
rect 14740 24352 14792 24361
rect 15016 24352 15068 24404
rect 15752 24395 15804 24404
rect 15752 24361 15761 24395
rect 15761 24361 15795 24395
rect 15795 24361 15804 24395
rect 15752 24352 15804 24361
rect 15936 24352 15988 24404
rect 16212 24284 16264 24336
rect 18420 24352 18472 24404
rect 20352 24352 20404 24404
rect 18696 24327 18748 24336
rect 10140 24191 10192 24200
rect 5908 24080 5960 24132
rect 5632 24012 5684 24064
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 11704 24148 11756 24200
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 6920 24123 6972 24132
rect 6920 24089 6929 24123
rect 6929 24089 6963 24123
rect 6963 24089 6972 24123
rect 6920 24080 6972 24089
rect 7656 24080 7708 24132
rect 8484 24123 8536 24132
rect 8484 24089 8493 24123
rect 8493 24089 8527 24123
rect 8527 24089 8536 24123
rect 8484 24080 8536 24089
rect 9588 24080 9640 24132
rect 13728 24216 13780 24268
rect 16396 24259 16448 24268
rect 13360 24148 13412 24200
rect 13912 24148 13964 24200
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 16764 24216 16816 24268
rect 18696 24293 18705 24327
rect 18705 24293 18739 24327
rect 18739 24293 18748 24327
rect 18696 24284 18748 24293
rect 19156 24284 19208 24336
rect 21456 24352 21508 24404
rect 21732 24352 21784 24404
rect 22928 24352 22980 24404
rect 24400 24352 24452 24404
rect 25044 24352 25096 24404
rect 26700 24352 26752 24404
rect 21824 24284 21876 24336
rect 22284 24259 22336 24268
rect 7748 24012 7800 24064
rect 9404 24012 9456 24064
rect 10968 24012 11020 24064
rect 12256 24012 12308 24064
rect 14004 24080 14056 24132
rect 14280 24080 14332 24132
rect 14372 24080 14424 24132
rect 13360 24012 13412 24064
rect 13912 24012 13964 24064
rect 14096 24012 14148 24064
rect 16304 24148 16356 24200
rect 16856 24148 16908 24200
rect 17316 24148 17368 24200
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 15568 24123 15620 24132
rect 15568 24089 15577 24123
rect 15577 24089 15611 24123
rect 15611 24089 15620 24123
rect 15568 24080 15620 24089
rect 15660 24080 15712 24132
rect 16948 24080 17000 24132
rect 15016 24012 15068 24064
rect 16672 24012 16724 24064
rect 17408 24012 17460 24064
rect 22284 24225 22293 24259
rect 22293 24225 22327 24259
rect 22327 24225 22336 24259
rect 22284 24216 22336 24225
rect 23572 24284 23624 24336
rect 24492 24284 24544 24336
rect 25872 24284 25924 24336
rect 27620 24352 27672 24404
rect 28264 24352 28316 24404
rect 28908 24352 28960 24404
rect 31024 24395 31076 24404
rect 31024 24361 31033 24395
rect 31033 24361 31067 24395
rect 31067 24361 31076 24395
rect 31024 24352 31076 24361
rect 29184 24327 29236 24336
rect 29184 24293 29193 24327
rect 29193 24293 29227 24327
rect 29227 24293 29236 24327
rect 29184 24284 29236 24293
rect 29920 24284 29972 24336
rect 31208 24284 31260 24336
rect 22928 24216 22980 24268
rect 25412 24216 25464 24268
rect 28724 24216 28776 24268
rect 28908 24216 28960 24268
rect 29644 24216 29696 24268
rect 31024 24259 31076 24268
rect 17960 24148 18012 24200
rect 18144 24148 18196 24200
rect 18328 24148 18380 24200
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 18880 24148 18932 24200
rect 18972 24148 19024 24200
rect 19340 24148 19392 24200
rect 19524 24148 19576 24200
rect 19984 24148 20036 24200
rect 20076 24148 20128 24200
rect 20260 24148 20312 24200
rect 22100 24148 22152 24200
rect 23664 24148 23716 24200
rect 24584 24191 24636 24200
rect 24584 24157 24593 24191
rect 24593 24157 24627 24191
rect 24627 24157 24636 24191
rect 24584 24148 24636 24157
rect 25964 24148 26016 24200
rect 17868 24012 17920 24064
rect 19248 24012 19300 24064
rect 19340 24012 19392 24064
rect 19708 24012 19760 24064
rect 19892 24012 19944 24064
rect 21088 24080 21140 24132
rect 21272 24080 21324 24132
rect 22836 24080 22888 24132
rect 23572 24012 23624 24064
rect 25044 24012 25096 24064
rect 26240 24012 26292 24064
rect 28540 24080 28592 24132
rect 27804 24012 27856 24064
rect 29828 24148 29880 24200
rect 31024 24225 31033 24259
rect 31033 24225 31067 24259
rect 31067 24225 31076 24259
rect 31024 24216 31076 24225
rect 29184 24080 29236 24132
rect 29460 24080 29512 24132
rect 30748 24148 30800 24200
rect 30840 24123 30892 24132
rect 30840 24089 30849 24123
rect 30849 24089 30883 24123
rect 30883 24089 30892 24123
rect 30840 24080 30892 24089
rect 28724 24012 28776 24064
rect 29736 24012 29788 24064
rect 29828 24012 29880 24064
rect 31576 24012 31628 24064
rect 8632 23910 8684 23962
rect 8696 23910 8748 23962
rect 8760 23910 8812 23962
rect 8824 23910 8876 23962
rect 8888 23910 8940 23962
rect 16314 23910 16366 23962
rect 16378 23910 16430 23962
rect 16442 23910 16494 23962
rect 16506 23910 16558 23962
rect 16570 23910 16622 23962
rect 23996 23910 24048 23962
rect 24060 23910 24112 23962
rect 24124 23910 24176 23962
rect 24188 23910 24240 23962
rect 24252 23910 24304 23962
rect 31678 23910 31730 23962
rect 31742 23910 31794 23962
rect 31806 23910 31858 23962
rect 31870 23910 31922 23962
rect 31934 23910 31986 23962
rect 4344 23851 4396 23860
rect 4344 23817 4353 23851
rect 4353 23817 4387 23851
rect 4387 23817 4396 23851
rect 4344 23808 4396 23817
rect 7012 23808 7064 23860
rect 7288 23851 7340 23860
rect 7288 23817 7297 23851
rect 7297 23817 7331 23851
rect 7331 23817 7340 23851
rect 7288 23808 7340 23817
rect 9404 23808 9456 23860
rect 10876 23808 10928 23860
rect 12164 23851 12216 23860
rect 10508 23740 10560 23792
rect 11152 23740 11204 23792
rect 12164 23817 12173 23851
rect 12173 23817 12207 23851
rect 12207 23817 12216 23851
rect 12164 23808 12216 23817
rect 15384 23851 15436 23860
rect 15384 23817 15393 23851
rect 15393 23817 15427 23851
rect 15427 23817 15436 23851
rect 15384 23808 15436 23817
rect 15476 23808 15528 23860
rect 10416 23672 10468 23724
rect 11060 23672 11112 23724
rect 11428 23672 11480 23724
rect 12348 23715 12400 23724
rect 12348 23681 12357 23715
rect 12357 23681 12391 23715
rect 12391 23681 12400 23715
rect 12348 23672 12400 23681
rect 1584 23647 1636 23656
rect 1584 23613 1593 23647
rect 1593 23613 1627 23647
rect 1627 23613 1636 23647
rect 1584 23604 1636 23613
rect 7104 23604 7156 23656
rect 9956 23647 10008 23656
rect 9956 23613 9965 23647
rect 9965 23613 9999 23647
rect 9999 23613 10008 23647
rect 9956 23604 10008 23613
rect 11152 23604 11204 23656
rect 14096 23740 14148 23792
rect 14280 23740 14332 23792
rect 14556 23740 14608 23792
rect 15660 23740 15712 23792
rect 13452 23715 13504 23724
rect 5356 23536 5408 23588
rect 7840 23511 7892 23520
rect 7840 23477 7849 23511
rect 7849 23477 7883 23511
rect 7883 23477 7892 23511
rect 7840 23468 7892 23477
rect 9588 23536 9640 23588
rect 13452 23681 13461 23715
rect 13461 23681 13495 23715
rect 13495 23681 13504 23715
rect 13452 23672 13504 23681
rect 14372 23672 14424 23724
rect 15108 23672 15160 23724
rect 15844 23715 15896 23724
rect 15844 23681 15853 23715
rect 15853 23681 15887 23715
rect 15887 23681 15896 23715
rect 15844 23672 15896 23681
rect 16672 23740 16724 23792
rect 16856 23740 16908 23792
rect 16120 23715 16172 23724
rect 16120 23681 16129 23715
rect 16129 23681 16163 23715
rect 16163 23681 16172 23715
rect 16120 23672 16172 23681
rect 16212 23672 16264 23724
rect 13360 23604 13412 23656
rect 14740 23604 14792 23656
rect 16764 23604 16816 23656
rect 17132 23672 17184 23724
rect 17316 23715 17368 23724
rect 17316 23681 17325 23715
rect 17325 23681 17359 23715
rect 17359 23681 17368 23715
rect 18144 23740 18196 23792
rect 18328 23740 18380 23792
rect 17316 23672 17368 23681
rect 17684 23672 17736 23724
rect 18420 23715 18472 23724
rect 18420 23681 18429 23715
rect 18429 23681 18463 23715
rect 18463 23681 18472 23715
rect 18420 23672 18472 23681
rect 19156 23740 19208 23792
rect 20628 23808 20680 23860
rect 21272 23808 21324 23860
rect 21548 23808 21600 23860
rect 22376 23808 22428 23860
rect 26884 23808 26936 23860
rect 27252 23808 27304 23860
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 14280 23536 14332 23588
rect 14832 23536 14884 23588
rect 15108 23536 15160 23588
rect 15292 23536 15344 23588
rect 16120 23536 16172 23588
rect 8852 23511 8904 23520
rect 8852 23477 8861 23511
rect 8861 23477 8895 23511
rect 8895 23477 8904 23511
rect 8852 23468 8904 23477
rect 10600 23511 10652 23520
rect 10600 23477 10609 23511
rect 10609 23477 10643 23511
rect 10643 23477 10652 23511
rect 10600 23468 10652 23477
rect 10784 23468 10836 23520
rect 11980 23468 12032 23520
rect 12164 23468 12216 23520
rect 12440 23468 12492 23520
rect 12992 23511 13044 23520
rect 12992 23477 13001 23511
rect 13001 23477 13035 23511
rect 13035 23477 13044 23511
rect 12992 23468 13044 23477
rect 13544 23511 13596 23520
rect 13544 23477 13553 23511
rect 13553 23477 13587 23511
rect 13587 23477 13596 23511
rect 13544 23468 13596 23477
rect 13636 23511 13688 23520
rect 13636 23477 13645 23511
rect 13645 23477 13679 23511
rect 13679 23477 13688 23511
rect 13636 23468 13688 23477
rect 13912 23468 13964 23520
rect 14096 23468 14148 23520
rect 14188 23468 14240 23520
rect 16396 23468 16448 23520
rect 16580 23536 16632 23588
rect 19064 23604 19116 23656
rect 19156 23604 19208 23656
rect 19248 23604 19300 23656
rect 19524 23715 19576 23724
rect 19524 23681 19533 23715
rect 19533 23681 19567 23715
rect 19567 23681 19576 23715
rect 19800 23740 19852 23792
rect 20996 23783 21048 23792
rect 19524 23672 19576 23681
rect 19898 23737 19950 23758
rect 19898 23706 19905 23737
rect 19905 23706 19939 23737
rect 19939 23706 19950 23737
rect 18144 23536 18196 23588
rect 18328 23536 18380 23588
rect 18052 23468 18104 23520
rect 19800 23536 19852 23588
rect 20996 23749 21005 23783
rect 21005 23749 21039 23783
rect 21039 23749 21048 23783
rect 20996 23740 21048 23749
rect 21364 23740 21416 23792
rect 21732 23740 21784 23792
rect 21088 23604 21140 23656
rect 21456 23604 21508 23656
rect 20260 23536 20312 23588
rect 22928 23740 22980 23792
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22468 23715 22520 23724
rect 22468 23681 22477 23715
rect 22477 23681 22511 23715
rect 22511 23681 22520 23715
rect 22468 23672 22520 23681
rect 23388 23740 23440 23792
rect 23756 23740 23808 23792
rect 24860 23740 24912 23792
rect 25688 23740 25740 23792
rect 25872 23740 25924 23792
rect 26240 23740 26292 23792
rect 26792 23740 26844 23792
rect 27528 23808 27580 23860
rect 25504 23672 25556 23724
rect 26056 23672 26108 23724
rect 22744 23604 22796 23656
rect 23480 23647 23532 23656
rect 23480 23613 23489 23647
rect 23489 23613 23523 23647
rect 23523 23613 23532 23647
rect 23480 23604 23532 23613
rect 23572 23604 23624 23656
rect 21916 23536 21968 23588
rect 22652 23536 22704 23588
rect 23204 23536 23256 23588
rect 26976 23672 27028 23724
rect 26516 23647 26568 23656
rect 26516 23613 26525 23647
rect 26525 23613 26559 23647
rect 26559 23613 26568 23647
rect 26516 23604 26568 23613
rect 26700 23604 26752 23656
rect 27712 23672 27764 23724
rect 28448 23740 28500 23792
rect 27988 23715 28040 23724
rect 27988 23681 27997 23715
rect 27997 23681 28031 23715
rect 28031 23681 28040 23715
rect 27988 23672 28040 23681
rect 28356 23672 28408 23724
rect 28540 23672 28592 23724
rect 29092 23808 29144 23860
rect 29644 23808 29696 23860
rect 30196 23808 30248 23860
rect 30656 23851 30708 23860
rect 30656 23817 30665 23851
rect 30665 23817 30699 23851
rect 30699 23817 30708 23851
rect 30656 23808 30708 23817
rect 28908 23672 28960 23724
rect 29552 23672 29604 23724
rect 30012 23715 30064 23724
rect 30012 23681 30021 23715
rect 30021 23681 30055 23715
rect 30055 23681 30064 23715
rect 30012 23672 30064 23681
rect 30564 23672 30616 23724
rect 30932 23715 30984 23724
rect 30932 23681 30941 23715
rect 30941 23681 30975 23715
rect 30975 23681 30984 23715
rect 30932 23672 30984 23681
rect 31392 23740 31444 23792
rect 32220 23672 32272 23724
rect 31300 23647 31352 23656
rect 21548 23468 21600 23520
rect 22376 23511 22428 23520
rect 22376 23477 22385 23511
rect 22385 23477 22419 23511
rect 22419 23477 22428 23511
rect 22376 23468 22428 23477
rect 22744 23511 22796 23520
rect 22744 23477 22753 23511
rect 22753 23477 22787 23511
rect 22787 23477 22796 23511
rect 22744 23468 22796 23477
rect 23112 23468 23164 23520
rect 24124 23468 24176 23520
rect 28540 23536 28592 23588
rect 28724 23536 28776 23588
rect 31300 23613 31309 23647
rect 31309 23613 31343 23647
rect 31343 23613 31352 23647
rect 31300 23604 31352 23613
rect 31392 23604 31444 23656
rect 32404 23604 32456 23656
rect 25044 23468 25096 23520
rect 25228 23468 25280 23520
rect 25320 23468 25372 23520
rect 29460 23536 29512 23588
rect 29736 23536 29788 23588
rect 30564 23536 30616 23588
rect 29368 23468 29420 23520
rect 30288 23468 30340 23520
rect 4791 23366 4843 23418
rect 4855 23366 4907 23418
rect 4919 23366 4971 23418
rect 4983 23366 5035 23418
rect 5047 23366 5099 23418
rect 12473 23366 12525 23418
rect 12537 23366 12589 23418
rect 12601 23366 12653 23418
rect 12665 23366 12717 23418
rect 12729 23366 12781 23418
rect 20155 23366 20207 23418
rect 20219 23366 20271 23418
rect 20283 23366 20335 23418
rect 20347 23366 20399 23418
rect 20411 23366 20463 23418
rect 27837 23366 27889 23418
rect 27901 23366 27953 23418
rect 27965 23366 28017 23418
rect 28029 23366 28081 23418
rect 28093 23366 28145 23418
rect 4252 23264 4304 23316
rect 5816 23307 5868 23316
rect 5816 23273 5825 23307
rect 5825 23273 5859 23307
rect 5859 23273 5868 23307
rect 5816 23264 5868 23273
rect 5908 23264 5960 23316
rect 8484 23264 8536 23316
rect 9588 23264 9640 23316
rect 10600 23264 10652 23316
rect 10140 23196 10192 23248
rect 11060 23196 11112 23248
rect 11428 23196 11480 23248
rect 12440 23264 12492 23316
rect 13636 23264 13688 23316
rect 14372 23264 14424 23316
rect 14832 23307 14884 23316
rect 5448 23128 5500 23180
rect 9588 23128 9640 23180
rect 13728 23196 13780 23248
rect 14188 23196 14240 23248
rect 14832 23273 14841 23307
rect 14841 23273 14875 23307
rect 14875 23273 14884 23307
rect 14832 23264 14884 23273
rect 14924 23264 14976 23316
rect 15292 23264 15344 23316
rect 15844 23264 15896 23316
rect 16580 23264 16632 23316
rect 16672 23264 16724 23316
rect 15384 23196 15436 23248
rect 1584 23103 1636 23112
rect 1584 23069 1593 23103
rect 1593 23069 1627 23103
rect 1627 23069 1636 23103
rect 1584 23060 1636 23069
rect 5080 23060 5132 23112
rect 8024 23060 8076 23112
rect 9404 23060 9456 23112
rect 10508 23060 10560 23112
rect 6552 22992 6604 23044
rect 6644 22992 6696 23044
rect 12992 23128 13044 23180
rect 11244 23060 11296 23112
rect 11428 23060 11480 23112
rect 11612 23060 11664 23112
rect 12164 23060 12216 23112
rect 12808 23103 12860 23112
rect 12808 23069 12817 23103
rect 12817 23069 12851 23103
rect 12851 23069 12860 23103
rect 12808 23060 12860 23069
rect 13452 23060 13504 23112
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 13912 23060 13964 23112
rect 14372 23060 14424 23112
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 14832 23128 14884 23180
rect 16120 23128 16172 23180
rect 15660 23103 15712 23112
rect 15292 23035 15344 23044
rect 15292 23001 15301 23035
rect 15301 23001 15335 23035
rect 15335 23001 15344 23035
rect 15292 22992 15344 23001
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 15844 23060 15896 23112
rect 16212 23103 16264 23112
rect 16212 23069 16221 23103
rect 16221 23069 16255 23103
rect 16255 23069 16264 23103
rect 16212 23060 16264 23069
rect 16396 23060 16448 23112
rect 17132 23128 17184 23180
rect 17868 23128 17920 23180
rect 18420 23196 18472 23248
rect 19984 23264 20036 23316
rect 15936 22992 15988 23044
rect 16120 22992 16172 23044
rect 16856 23060 16908 23112
rect 16948 23060 17000 23112
rect 17316 23103 17368 23112
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17500 23103 17552 23112
rect 17316 23060 17368 23069
rect 17500 23069 17509 23103
rect 17509 23069 17543 23103
rect 17543 23069 17552 23103
rect 17500 23060 17552 23069
rect 17684 23060 17736 23112
rect 19340 23128 19392 23180
rect 19524 23196 19576 23248
rect 20812 23196 20864 23248
rect 21272 23264 21324 23316
rect 24860 23264 24912 23316
rect 22560 23196 22612 23248
rect 24032 23196 24084 23248
rect 26792 23264 26844 23316
rect 27712 23264 27764 23316
rect 28540 23264 28592 23316
rect 28816 23307 28868 23316
rect 28816 23273 28825 23307
rect 28825 23273 28859 23307
rect 28859 23273 28868 23307
rect 28816 23264 28868 23273
rect 29736 23264 29788 23316
rect 30104 23264 30156 23316
rect 30196 23264 30248 23316
rect 26976 23239 27028 23248
rect 26976 23205 26985 23239
rect 26985 23205 27019 23239
rect 27019 23205 27028 23239
rect 26976 23196 27028 23205
rect 27804 23196 27856 23248
rect 17132 22992 17184 23044
rect 17868 22992 17920 23044
rect 19524 23060 19576 23112
rect 19800 23060 19852 23112
rect 20352 23128 20404 23180
rect 21456 23128 21508 23180
rect 22100 23128 22152 23180
rect 19064 22992 19116 23044
rect 19156 22992 19208 23044
rect 6092 22924 6144 22976
rect 7472 22924 7524 22976
rect 7656 22924 7708 22976
rect 9036 22924 9088 22976
rect 10876 22967 10928 22976
rect 10876 22933 10885 22967
rect 10885 22933 10919 22967
rect 10919 22933 10928 22967
rect 10876 22924 10928 22933
rect 11704 22924 11756 22976
rect 12072 22967 12124 22976
rect 12072 22933 12081 22967
rect 12081 22933 12115 22967
rect 12115 22933 12124 22967
rect 12072 22924 12124 22933
rect 12164 22924 12216 22976
rect 13268 22924 13320 22976
rect 14096 22924 14148 22976
rect 16672 22924 16724 22976
rect 16764 22924 16816 22976
rect 20444 23060 20496 23112
rect 21272 23103 21324 23112
rect 21272 23069 21281 23103
rect 21281 23069 21315 23103
rect 21315 23069 21324 23103
rect 21272 23060 21324 23069
rect 21364 23060 21416 23112
rect 21640 23060 21692 23112
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 22192 23060 22244 23112
rect 23112 23128 23164 23180
rect 23664 23128 23716 23180
rect 24124 23060 24176 23112
rect 25044 23128 25096 23180
rect 26332 23103 26384 23112
rect 26332 23069 26341 23103
rect 26341 23069 26375 23103
rect 26375 23069 26384 23103
rect 26332 23060 26384 23069
rect 26700 23060 26752 23112
rect 27068 23103 27120 23112
rect 27068 23069 27077 23103
rect 27077 23069 27111 23103
rect 27111 23069 27120 23103
rect 27068 23060 27120 23069
rect 27620 23103 27672 23112
rect 27620 23069 27629 23103
rect 27629 23069 27663 23103
rect 27663 23069 27672 23103
rect 27620 23060 27672 23069
rect 27712 23060 27764 23112
rect 28816 23060 28868 23112
rect 29276 23128 29328 23180
rect 29736 23171 29788 23180
rect 29736 23137 29745 23171
rect 29745 23137 29779 23171
rect 29779 23137 29788 23171
rect 29736 23128 29788 23137
rect 29552 23060 29604 23112
rect 29644 23060 29696 23112
rect 31116 23196 31168 23248
rect 30288 23128 30340 23180
rect 31024 23128 31076 23180
rect 21456 22992 21508 23044
rect 22100 22992 22152 23044
rect 24676 22992 24728 23044
rect 26056 23035 26108 23044
rect 26056 23001 26065 23035
rect 26065 23001 26099 23035
rect 26099 23001 26108 23035
rect 26056 22992 26108 23001
rect 20628 22924 20680 22976
rect 21088 22924 21140 22976
rect 24032 22924 24084 22976
rect 25412 22924 25464 22976
rect 25688 22924 25740 22976
rect 30288 22992 30340 23044
rect 30932 23060 30984 23112
rect 32772 23060 32824 23112
rect 31024 22992 31076 23044
rect 26424 22924 26476 22976
rect 27068 22924 27120 22976
rect 27252 22924 27304 22976
rect 30748 22924 30800 22976
rect 31484 22924 31536 22976
rect 8632 22822 8684 22874
rect 8696 22822 8748 22874
rect 8760 22822 8812 22874
rect 8824 22822 8876 22874
rect 8888 22822 8940 22874
rect 16314 22822 16366 22874
rect 16378 22822 16430 22874
rect 16442 22822 16494 22874
rect 16506 22822 16558 22874
rect 16570 22822 16622 22874
rect 23996 22822 24048 22874
rect 24060 22822 24112 22874
rect 24124 22822 24176 22874
rect 24188 22822 24240 22874
rect 24252 22822 24304 22874
rect 31678 22822 31730 22874
rect 31742 22822 31794 22874
rect 31806 22822 31858 22874
rect 31870 22822 31922 22874
rect 31934 22822 31986 22874
rect 5632 22720 5684 22772
rect 7104 22763 7156 22772
rect 7104 22729 7113 22763
rect 7113 22729 7147 22763
rect 7147 22729 7156 22763
rect 7104 22720 7156 22729
rect 8208 22763 8260 22772
rect 8208 22729 8217 22763
rect 8217 22729 8251 22763
rect 8251 22729 8260 22763
rect 8208 22720 8260 22729
rect 11980 22720 12032 22772
rect 12348 22720 12400 22772
rect 12716 22720 12768 22772
rect 12900 22720 12952 22772
rect 13544 22720 13596 22772
rect 4436 22652 4488 22704
rect 5172 22652 5224 22704
rect 8116 22652 8168 22704
rect 10416 22695 10468 22704
rect 10416 22661 10425 22695
rect 10425 22661 10459 22695
rect 10459 22661 10468 22695
rect 10416 22652 10468 22661
rect 11428 22652 11480 22704
rect 14096 22720 14148 22772
rect 16028 22720 16080 22772
rect 16120 22720 16172 22772
rect 16580 22720 16632 22772
rect 19708 22720 19760 22772
rect 19800 22720 19852 22772
rect 21180 22720 21232 22772
rect 21272 22720 21324 22772
rect 22008 22720 22060 22772
rect 22744 22720 22796 22772
rect 10324 22627 10376 22636
rect 10324 22593 10333 22627
rect 10333 22593 10367 22627
rect 10367 22593 10376 22627
rect 10324 22584 10376 22593
rect 10508 22627 10560 22636
rect 10508 22593 10517 22627
rect 10517 22593 10551 22627
rect 10551 22593 10560 22627
rect 10508 22584 10560 22593
rect 5908 22516 5960 22568
rect 5816 22448 5868 22500
rect 6368 22448 6420 22500
rect 9312 22448 9364 22500
rect 6092 22380 6144 22432
rect 8760 22423 8812 22432
rect 8760 22389 8769 22423
rect 8769 22389 8803 22423
rect 8803 22389 8812 22423
rect 8760 22380 8812 22389
rect 9864 22491 9916 22500
rect 9864 22457 9873 22491
rect 9873 22457 9907 22491
rect 9907 22457 9916 22491
rect 9864 22448 9916 22457
rect 11612 22584 11664 22636
rect 12440 22516 12492 22568
rect 12808 22584 12860 22636
rect 12900 22584 12952 22636
rect 13084 22584 13136 22636
rect 13360 22627 13412 22636
rect 13360 22593 13411 22627
rect 13411 22593 13412 22627
rect 13360 22584 13412 22593
rect 13820 22584 13872 22636
rect 14648 22652 14700 22704
rect 15016 22652 15068 22704
rect 15476 22652 15528 22704
rect 15844 22652 15896 22704
rect 16856 22652 16908 22704
rect 17408 22652 17460 22704
rect 17868 22652 17920 22704
rect 18144 22652 18196 22704
rect 20352 22695 20404 22704
rect 20352 22661 20361 22695
rect 20361 22661 20395 22695
rect 20395 22661 20404 22695
rect 20352 22652 20404 22661
rect 21548 22652 21600 22704
rect 15108 22627 15160 22636
rect 15108 22593 15117 22627
rect 15117 22593 15151 22627
rect 15151 22593 15160 22627
rect 15108 22584 15160 22593
rect 13912 22516 13964 22568
rect 10784 22380 10836 22432
rect 11060 22380 11112 22432
rect 13268 22448 13320 22500
rect 14096 22516 14148 22568
rect 16304 22584 16356 22636
rect 16764 22584 16816 22636
rect 17592 22584 17644 22636
rect 18236 22584 18288 22636
rect 18696 22627 18748 22636
rect 15568 22516 15620 22568
rect 16028 22516 16080 22568
rect 15016 22448 15068 22500
rect 16212 22448 16264 22500
rect 16488 22448 16540 22500
rect 16764 22448 16816 22500
rect 16948 22448 17000 22500
rect 17040 22448 17092 22500
rect 17316 22448 17368 22500
rect 12348 22380 12400 22432
rect 12716 22380 12768 22432
rect 17408 22380 17460 22432
rect 17776 22516 17828 22568
rect 18696 22593 18705 22627
rect 18705 22593 18739 22627
rect 18739 22593 18748 22627
rect 18696 22584 18748 22593
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 18972 22584 19024 22636
rect 19248 22559 19300 22568
rect 19248 22525 19257 22559
rect 19257 22525 19291 22559
rect 19291 22525 19300 22559
rect 19248 22516 19300 22525
rect 19524 22559 19576 22568
rect 19524 22525 19533 22559
rect 19533 22525 19567 22559
rect 19567 22525 19576 22559
rect 19524 22516 19576 22525
rect 19984 22584 20036 22636
rect 20720 22584 20772 22636
rect 21916 22584 21968 22636
rect 22652 22584 22704 22636
rect 17960 22448 18012 22500
rect 18512 22448 18564 22500
rect 19340 22448 19392 22500
rect 19984 22448 20036 22500
rect 19524 22380 19576 22432
rect 20076 22380 20128 22432
rect 21548 22516 21600 22568
rect 21640 22516 21692 22568
rect 22376 22516 22428 22568
rect 22744 22516 22796 22568
rect 22928 22559 22980 22568
rect 22928 22525 22937 22559
rect 22937 22525 22971 22559
rect 22971 22525 22980 22559
rect 22928 22516 22980 22525
rect 25320 22652 25372 22704
rect 25964 22652 26016 22704
rect 29644 22652 29696 22704
rect 23756 22627 23808 22636
rect 23756 22593 23765 22627
rect 23765 22593 23799 22627
rect 23799 22593 23808 22627
rect 23756 22584 23808 22593
rect 24584 22584 24636 22636
rect 26332 22627 26384 22636
rect 26332 22593 26341 22627
rect 26341 22593 26375 22627
rect 26375 22593 26384 22627
rect 26332 22584 26384 22593
rect 26516 22584 26568 22636
rect 26976 22584 27028 22636
rect 27252 22627 27304 22636
rect 25964 22516 26016 22568
rect 21088 22448 21140 22500
rect 21180 22380 21232 22432
rect 21824 22448 21876 22500
rect 23664 22448 23716 22500
rect 24860 22448 24912 22500
rect 26424 22516 26476 22568
rect 27252 22593 27271 22627
rect 27271 22593 27304 22627
rect 27252 22584 27304 22593
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 28264 22584 28316 22636
rect 28080 22516 28132 22568
rect 28448 22584 28500 22636
rect 29184 22584 29236 22636
rect 29552 22627 29604 22636
rect 29552 22593 29561 22627
rect 29561 22593 29595 22627
rect 29595 22593 29604 22627
rect 29552 22584 29604 22593
rect 30288 22720 30340 22772
rect 31024 22763 31076 22772
rect 31024 22729 31033 22763
rect 31033 22729 31067 22763
rect 31067 22729 31076 22763
rect 31024 22720 31076 22729
rect 31116 22695 31168 22704
rect 31116 22661 31125 22695
rect 31125 22661 31159 22695
rect 31159 22661 31168 22695
rect 31116 22652 31168 22661
rect 30380 22584 30432 22636
rect 30932 22584 30984 22636
rect 32864 22584 32916 22636
rect 29828 22559 29880 22568
rect 29828 22525 29837 22559
rect 29837 22525 29871 22559
rect 29871 22525 29880 22559
rect 30748 22559 30800 22568
rect 29828 22516 29880 22525
rect 30748 22525 30757 22559
rect 30757 22525 30791 22559
rect 30791 22525 30800 22559
rect 30748 22516 30800 22525
rect 30840 22516 30892 22568
rect 32680 22516 32732 22568
rect 28724 22491 28776 22500
rect 22192 22380 22244 22432
rect 22468 22380 22520 22432
rect 23112 22380 23164 22432
rect 23940 22380 23992 22432
rect 26424 22380 26476 22432
rect 28724 22457 28733 22491
rect 28733 22457 28767 22491
rect 28767 22457 28776 22491
rect 28724 22448 28776 22457
rect 29276 22448 29328 22500
rect 29644 22448 29696 22500
rect 26700 22380 26752 22432
rect 27252 22380 27304 22432
rect 27528 22423 27580 22432
rect 27528 22389 27537 22423
rect 27537 22389 27571 22423
rect 27571 22389 27580 22423
rect 27528 22380 27580 22389
rect 28632 22380 28684 22432
rect 29000 22380 29052 22432
rect 30104 22380 30156 22432
rect 30288 22423 30340 22432
rect 30288 22389 30297 22423
rect 30297 22389 30331 22423
rect 30331 22389 30340 22423
rect 30288 22380 30340 22389
rect 30748 22380 30800 22432
rect 32128 22380 32180 22432
rect 4791 22278 4843 22330
rect 4855 22278 4907 22330
rect 4919 22278 4971 22330
rect 4983 22278 5035 22330
rect 5047 22278 5099 22330
rect 12473 22278 12525 22330
rect 12537 22278 12589 22330
rect 12601 22278 12653 22330
rect 12665 22278 12717 22330
rect 12729 22278 12781 22330
rect 20155 22278 20207 22330
rect 20219 22278 20271 22330
rect 20283 22278 20335 22330
rect 20347 22278 20399 22330
rect 20411 22278 20463 22330
rect 27837 22278 27889 22330
rect 27901 22278 27953 22330
rect 27965 22278 28017 22330
rect 28029 22278 28081 22330
rect 28093 22278 28145 22330
rect 5540 22176 5592 22228
rect 5908 22176 5960 22228
rect 6368 22219 6420 22228
rect 6368 22185 6377 22219
rect 6377 22185 6411 22219
rect 6411 22185 6420 22219
rect 6368 22176 6420 22185
rect 6552 22176 6604 22228
rect 9588 22176 9640 22228
rect 9772 22176 9824 22228
rect 11152 22176 11204 22228
rect 11980 22219 12032 22228
rect 11980 22185 11989 22219
rect 11989 22185 12023 22219
rect 12023 22185 12032 22219
rect 11980 22176 12032 22185
rect 11060 22151 11112 22160
rect 5356 22040 5408 22092
rect 9312 22040 9364 22092
rect 10784 22040 10836 22092
rect 11060 22117 11069 22151
rect 11069 22117 11103 22151
rect 11103 22117 11112 22151
rect 14096 22176 14148 22228
rect 14280 22219 14332 22228
rect 14280 22185 14289 22219
rect 14289 22185 14323 22219
rect 14323 22185 14332 22219
rect 14280 22176 14332 22185
rect 14464 22219 14516 22228
rect 14464 22185 14473 22219
rect 14473 22185 14507 22219
rect 14507 22185 14516 22219
rect 14464 22176 14516 22185
rect 11060 22108 11112 22117
rect 13084 22108 13136 22160
rect 17132 22176 17184 22228
rect 4712 22015 4764 22024
rect 4712 21981 4721 22015
rect 4721 21981 4755 22015
rect 4755 21981 4764 22015
rect 4712 21972 4764 21981
rect 9588 22015 9640 22024
rect 4252 21904 4304 21956
rect 9128 21904 9180 21956
rect 6552 21836 6604 21888
rect 7564 21836 7616 21888
rect 8484 21879 8536 21888
rect 8484 21845 8493 21879
rect 8493 21845 8527 21879
rect 8527 21845 8536 21879
rect 8484 21836 8536 21845
rect 9588 21981 9597 22015
rect 9597 21981 9631 22015
rect 9631 21981 9640 22015
rect 9588 21972 9640 21981
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10324 22015 10376 22024
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 10324 21972 10376 21981
rect 9956 21904 10008 21956
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 12348 22040 12400 22092
rect 11336 21904 11388 21956
rect 11428 21904 11480 21956
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 13636 22040 13688 22092
rect 13084 21972 13136 22024
rect 13452 22015 13504 22024
rect 13452 21981 13461 22015
rect 13461 21981 13495 22015
rect 13495 21981 13504 22015
rect 13452 21972 13504 21981
rect 16580 22108 16632 22160
rect 19156 22176 19208 22228
rect 17408 22108 17460 22160
rect 18052 22108 18104 22160
rect 18328 22108 18380 22160
rect 18420 22108 18472 22160
rect 20720 22176 20772 22228
rect 20996 22176 21048 22228
rect 23664 22176 23716 22228
rect 24676 22176 24728 22228
rect 25136 22176 25188 22228
rect 25780 22176 25832 22228
rect 26148 22176 26200 22228
rect 26700 22176 26752 22228
rect 26976 22176 27028 22228
rect 28448 22176 28500 22228
rect 28632 22176 28684 22228
rect 29092 22219 29144 22228
rect 15660 22083 15712 22092
rect 15660 22049 15669 22083
rect 15669 22049 15703 22083
rect 15703 22049 15712 22083
rect 15660 22040 15712 22049
rect 16120 22040 16172 22092
rect 16948 22040 17000 22092
rect 15936 21972 15988 22024
rect 12256 21904 12308 21956
rect 14556 21904 14608 21956
rect 15200 21904 15252 21956
rect 15384 21904 15436 21956
rect 16028 21904 16080 21956
rect 16488 21904 16540 21956
rect 17316 22040 17368 22092
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 17776 22015 17828 22024
rect 17776 21981 17785 22015
rect 17785 21981 17819 22015
rect 17819 21981 17828 22015
rect 17776 21972 17828 21981
rect 18052 21972 18104 22024
rect 18144 21972 18196 22024
rect 18328 21972 18380 22024
rect 19524 22108 19576 22160
rect 21916 22151 21968 22160
rect 18880 22083 18932 22092
rect 18880 22049 18889 22083
rect 18889 22049 18923 22083
rect 18923 22049 18932 22083
rect 18880 22040 18932 22049
rect 19248 22040 19300 22092
rect 21916 22117 21925 22151
rect 21925 22117 21959 22151
rect 21959 22117 21968 22151
rect 21916 22108 21968 22117
rect 26424 22108 26476 22160
rect 20996 22040 21048 22092
rect 21456 22040 21508 22092
rect 25596 22040 25648 22092
rect 26148 22083 26200 22092
rect 26148 22049 26157 22083
rect 26157 22049 26191 22083
rect 26191 22049 26200 22083
rect 26148 22040 26200 22049
rect 19708 21972 19760 22024
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 23664 22015 23716 22024
rect 23664 21981 23666 22015
rect 23666 21981 23700 22015
rect 23700 21981 23716 22015
rect 23664 21972 23716 21981
rect 26608 22108 26660 22160
rect 29092 22185 29101 22219
rect 29101 22185 29135 22219
rect 29135 22185 29144 22219
rect 29092 22176 29144 22185
rect 29276 22176 29328 22228
rect 26700 22040 26752 22092
rect 12900 21836 12952 21888
rect 13268 21879 13320 21888
rect 13268 21845 13277 21879
rect 13277 21845 13311 21879
rect 13311 21845 13320 21879
rect 13268 21836 13320 21845
rect 13636 21879 13688 21888
rect 13636 21845 13645 21879
rect 13645 21845 13679 21879
rect 13679 21845 13688 21879
rect 13636 21836 13688 21845
rect 14188 21836 14240 21888
rect 17316 21836 17368 21888
rect 17960 21904 18012 21956
rect 18788 21904 18840 21956
rect 18880 21904 18932 21956
rect 19524 21904 19576 21956
rect 21180 21904 21232 21956
rect 22376 21904 22428 21956
rect 23296 21904 23348 21956
rect 24492 21904 24544 21956
rect 24768 21904 24820 21956
rect 25872 21904 25924 21956
rect 22100 21836 22152 21888
rect 23020 21836 23072 21888
rect 24584 21836 24636 21888
rect 27528 22040 27580 22092
rect 28540 22040 28592 22092
rect 28632 22040 28684 22092
rect 27252 22015 27304 22024
rect 27252 21981 27261 22015
rect 27261 21981 27295 22015
rect 27295 21981 27304 22015
rect 27252 21972 27304 21981
rect 27988 22015 28040 22018
rect 27988 21981 27997 22015
rect 27997 21981 28031 22015
rect 28031 21981 28040 22015
rect 30288 22108 30340 22160
rect 27988 21966 28040 21981
rect 27344 21904 27396 21956
rect 27160 21836 27212 21888
rect 27436 21836 27488 21888
rect 28172 21904 28224 21956
rect 28908 21972 28960 22024
rect 29000 22015 29052 22024
rect 29000 21981 29009 22015
rect 29009 21981 29043 22015
rect 29043 21981 29052 22015
rect 29000 21972 29052 21981
rect 28908 21836 28960 21888
rect 29092 21904 29144 21956
rect 30564 22040 30616 22092
rect 29276 21972 29328 22024
rect 29552 21972 29604 22024
rect 29644 21972 29696 22024
rect 30104 22015 30156 22024
rect 30104 21981 30113 22015
rect 30113 21981 30147 22015
rect 30147 21981 30156 22015
rect 30104 21972 30156 21981
rect 29828 21947 29880 21956
rect 29828 21913 29837 21947
rect 29837 21913 29871 21947
rect 29871 21913 29880 21947
rect 29828 21904 29880 21913
rect 30104 21836 30156 21888
rect 30380 21972 30432 22024
rect 31024 22015 31076 22024
rect 31024 21981 31033 22015
rect 31033 21981 31067 22015
rect 31067 21981 31076 22015
rect 31024 21972 31076 21981
rect 31484 21972 31536 22024
rect 30288 21836 30340 21888
rect 31116 21879 31168 21888
rect 31116 21845 31125 21879
rect 31125 21845 31159 21879
rect 31159 21845 31168 21879
rect 31116 21836 31168 21845
rect 8632 21734 8684 21786
rect 8696 21734 8748 21786
rect 8760 21734 8812 21786
rect 8824 21734 8876 21786
rect 8888 21734 8940 21786
rect 16314 21734 16366 21786
rect 16378 21734 16430 21786
rect 16442 21734 16494 21786
rect 16506 21734 16558 21786
rect 16570 21734 16622 21786
rect 23996 21734 24048 21786
rect 24060 21734 24112 21786
rect 24124 21734 24176 21786
rect 24188 21734 24240 21786
rect 24252 21734 24304 21786
rect 31678 21734 31730 21786
rect 31742 21734 31794 21786
rect 31806 21734 31858 21786
rect 31870 21734 31922 21786
rect 31934 21734 31986 21786
rect 5448 21675 5500 21684
rect 5448 21641 5457 21675
rect 5457 21641 5491 21675
rect 5491 21641 5500 21675
rect 5448 21632 5500 21641
rect 5816 21632 5868 21684
rect 9864 21632 9916 21684
rect 11244 21632 11296 21684
rect 11336 21632 11388 21684
rect 11980 21632 12032 21684
rect 13268 21632 13320 21684
rect 13452 21632 13504 21684
rect 5540 21564 5592 21616
rect 7564 21564 7616 21616
rect 11428 21564 11480 21616
rect 11796 21564 11848 21616
rect 9772 21539 9824 21548
rect 9772 21505 9781 21539
rect 9781 21505 9815 21539
rect 9815 21505 9824 21539
rect 9772 21496 9824 21505
rect 10600 21496 10652 21548
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 9680 21471 9732 21480
rect 9680 21437 9689 21471
rect 9689 21437 9723 21471
rect 9723 21437 9732 21471
rect 9680 21428 9732 21437
rect 9864 21428 9916 21480
rect 12716 21496 12768 21548
rect 12992 21607 13044 21616
rect 12992 21573 13001 21607
rect 13001 21573 13035 21607
rect 13035 21573 13044 21607
rect 12992 21564 13044 21573
rect 14004 21564 14056 21616
rect 14924 21632 14976 21684
rect 16028 21632 16080 21684
rect 16120 21632 16172 21684
rect 16580 21632 16632 21684
rect 16844 21632 16896 21684
rect 17040 21632 17092 21684
rect 17316 21632 17368 21684
rect 17408 21632 17460 21684
rect 18144 21632 18196 21684
rect 18236 21632 18288 21684
rect 9312 21360 9364 21412
rect 10968 21360 11020 21412
rect 12256 21360 12308 21412
rect 12532 21403 12584 21412
rect 12532 21369 12541 21403
rect 12541 21369 12575 21403
rect 12575 21369 12584 21403
rect 12532 21360 12584 21369
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 7932 21292 7984 21344
rect 8944 21292 8996 21344
rect 9220 21292 9272 21344
rect 10508 21292 10560 21344
rect 12992 21292 13044 21344
rect 13360 21335 13412 21344
rect 13360 21301 13369 21335
rect 13369 21301 13403 21335
rect 13403 21301 13412 21335
rect 13360 21292 13412 21301
rect 13912 21471 13964 21480
rect 13912 21437 13921 21471
rect 13921 21437 13955 21471
rect 13955 21437 13964 21471
rect 13912 21428 13964 21437
rect 15292 21496 15344 21548
rect 14648 21428 14700 21480
rect 16304 21564 16356 21616
rect 16672 21564 16724 21616
rect 19340 21632 19392 21684
rect 19892 21632 19944 21684
rect 21364 21632 21416 21684
rect 22284 21632 22336 21684
rect 22560 21632 22612 21684
rect 22744 21632 22796 21684
rect 23388 21632 23440 21684
rect 23664 21632 23716 21684
rect 18696 21564 18748 21616
rect 19156 21564 19208 21616
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 16028 21496 16080 21548
rect 17684 21496 17736 21548
rect 18972 21496 19024 21548
rect 19340 21496 19392 21548
rect 19984 21564 20036 21616
rect 20996 21564 21048 21616
rect 23848 21632 23900 21684
rect 29828 21632 29880 21684
rect 30748 21632 30800 21684
rect 22100 21496 22152 21548
rect 26332 21564 26384 21616
rect 26700 21564 26752 21616
rect 26792 21564 26844 21616
rect 26976 21564 27028 21616
rect 27160 21564 27212 21616
rect 28172 21564 28224 21616
rect 28816 21564 28868 21616
rect 24676 21496 24728 21548
rect 26608 21539 26660 21548
rect 26608 21505 26617 21539
rect 26617 21505 26651 21539
rect 26651 21505 26660 21539
rect 26608 21496 26660 21505
rect 17592 21428 17644 21480
rect 18236 21428 18288 21480
rect 18420 21471 18472 21480
rect 18420 21437 18429 21471
rect 18429 21437 18463 21471
rect 18463 21437 18472 21471
rect 18420 21428 18472 21437
rect 18512 21428 18564 21480
rect 18696 21428 18748 21480
rect 18788 21428 18840 21480
rect 19800 21428 19852 21480
rect 26976 21428 27028 21480
rect 28908 21496 28960 21548
rect 29552 21564 29604 21616
rect 29920 21564 29972 21616
rect 30288 21496 30340 21548
rect 30656 21539 30708 21548
rect 15936 21360 15988 21412
rect 17684 21360 17736 21412
rect 17776 21360 17828 21412
rect 18420 21292 18472 21344
rect 19248 21360 19300 21412
rect 19432 21360 19484 21412
rect 20720 21360 20772 21412
rect 20812 21292 20864 21344
rect 20996 21360 21048 21412
rect 21824 21360 21876 21412
rect 22468 21360 22520 21412
rect 24952 21360 25004 21412
rect 30380 21428 30432 21480
rect 23020 21292 23072 21344
rect 23204 21292 23256 21344
rect 28448 21360 28500 21412
rect 29368 21360 29420 21412
rect 30656 21505 30665 21539
rect 30665 21505 30699 21539
rect 30699 21505 30708 21539
rect 30656 21496 30708 21505
rect 30840 21539 30892 21548
rect 30840 21505 30849 21539
rect 30849 21505 30883 21539
rect 30883 21505 30892 21539
rect 30840 21496 30892 21505
rect 30656 21360 30708 21412
rect 26976 21292 27028 21344
rect 28816 21292 28868 21344
rect 28908 21335 28960 21344
rect 28908 21301 28917 21335
rect 28917 21301 28951 21335
rect 28951 21301 28960 21335
rect 28908 21292 28960 21301
rect 29460 21292 29512 21344
rect 31116 21335 31168 21344
rect 31116 21301 31125 21335
rect 31125 21301 31159 21335
rect 31159 21301 31168 21335
rect 31116 21292 31168 21301
rect 4791 21190 4843 21242
rect 4855 21190 4907 21242
rect 4919 21190 4971 21242
rect 4983 21190 5035 21242
rect 5047 21190 5099 21242
rect 12473 21190 12525 21242
rect 12537 21190 12589 21242
rect 12601 21190 12653 21242
rect 12665 21190 12717 21242
rect 12729 21190 12781 21242
rect 20155 21190 20207 21242
rect 20219 21190 20271 21242
rect 20283 21190 20335 21242
rect 20347 21190 20399 21242
rect 20411 21190 20463 21242
rect 27837 21190 27889 21242
rect 27901 21190 27953 21242
rect 27965 21190 28017 21242
rect 28029 21190 28081 21242
rect 28093 21190 28145 21242
rect 7472 21088 7524 21140
rect 7656 21088 7708 21140
rect 8300 21088 8352 21140
rect 9128 21088 9180 21140
rect 11796 21088 11848 21140
rect 12440 21088 12492 21140
rect 13360 21088 13412 21140
rect 15384 21088 15436 21140
rect 16488 21088 16540 21140
rect 17868 21088 17920 21140
rect 18052 21088 18104 21140
rect 10600 21020 10652 21072
rect 8300 20952 8352 21004
rect 9312 20952 9364 21004
rect 9956 20884 10008 20936
rect 10232 20884 10284 20936
rect 10508 20927 10560 20936
rect 8300 20816 8352 20868
rect 8944 20816 8996 20868
rect 6000 20748 6052 20800
rect 7380 20791 7432 20800
rect 7380 20757 7389 20791
rect 7389 20757 7423 20791
rect 7423 20757 7432 20791
rect 7380 20748 7432 20757
rect 8024 20791 8076 20800
rect 8024 20757 8033 20791
rect 8033 20757 8067 20791
rect 8067 20757 8076 20791
rect 8024 20748 8076 20757
rect 8116 20748 8168 20800
rect 8392 20748 8444 20800
rect 9036 20748 9088 20800
rect 9496 20816 9548 20868
rect 10508 20893 10517 20927
rect 10517 20893 10551 20927
rect 10551 20893 10560 20927
rect 10508 20884 10560 20893
rect 10876 20884 10928 20936
rect 11428 20952 11480 21004
rect 11980 20952 12032 21004
rect 11152 20816 11204 20868
rect 11796 20884 11848 20936
rect 12072 20927 12124 20936
rect 12072 20893 12081 20927
rect 12081 20893 12115 20927
rect 12115 20893 12124 20927
rect 12072 20884 12124 20893
rect 12532 20927 12584 20936
rect 12532 20893 12541 20927
rect 12541 20893 12575 20927
rect 12575 20893 12584 20927
rect 12532 20884 12584 20893
rect 13176 20952 13228 21004
rect 13452 20952 13504 21004
rect 15016 21020 15068 21072
rect 14464 20952 14516 21004
rect 16120 21020 16172 21072
rect 16304 21020 16356 21072
rect 16856 21020 16908 21072
rect 16396 20995 16448 21004
rect 16396 20961 16405 20995
rect 16405 20961 16439 20995
rect 16439 20961 16448 20995
rect 16396 20952 16448 20961
rect 16488 20952 16540 21004
rect 17776 21020 17828 21072
rect 18696 21088 18748 21140
rect 19984 21088 20036 21140
rect 18788 21020 18840 21072
rect 21456 21088 21508 21140
rect 25504 21088 25556 21140
rect 25596 21088 25648 21140
rect 29000 21088 29052 21140
rect 29368 21088 29420 21140
rect 31300 21131 31352 21140
rect 31300 21097 31309 21131
rect 31309 21097 31343 21131
rect 31343 21097 31352 21131
rect 31300 21088 31352 21097
rect 29736 21063 29788 21072
rect 9588 20748 9640 20800
rect 9772 20791 9824 20800
rect 9772 20757 9781 20791
rect 9781 20757 9815 20791
rect 9815 20757 9824 20791
rect 9772 20748 9824 20757
rect 10416 20791 10468 20800
rect 10416 20757 10425 20791
rect 10425 20757 10459 20791
rect 10459 20757 10468 20791
rect 10416 20748 10468 20757
rect 11060 20748 11112 20800
rect 11244 20791 11296 20800
rect 11244 20757 11253 20791
rect 11253 20757 11287 20791
rect 11287 20757 11296 20791
rect 11244 20748 11296 20757
rect 11796 20748 11848 20800
rect 12624 20748 12676 20800
rect 13084 20748 13136 20800
rect 13636 20748 13688 20800
rect 15200 20816 15252 20868
rect 15752 20884 15804 20936
rect 16580 20884 16632 20936
rect 17592 20952 17644 21004
rect 18236 20927 18288 20936
rect 15844 20816 15896 20868
rect 16028 20816 16080 20868
rect 16764 20816 16816 20868
rect 14464 20791 14516 20800
rect 14464 20757 14491 20791
rect 14491 20757 14516 20791
rect 14464 20748 14516 20757
rect 14740 20748 14792 20800
rect 15476 20748 15528 20800
rect 15660 20791 15712 20800
rect 15660 20757 15669 20791
rect 15669 20757 15703 20791
rect 15703 20757 15712 20791
rect 15660 20748 15712 20757
rect 15936 20748 15988 20800
rect 17224 20748 17276 20800
rect 17684 20816 17736 20868
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 18328 20884 18380 20936
rect 20720 20952 20772 21004
rect 20812 20952 20864 21004
rect 21548 20952 21600 21004
rect 29736 21029 29745 21063
rect 29745 21029 29779 21063
rect 29779 21029 29788 21063
rect 29736 21020 29788 21029
rect 30012 21020 30064 21072
rect 27344 20952 27396 21004
rect 27620 20952 27672 21004
rect 18604 20927 18656 20936
rect 18604 20893 18613 20927
rect 18613 20893 18647 20927
rect 18647 20893 18656 20927
rect 18604 20884 18656 20893
rect 18788 20884 18840 20936
rect 19800 20884 19852 20936
rect 19892 20884 19944 20936
rect 18144 20816 18196 20868
rect 18328 20748 18380 20800
rect 20076 20748 20128 20800
rect 20536 20816 20588 20868
rect 20996 20816 21048 20868
rect 20628 20748 20680 20800
rect 20904 20748 20956 20800
rect 26700 20884 26752 20936
rect 25228 20816 25280 20868
rect 26240 20859 26292 20868
rect 26240 20825 26249 20859
rect 26249 20825 26283 20859
rect 26283 20825 26292 20859
rect 26240 20816 26292 20825
rect 26608 20816 26660 20868
rect 28540 20952 28592 21004
rect 29828 20952 29880 21004
rect 30196 20952 30248 21004
rect 27252 20859 27304 20868
rect 27252 20825 27261 20859
rect 27261 20825 27295 20859
rect 27295 20825 27304 20859
rect 27252 20816 27304 20825
rect 28540 20816 28592 20868
rect 29644 20816 29696 20868
rect 30288 20884 30340 20936
rect 31300 20884 31352 20936
rect 30840 20859 30892 20868
rect 30840 20825 30849 20859
rect 30849 20825 30883 20859
rect 30883 20825 30892 20859
rect 30840 20816 30892 20825
rect 25964 20748 26016 20800
rect 26056 20748 26108 20800
rect 28632 20748 28684 20800
rect 29368 20748 29420 20800
rect 29736 20748 29788 20800
rect 30196 20748 30248 20800
rect 8632 20646 8684 20698
rect 8696 20646 8748 20698
rect 8760 20646 8812 20698
rect 8824 20646 8876 20698
rect 8888 20646 8940 20698
rect 16314 20646 16366 20698
rect 16378 20646 16430 20698
rect 16442 20646 16494 20698
rect 16506 20646 16558 20698
rect 16570 20646 16622 20698
rect 23996 20646 24048 20698
rect 24060 20646 24112 20698
rect 24124 20646 24176 20698
rect 24188 20646 24240 20698
rect 24252 20646 24304 20698
rect 31678 20646 31730 20698
rect 31742 20646 31794 20698
rect 31806 20646 31858 20698
rect 31870 20646 31922 20698
rect 31934 20646 31986 20698
rect 8300 20544 8352 20596
rect 9864 20544 9916 20596
rect 12900 20544 12952 20596
rect 9680 20476 9732 20528
rect 14004 20544 14056 20596
rect 16948 20544 17000 20596
rect 17960 20544 18012 20596
rect 22376 20544 22428 20596
rect 9956 20408 10008 20460
rect 10232 20451 10284 20460
rect 10232 20417 10241 20451
rect 10241 20417 10275 20451
rect 10275 20417 10284 20451
rect 10232 20408 10284 20417
rect 10600 20408 10652 20460
rect 10876 20451 10928 20460
rect 10876 20417 10885 20451
rect 10885 20417 10919 20451
rect 10919 20417 10928 20451
rect 10876 20408 10928 20417
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 7380 20340 7432 20392
rect 11336 20408 11388 20460
rect 11796 20408 11848 20460
rect 13084 20519 13136 20528
rect 13084 20485 13093 20519
rect 13093 20485 13127 20519
rect 13127 20485 13136 20519
rect 13084 20476 13136 20485
rect 13452 20476 13504 20528
rect 13544 20476 13596 20528
rect 14096 20408 14148 20460
rect 14280 20408 14332 20460
rect 15660 20408 15712 20460
rect 7472 20272 7524 20324
rect 9680 20315 9732 20324
rect 9680 20281 9689 20315
rect 9689 20281 9723 20315
rect 9723 20281 9732 20315
rect 9680 20272 9732 20281
rect 7656 20204 7708 20256
rect 7932 20204 7984 20256
rect 9036 20247 9088 20256
rect 9036 20213 9045 20247
rect 9045 20213 9079 20247
rect 9079 20213 9088 20247
rect 9036 20204 9088 20213
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 12164 20340 12216 20392
rect 13544 20340 13596 20392
rect 13728 20340 13780 20392
rect 14740 20340 14792 20392
rect 15292 20383 15344 20392
rect 12716 20272 12768 20324
rect 12808 20272 12860 20324
rect 14648 20272 14700 20324
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 15476 20340 15528 20392
rect 15936 20340 15988 20392
rect 16764 20340 16816 20392
rect 17224 20476 17276 20528
rect 18328 20476 18380 20528
rect 17132 20408 17184 20460
rect 17408 20408 17460 20460
rect 16212 20272 16264 20324
rect 17408 20272 17460 20324
rect 12072 20204 12124 20256
rect 12532 20204 12584 20256
rect 12900 20204 12952 20256
rect 13912 20204 13964 20256
rect 14096 20247 14148 20256
rect 14096 20213 14105 20247
rect 14105 20213 14139 20247
rect 14139 20213 14148 20247
rect 14096 20204 14148 20213
rect 14464 20204 14516 20256
rect 14832 20204 14884 20256
rect 15016 20204 15068 20256
rect 16028 20204 16080 20256
rect 16120 20204 16172 20256
rect 17500 20204 17552 20256
rect 17960 20408 18012 20460
rect 18236 20408 18288 20460
rect 18420 20408 18472 20460
rect 19156 20476 19208 20528
rect 19248 20408 19300 20460
rect 19892 20476 19944 20528
rect 20720 20476 20772 20528
rect 21272 20476 21324 20528
rect 25596 20544 25648 20596
rect 26424 20544 26476 20596
rect 29736 20544 29788 20596
rect 25688 20476 25740 20528
rect 26148 20476 26200 20528
rect 27712 20476 27764 20528
rect 29092 20476 29144 20528
rect 29920 20476 29972 20528
rect 30564 20476 30616 20528
rect 18696 20272 18748 20324
rect 18788 20272 18840 20324
rect 18880 20272 18932 20324
rect 21640 20408 21692 20460
rect 21916 20408 21968 20460
rect 20812 20340 20864 20392
rect 19616 20272 19668 20324
rect 17684 20204 17736 20256
rect 17868 20204 17920 20256
rect 18052 20247 18104 20256
rect 18052 20213 18061 20247
rect 18061 20213 18095 20247
rect 18095 20213 18104 20247
rect 18052 20204 18104 20213
rect 18236 20204 18288 20256
rect 19984 20272 20036 20324
rect 21456 20383 21508 20392
rect 21456 20349 21465 20383
rect 21465 20349 21499 20383
rect 21499 20349 21508 20383
rect 21456 20340 21508 20349
rect 22284 20383 22336 20392
rect 21640 20272 21692 20324
rect 19892 20204 19944 20256
rect 21548 20204 21600 20256
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22284 20340 22336 20349
rect 22376 20340 22428 20392
rect 26700 20408 26752 20460
rect 26976 20408 27028 20460
rect 23480 20340 23532 20392
rect 25872 20340 25924 20392
rect 23756 20272 23808 20324
rect 22744 20204 22796 20256
rect 25780 20204 25832 20256
rect 26608 20340 26660 20392
rect 28540 20408 28592 20460
rect 28816 20408 28868 20460
rect 29460 20408 29512 20460
rect 32036 20476 32088 20528
rect 27528 20340 27580 20392
rect 27896 20340 27948 20392
rect 28724 20340 28776 20392
rect 29644 20340 29696 20392
rect 30564 20340 30616 20392
rect 30012 20272 30064 20324
rect 30840 20408 30892 20460
rect 31576 20408 31628 20460
rect 32864 20408 32916 20460
rect 30932 20383 30984 20392
rect 30932 20349 30941 20383
rect 30941 20349 30975 20383
rect 30975 20349 30984 20383
rect 30932 20340 30984 20349
rect 28724 20204 28776 20256
rect 30288 20204 30340 20256
rect 30472 20247 30524 20256
rect 30472 20213 30481 20247
rect 30481 20213 30515 20247
rect 30515 20213 30524 20247
rect 30472 20204 30524 20213
rect 32864 20272 32916 20324
rect 32588 20204 32640 20256
rect 4791 20102 4843 20154
rect 4855 20102 4907 20154
rect 4919 20102 4971 20154
rect 4983 20102 5035 20154
rect 5047 20102 5099 20154
rect 12473 20102 12525 20154
rect 12537 20102 12589 20154
rect 12601 20102 12653 20154
rect 12665 20102 12717 20154
rect 12729 20102 12781 20154
rect 20155 20102 20207 20154
rect 20219 20102 20271 20154
rect 20283 20102 20335 20154
rect 20347 20102 20399 20154
rect 20411 20102 20463 20154
rect 27837 20102 27889 20154
rect 27901 20102 27953 20154
rect 27965 20102 28017 20154
rect 28029 20102 28081 20154
rect 28093 20102 28145 20154
rect 32864 20136 32916 20188
rect 7932 20000 7984 20052
rect 11520 19932 11572 19984
rect 11980 19932 12032 19984
rect 12164 20000 12216 20052
rect 13728 20043 13780 20052
rect 13176 19932 13228 19984
rect 13728 20009 13737 20043
rect 13737 20009 13771 20043
rect 13771 20009 13780 20043
rect 13728 20000 13780 20009
rect 13912 20000 13964 20052
rect 14280 19932 14332 19984
rect 17960 19932 18012 19984
rect 18236 20000 18288 20052
rect 19708 20000 19760 20052
rect 10876 19864 10928 19916
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 7932 19796 7984 19848
rect 10232 19796 10284 19848
rect 8024 19728 8076 19780
rect 9864 19728 9916 19780
rect 10600 19796 10652 19848
rect 11520 19796 11572 19848
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 12348 19864 12400 19916
rect 13636 19864 13688 19916
rect 13820 19864 13872 19916
rect 16212 19907 16264 19916
rect 12256 19796 12308 19848
rect 12624 19796 12676 19848
rect 13268 19796 13320 19848
rect 13452 19796 13504 19848
rect 14280 19796 14332 19848
rect 12716 19771 12768 19780
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 7380 19660 7432 19712
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 11244 19703 11296 19712
rect 11244 19669 11253 19703
rect 11253 19669 11287 19703
rect 11287 19669 11296 19703
rect 11244 19660 11296 19669
rect 12716 19737 12725 19771
rect 12725 19737 12759 19771
rect 12759 19737 12768 19771
rect 12716 19728 12768 19737
rect 12992 19728 13044 19780
rect 14740 19796 14792 19848
rect 14832 19839 14884 19848
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 15016 19796 15068 19848
rect 15476 19839 15528 19848
rect 15476 19805 15485 19839
rect 15485 19805 15519 19839
rect 15519 19805 15528 19839
rect 15476 19796 15528 19805
rect 15568 19796 15620 19848
rect 16212 19873 16221 19907
rect 16221 19873 16255 19907
rect 16255 19873 16264 19907
rect 16212 19864 16264 19873
rect 17224 19864 17276 19916
rect 17132 19796 17184 19848
rect 14648 19771 14700 19780
rect 14648 19737 14657 19771
rect 14657 19737 14691 19771
rect 14691 19737 14700 19771
rect 14648 19728 14700 19737
rect 15108 19728 15160 19780
rect 15660 19728 15712 19780
rect 18696 19932 18748 19984
rect 21640 20000 21692 20052
rect 23020 20000 23072 20052
rect 25044 20000 25096 20052
rect 25320 20000 25372 20052
rect 26516 20000 26568 20052
rect 26792 20000 26844 20052
rect 21916 19932 21968 19984
rect 22468 19932 22520 19984
rect 23480 19932 23532 19984
rect 26148 19932 26200 19984
rect 27712 20000 27764 20052
rect 27436 19975 27488 19984
rect 27436 19941 27445 19975
rect 27445 19941 27479 19975
rect 27479 19941 27488 19975
rect 29000 20000 29052 20052
rect 30840 20000 30892 20052
rect 27436 19932 27488 19941
rect 17684 19796 17736 19848
rect 18144 19796 18196 19848
rect 12532 19660 12584 19712
rect 12808 19703 12860 19712
rect 12808 19669 12817 19703
rect 12817 19669 12851 19703
rect 12851 19669 12860 19703
rect 12808 19660 12860 19669
rect 13636 19660 13688 19712
rect 14188 19660 14240 19712
rect 14280 19660 14332 19712
rect 15936 19660 15988 19712
rect 16028 19660 16080 19712
rect 17408 19660 17460 19712
rect 17960 19728 18012 19780
rect 18972 19796 19024 19848
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 18696 19728 18748 19780
rect 19708 19728 19760 19780
rect 22744 19839 22796 19848
rect 22744 19805 22753 19839
rect 22753 19805 22787 19839
rect 22787 19805 22796 19839
rect 22744 19796 22796 19805
rect 22836 19796 22888 19848
rect 23756 19864 23808 19916
rect 24860 19864 24912 19916
rect 23388 19796 23440 19848
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 26424 19864 26476 19916
rect 26884 19864 26936 19916
rect 27712 19864 27764 19916
rect 26792 19796 26844 19848
rect 19892 19728 19944 19780
rect 20260 19728 20312 19780
rect 22100 19771 22152 19780
rect 18512 19660 18564 19712
rect 19340 19660 19392 19712
rect 19800 19660 19852 19712
rect 21364 19660 21416 19712
rect 22100 19737 22109 19771
rect 22109 19737 22143 19771
rect 22143 19737 22152 19771
rect 22100 19728 22152 19737
rect 22928 19728 22980 19780
rect 24860 19771 24912 19780
rect 23296 19660 23348 19712
rect 24860 19737 24869 19771
rect 24869 19737 24903 19771
rect 24903 19737 24912 19771
rect 24860 19728 24912 19737
rect 25872 19728 25924 19780
rect 26516 19728 26568 19780
rect 27896 19796 27948 19848
rect 31116 19932 31168 19984
rect 30196 19907 30248 19916
rect 30196 19873 30205 19907
rect 30205 19873 30239 19907
rect 30239 19873 30248 19907
rect 30196 19864 30248 19873
rect 30748 19907 30800 19916
rect 30748 19873 30757 19907
rect 30757 19873 30791 19907
rect 30791 19873 30800 19907
rect 30748 19864 30800 19873
rect 31576 19864 31628 19916
rect 27252 19660 27304 19712
rect 29736 19771 29788 19780
rect 29736 19737 29745 19771
rect 29745 19737 29779 19771
rect 29779 19737 29788 19771
rect 29736 19728 29788 19737
rect 30472 19796 30524 19848
rect 31116 19839 31168 19848
rect 31116 19805 31125 19839
rect 31125 19805 31159 19839
rect 31159 19805 31168 19839
rect 31116 19796 31168 19805
rect 28264 19703 28316 19712
rect 28264 19669 28273 19703
rect 28273 19669 28307 19703
rect 28307 19669 28316 19703
rect 28264 19660 28316 19669
rect 30012 19660 30064 19712
rect 30288 19660 30340 19712
rect 30472 19660 30524 19712
rect 8632 19558 8684 19610
rect 8696 19558 8748 19610
rect 8760 19558 8812 19610
rect 8824 19558 8876 19610
rect 8888 19558 8940 19610
rect 16314 19558 16366 19610
rect 16378 19558 16430 19610
rect 16442 19558 16494 19610
rect 16506 19558 16558 19610
rect 16570 19558 16622 19610
rect 23996 19558 24048 19610
rect 24060 19558 24112 19610
rect 24124 19558 24176 19610
rect 24188 19558 24240 19610
rect 24252 19558 24304 19610
rect 31678 19558 31730 19610
rect 31742 19558 31794 19610
rect 31806 19558 31858 19610
rect 31870 19558 31922 19610
rect 31934 19558 31986 19610
rect 9036 19456 9088 19508
rect 11428 19456 11480 19508
rect 12164 19456 12216 19508
rect 13268 19456 13320 19508
rect 14096 19456 14148 19508
rect 16764 19456 16816 19508
rect 16948 19456 17000 19508
rect 17960 19456 18012 19508
rect 18880 19456 18932 19508
rect 19156 19499 19208 19508
rect 19156 19465 19165 19499
rect 19165 19465 19199 19499
rect 19199 19465 19208 19499
rect 19156 19456 19208 19465
rect 8024 19388 8076 19440
rect 9496 19388 9548 19440
rect 11336 19388 11388 19440
rect 11520 19388 11572 19440
rect 11704 19388 11756 19440
rect 12072 19431 12124 19440
rect 12072 19397 12081 19431
rect 12081 19397 12115 19431
rect 12115 19397 12124 19431
rect 12072 19388 12124 19397
rect 10876 19320 10928 19372
rect 9588 19252 9640 19304
rect 10048 19252 10100 19304
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 12532 19388 12584 19440
rect 12900 19431 12952 19440
rect 12900 19397 12909 19431
rect 12909 19397 12943 19431
rect 12943 19397 12952 19431
rect 12900 19388 12952 19397
rect 13176 19388 13228 19440
rect 12348 19320 12400 19372
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 12808 19320 12860 19372
rect 13084 19320 13136 19372
rect 11336 19252 11388 19304
rect 12900 19252 12952 19304
rect 13176 19252 13228 19304
rect 13728 19388 13780 19440
rect 17316 19388 17368 19440
rect 17408 19388 17460 19440
rect 13636 19363 13688 19372
rect 13636 19329 13645 19363
rect 13645 19329 13679 19363
rect 13679 19329 13688 19363
rect 13636 19320 13688 19329
rect 14280 19363 14332 19372
rect 14280 19329 14289 19363
rect 14289 19329 14323 19363
rect 14323 19329 14332 19363
rect 14280 19320 14332 19329
rect 14740 19320 14792 19372
rect 15844 19363 15896 19372
rect 15844 19329 15853 19363
rect 15853 19329 15887 19363
rect 15887 19329 15896 19363
rect 15844 19320 15896 19329
rect 15936 19320 15988 19372
rect 16304 19363 16356 19372
rect 16304 19329 16313 19363
rect 16313 19329 16347 19363
rect 16347 19329 16356 19363
rect 16304 19320 16356 19329
rect 17040 19363 17092 19372
rect 9680 19184 9732 19236
rect 9772 19184 9824 19236
rect 13728 19184 13780 19236
rect 13912 19252 13964 19304
rect 15200 19252 15252 19304
rect 15476 19252 15528 19304
rect 16764 19252 16816 19304
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 17224 19320 17276 19372
rect 17500 19320 17552 19372
rect 18420 19388 18472 19440
rect 19616 19456 19668 19508
rect 20628 19456 20680 19508
rect 20812 19456 20864 19508
rect 17960 19320 18012 19372
rect 18328 19320 18380 19372
rect 18788 19363 18840 19372
rect 15292 19227 15344 19236
rect 6000 19116 6052 19168
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 6644 19116 6696 19125
rect 7656 19159 7708 19168
rect 7656 19125 7665 19159
rect 7665 19125 7699 19159
rect 7699 19125 7708 19159
rect 7656 19116 7708 19125
rect 9220 19116 9272 19168
rect 9864 19116 9916 19168
rect 10784 19116 10836 19168
rect 11520 19116 11572 19168
rect 13268 19116 13320 19168
rect 13360 19116 13412 19168
rect 14924 19159 14976 19168
rect 14924 19125 14933 19159
rect 14933 19125 14967 19159
rect 14967 19125 14976 19159
rect 14924 19116 14976 19125
rect 15292 19193 15301 19227
rect 15301 19193 15335 19227
rect 15335 19193 15344 19227
rect 15292 19184 15344 19193
rect 15384 19184 15436 19236
rect 16856 19184 16908 19236
rect 17776 19295 17828 19304
rect 17776 19261 17785 19295
rect 17785 19261 17819 19295
rect 17819 19261 17828 19295
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 19984 19388 20036 19440
rect 21272 19456 21324 19508
rect 22652 19456 22704 19508
rect 23204 19456 23256 19508
rect 23388 19456 23440 19508
rect 25412 19456 25464 19508
rect 25596 19456 25648 19508
rect 26608 19456 26660 19508
rect 26700 19456 26752 19508
rect 27436 19456 27488 19508
rect 27528 19456 27580 19508
rect 27804 19456 27856 19508
rect 28448 19456 28500 19508
rect 22192 19388 22244 19440
rect 23848 19388 23900 19440
rect 25688 19388 25740 19440
rect 26332 19388 26384 19440
rect 28632 19456 28684 19508
rect 32312 19456 32364 19508
rect 22100 19320 22152 19372
rect 26976 19320 27028 19372
rect 27252 19320 27304 19372
rect 27436 19320 27488 19372
rect 27804 19363 27856 19372
rect 27804 19329 27813 19363
rect 27813 19329 27847 19363
rect 27847 19329 27856 19363
rect 27804 19320 27856 19329
rect 28172 19320 28224 19372
rect 29920 19388 29972 19440
rect 30288 19388 30340 19440
rect 29000 19320 29052 19372
rect 30472 19363 30524 19372
rect 30472 19329 30481 19363
rect 30481 19329 30515 19363
rect 30515 19329 30524 19363
rect 32220 19388 32272 19440
rect 30472 19320 30524 19329
rect 17776 19252 17828 19261
rect 18328 19184 18380 19236
rect 18144 19116 18196 19168
rect 18420 19116 18472 19168
rect 18604 19252 18656 19304
rect 19156 19252 19208 19304
rect 19898 19295 19950 19304
rect 19898 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19950 19295
rect 19064 19184 19116 19236
rect 19898 19252 19950 19261
rect 20352 19252 20404 19304
rect 21456 19252 21508 19304
rect 21180 19184 21232 19236
rect 21272 19116 21324 19168
rect 21732 19116 21784 19168
rect 27896 19252 27948 19304
rect 29184 19252 29236 19304
rect 29460 19252 29512 19304
rect 29920 19252 29972 19304
rect 30288 19252 30340 19304
rect 24860 19227 24912 19236
rect 24860 19193 24869 19227
rect 24869 19193 24903 19227
rect 24903 19193 24912 19227
rect 24860 19184 24912 19193
rect 26700 19184 26752 19236
rect 27252 19184 27304 19236
rect 27620 19184 27672 19236
rect 28172 19184 28224 19236
rect 24032 19159 24084 19168
rect 24032 19125 24041 19159
rect 24041 19125 24075 19159
rect 24075 19125 24084 19159
rect 24032 19116 24084 19125
rect 24216 19116 24268 19168
rect 26240 19116 26292 19168
rect 30748 19184 30800 19236
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 29184 19116 29236 19168
rect 30656 19116 30708 19168
rect 30932 19159 30984 19168
rect 30932 19125 30941 19159
rect 30941 19125 30975 19159
rect 30975 19125 30984 19159
rect 30932 19116 30984 19125
rect 4791 19014 4843 19066
rect 4855 19014 4907 19066
rect 4919 19014 4971 19066
rect 4983 19014 5035 19066
rect 5047 19014 5099 19066
rect 12473 19014 12525 19066
rect 12537 19014 12589 19066
rect 12601 19014 12653 19066
rect 12665 19014 12717 19066
rect 12729 19014 12781 19066
rect 20155 19014 20207 19066
rect 20219 19014 20271 19066
rect 20283 19014 20335 19066
rect 20347 19014 20399 19066
rect 20411 19014 20463 19066
rect 27837 19014 27889 19066
rect 27901 19014 27953 19066
rect 27965 19014 28017 19066
rect 28029 19014 28081 19066
rect 28093 19014 28145 19066
rect 12256 18912 12308 18964
rect 13728 18912 13780 18964
rect 14280 18912 14332 18964
rect 15016 18912 15068 18964
rect 15476 18912 15528 18964
rect 15936 18912 15988 18964
rect 12624 18844 12676 18896
rect 13452 18887 13504 18896
rect 13452 18853 13461 18887
rect 13461 18853 13495 18887
rect 13495 18853 13504 18887
rect 13452 18844 13504 18853
rect 13544 18844 13596 18896
rect 17132 18844 17184 18896
rect 9956 18819 10008 18828
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 10968 18776 11020 18828
rect 11060 18776 11112 18828
rect 1584 18751 1636 18760
rect 1584 18717 1593 18751
rect 1593 18717 1627 18751
rect 1627 18717 1636 18751
rect 1584 18708 1636 18717
rect 10048 18640 10100 18692
rect 7932 18615 7984 18624
rect 7932 18581 7941 18615
rect 7941 18581 7975 18615
rect 7975 18581 7984 18615
rect 7932 18572 7984 18581
rect 9220 18572 9272 18624
rect 11336 18708 11388 18760
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 12256 18708 12308 18760
rect 12992 18708 13044 18760
rect 13268 18776 13320 18828
rect 14004 18776 14056 18828
rect 15660 18776 15712 18828
rect 17500 18912 17552 18964
rect 17776 18912 17828 18964
rect 19340 18912 19392 18964
rect 19616 18912 19668 18964
rect 19984 18912 20036 18964
rect 18144 18844 18196 18896
rect 18328 18844 18380 18896
rect 11152 18640 11204 18692
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 16120 18708 16172 18760
rect 16212 18708 16264 18760
rect 16856 18708 16908 18760
rect 14924 18683 14976 18692
rect 14924 18649 14933 18683
rect 14933 18649 14967 18683
rect 14967 18649 14976 18683
rect 14924 18640 14976 18649
rect 15108 18683 15160 18692
rect 15108 18649 15117 18683
rect 15117 18649 15151 18683
rect 15151 18649 15160 18683
rect 15108 18640 15160 18649
rect 15568 18683 15620 18692
rect 15568 18649 15577 18683
rect 15577 18649 15611 18683
rect 15611 18649 15620 18683
rect 15568 18640 15620 18649
rect 16028 18640 16080 18692
rect 10968 18615 11020 18624
rect 10968 18581 10977 18615
rect 10977 18581 11011 18615
rect 11011 18581 11020 18615
rect 10968 18572 11020 18581
rect 11428 18572 11480 18624
rect 12072 18572 12124 18624
rect 12808 18572 12860 18624
rect 13544 18572 13596 18624
rect 13728 18572 13780 18624
rect 17132 18640 17184 18692
rect 17868 18776 17920 18828
rect 18420 18819 18472 18828
rect 17408 18708 17460 18760
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 17776 18708 17828 18760
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 20904 18912 20956 18964
rect 21824 18912 21876 18964
rect 22468 18887 22520 18896
rect 22468 18853 22477 18887
rect 22477 18853 22511 18887
rect 22511 18853 22520 18887
rect 22468 18844 22520 18853
rect 22744 18844 22796 18896
rect 20352 18776 20404 18828
rect 23204 18776 23256 18828
rect 26332 18912 26384 18964
rect 26976 18912 27028 18964
rect 24952 18844 25004 18896
rect 27436 18887 27488 18896
rect 26332 18819 26384 18828
rect 26332 18785 26341 18819
rect 26341 18785 26375 18819
rect 26375 18785 26384 18819
rect 26332 18776 26384 18785
rect 26608 18776 26660 18828
rect 26792 18819 26844 18828
rect 26792 18785 26801 18819
rect 26801 18785 26835 18819
rect 26835 18785 26844 18819
rect 26792 18776 26844 18785
rect 27436 18853 27445 18887
rect 27445 18853 27479 18887
rect 27479 18853 27488 18887
rect 27436 18844 27488 18853
rect 27712 18912 27764 18964
rect 28080 18912 28132 18964
rect 27896 18776 27948 18828
rect 27988 18776 28040 18828
rect 28356 18912 28408 18964
rect 28448 18912 28500 18964
rect 29552 18912 29604 18964
rect 28540 18776 28592 18828
rect 31116 18844 31168 18896
rect 30012 18776 30064 18828
rect 30932 18776 30984 18828
rect 18052 18708 18104 18760
rect 18788 18708 18840 18760
rect 18880 18708 18932 18760
rect 19616 18708 19668 18760
rect 21640 18708 21692 18760
rect 16488 18572 16540 18624
rect 18880 18572 18932 18624
rect 20536 18640 20588 18692
rect 21272 18640 21324 18692
rect 22008 18683 22060 18692
rect 22008 18649 22017 18683
rect 22017 18649 22051 18683
rect 22051 18649 22060 18683
rect 22008 18640 22060 18649
rect 24216 18708 24268 18760
rect 24952 18708 25004 18760
rect 27436 18708 27488 18760
rect 30104 18751 30156 18760
rect 21824 18572 21876 18624
rect 22284 18572 22336 18624
rect 23664 18572 23716 18624
rect 26148 18640 26200 18692
rect 25228 18572 25280 18624
rect 25964 18572 26016 18624
rect 26976 18640 27028 18692
rect 26792 18572 26844 18624
rect 28080 18640 28132 18692
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 30748 18751 30800 18760
rect 30748 18717 30757 18751
rect 30757 18717 30791 18751
rect 30791 18717 30800 18751
rect 30748 18708 30800 18717
rect 31668 18708 31720 18760
rect 30656 18640 30708 18692
rect 32496 18640 32548 18692
rect 28448 18572 28500 18624
rect 29184 18572 29236 18624
rect 29368 18572 29420 18624
rect 8632 18470 8684 18522
rect 8696 18470 8748 18522
rect 8760 18470 8812 18522
rect 8824 18470 8876 18522
rect 8888 18470 8940 18522
rect 16314 18470 16366 18522
rect 16378 18470 16430 18522
rect 16442 18470 16494 18522
rect 16506 18470 16558 18522
rect 16570 18470 16622 18522
rect 23996 18470 24048 18522
rect 24060 18470 24112 18522
rect 24124 18470 24176 18522
rect 24188 18470 24240 18522
rect 24252 18470 24304 18522
rect 31678 18470 31730 18522
rect 31742 18470 31794 18522
rect 31806 18470 31858 18522
rect 31870 18470 31922 18522
rect 31934 18470 31986 18522
rect 10048 18411 10100 18420
rect 10048 18377 10057 18411
rect 10057 18377 10091 18411
rect 10091 18377 10100 18411
rect 10048 18368 10100 18377
rect 15016 18368 15068 18420
rect 15476 18368 15528 18420
rect 11520 18300 11572 18352
rect 11796 18300 11848 18352
rect 9588 18232 9640 18284
rect 11244 18232 11296 18284
rect 14096 18300 14148 18352
rect 14280 18300 14332 18352
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 14464 18300 14516 18352
rect 14924 18300 14976 18352
rect 13636 18232 13688 18241
rect 10876 18164 10928 18216
rect 12624 18164 12676 18216
rect 14004 18164 14056 18216
rect 6644 18096 6696 18148
rect 9864 18096 9916 18148
rect 11060 18096 11112 18148
rect 12256 18096 12308 18148
rect 13912 18096 13964 18148
rect 14556 18232 14608 18284
rect 16028 18368 16080 18420
rect 17224 18368 17276 18420
rect 14188 18164 14240 18216
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 16580 18300 16632 18352
rect 16856 18300 16908 18352
rect 17316 18300 17368 18352
rect 17684 18343 17736 18352
rect 17684 18309 17693 18343
rect 17693 18309 17727 18343
rect 17727 18309 17736 18343
rect 17684 18300 17736 18309
rect 18328 18368 18380 18420
rect 17960 18300 18012 18352
rect 18144 18300 18196 18352
rect 19340 18300 19392 18352
rect 19892 18343 19944 18352
rect 19892 18309 19901 18343
rect 19901 18309 19935 18343
rect 19935 18309 19944 18343
rect 19892 18300 19944 18309
rect 19984 18300 20036 18352
rect 21456 18368 21508 18420
rect 25780 18368 25832 18420
rect 26884 18368 26936 18420
rect 21824 18300 21876 18352
rect 22192 18300 22244 18352
rect 22744 18300 22796 18352
rect 23572 18300 23624 18352
rect 16120 18164 16172 18216
rect 16396 18164 16448 18216
rect 19156 18232 19208 18284
rect 19616 18275 19668 18284
rect 19616 18241 19625 18275
rect 19625 18241 19659 18275
rect 19659 18241 19668 18275
rect 19616 18232 19668 18241
rect 23756 18232 23808 18284
rect 24400 18232 24452 18284
rect 25044 18232 25096 18284
rect 26148 18300 26200 18352
rect 26240 18300 26292 18352
rect 26700 18300 26752 18352
rect 17684 18164 17736 18216
rect 14464 18096 14516 18148
rect 18052 18096 18104 18148
rect 21640 18164 21692 18216
rect 21088 18096 21140 18148
rect 22376 18164 22428 18216
rect 23020 18164 23072 18216
rect 25320 18164 25372 18216
rect 25780 18164 25832 18216
rect 25964 18207 26016 18216
rect 25964 18173 25973 18207
rect 25973 18173 26007 18207
rect 26007 18173 26016 18207
rect 25964 18164 26016 18173
rect 26976 18232 27028 18284
rect 27436 18275 27488 18284
rect 27436 18241 27445 18275
rect 27445 18241 27479 18275
rect 27479 18241 27488 18275
rect 27436 18232 27488 18241
rect 27712 18411 27764 18420
rect 27712 18377 27721 18411
rect 27721 18377 27755 18411
rect 27755 18377 27764 18411
rect 27712 18368 27764 18377
rect 30196 18368 30248 18420
rect 30840 18368 30892 18420
rect 27896 18300 27948 18352
rect 27988 18232 28040 18284
rect 28264 18232 28316 18284
rect 28448 18232 28500 18284
rect 23480 18096 23532 18148
rect 26516 18096 26568 18148
rect 28080 18164 28132 18216
rect 28172 18207 28224 18216
rect 28172 18173 28181 18207
rect 28181 18173 28215 18207
rect 28215 18173 28224 18207
rect 28172 18164 28224 18173
rect 28816 18164 28868 18216
rect 32772 18300 32824 18352
rect 29000 18232 29052 18284
rect 29184 18164 29236 18216
rect 29460 18275 29512 18284
rect 29460 18241 29469 18275
rect 29469 18241 29503 18275
rect 29503 18241 29512 18275
rect 29644 18275 29696 18284
rect 29460 18232 29512 18241
rect 29644 18241 29653 18275
rect 29653 18241 29687 18275
rect 29687 18241 29696 18275
rect 29644 18232 29696 18241
rect 30012 18232 30064 18284
rect 30196 18275 30248 18284
rect 30196 18241 30205 18275
rect 30205 18241 30239 18275
rect 30239 18241 30248 18275
rect 30196 18232 30248 18241
rect 30472 18232 30524 18284
rect 31668 18232 31720 18284
rect 30288 18164 30340 18216
rect 32404 18164 32456 18216
rect 27804 18096 27856 18148
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 9496 18071 9548 18080
rect 9496 18037 9505 18071
rect 9505 18037 9539 18071
rect 9539 18037 9548 18071
rect 9496 18028 9548 18037
rect 10876 18028 10928 18080
rect 11244 18028 11296 18080
rect 12164 18028 12216 18080
rect 13728 18028 13780 18080
rect 13820 18028 13872 18080
rect 14832 18028 14884 18080
rect 15016 18071 15068 18080
rect 15016 18037 15025 18071
rect 15025 18037 15059 18071
rect 15059 18037 15068 18071
rect 15016 18028 15068 18037
rect 15154 18028 15206 18080
rect 15292 18028 15344 18080
rect 15660 18028 15712 18080
rect 15936 18028 15988 18080
rect 16304 18028 16356 18080
rect 17408 18028 17460 18080
rect 20352 18028 20404 18080
rect 21824 18028 21876 18080
rect 22928 18028 22980 18080
rect 23756 18071 23808 18080
rect 23756 18037 23765 18071
rect 23765 18037 23799 18071
rect 23799 18037 23808 18071
rect 23756 18028 23808 18037
rect 24676 18071 24728 18080
rect 24676 18037 24685 18071
rect 24685 18037 24719 18071
rect 24719 18037 24728 18071
rect 24676 18028 24728 18037
rect 29828 18096 29880 18148
rect 30748 18096 30800 18148
rect 32220 18096 32272 18148
rect 29276 18028 29328 18080
rect 32312 18028 32364 18080
rect 4791 17926 4843 17978
rect 4855 17926 4907 17978
rect 4919 17926 4971 17978
rect 4983 17926 5035 17978
rect 5047 17926 5099 17978
rect 12473 17926 12525 17978
rect 12537 17926 12589 17978
rect 12601 17926 12653 17978
rect 12665 17926 12717 17978
rect 12729 17926 12781 17978
rect 20155 17926 20207 17978
rect 20219 17926 20271 17978
rect 20283 17926 20335 17978
rect 20347 17926 20399 17978
rect 20411 17926 20463 17978
rect 27837 17926 27889 17978
rect 27901 17926 27953 17978
rect 27965 17926 28017 17978
rect 28029 17926 28081 17978
rect 28093 17926 28145 17978
rect 9956 17824 10008 17876
rect 14556 17824 14608 17876
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 15108 17756 15160 17808
rect 15200 17756 15252 17808
rect 12992 17688 13044 17740
rect 15568 17824 15620 17876
rect 15936 17824 15988 17876
rect 16672 17824 16724 17876
rect 16856 17824 16908 17876
rect 17960 17824 18012 17876
rect 22008 17824 22060 17876
rect 23112 17824 23164 17876
rect 25044 17824 25096 17876
rect 25504 17824 25556 17876
rect 26884 17824 26936 17876
rect 28172 17867 28224 17876
rect 16120 17756 16172 17808
rect 15568 17688 15620 17740
rect 16580 17756 16632 17808
rect 17592 17756 17644 17808
rect 19616 17756 19668 17808
rect 21088 17756 21140 17808
rect 19248 17688 19300 17740
rect 22376 17731 22428 17740
rect 22376 17697 22385 17731
rect 22385 17697 22419 17731
rect 22419 17697 22428 17731
rect 22376 17688 22428 17697
rect 22468 17688 22520 17740
rect 15016 17620 15068 17672
rect 15752 17620 15804 17672
rect 15844 17620 15896 17672
rect 16304 17663 16356 17672
rect 16304 17629 16321 17663
rect 16321 17629 16356 17663
rect 16304 17620 16356 17629
rect 13452 17552 13504 17604
rect 13636 17595 13688 17604
rect 13636 17561 13645 17595
rect 13645 17561 13679 17595
rect 13679 17561 13688 17595
rect 13636 17552 13688 17561
rect 14280 17552 14332 17604
rect 14556 17595 14608 17604
rect 14556 17561 14565 17595
rect 14565 17561 14599 17595
rect 14599 17561 14608 17595
rect 14556 17552 14608 17561
rect 9864 17527 9916 17536
rect 9864 17493 9873 17527
rect 9873 17493 9907 17527
rect 9907 17493 9916 17527
rect 9864 17484 9916 17493
rect 10416 17527 10468 17536
rect 10416 17493 10425 17527
rect 10425 17493 10459 17527
rect 10459 17493 10468 17527
rect 10416 17484 10468 17493
rect 11612 17527 11664 17536
rect 11612 17493 11621 17527
rect 11621 17493 11655 17527
rect 11655 17493 11664 17527
rect 11612 17484 11664 17493
rect 12992 17527 13044 17536
rect 12992 17493 13001 17527
rect 13001 17493 13035 17527
rect 13035 17493 13044 17527
rect 12992 17484 13044 17493
rect 13268 17484 13320 17536
rect 13728 17484 13780 17536
rect 15200 17527 15252 17536
rect 15200 17493 15209 17527
rect 15209 17493 15243 17527
rect 15243 17493 15252 17527
rect 15200 17484 15252 17493
rect 15568 17552 15620 17604
rect 15936 17552 15988 17604
rect 17316 17620 17368 17672
rect 19340 17620 19392 17672
rect 16764 17552 16816 17604
rect 16948 17552 17000 17604
rect 19800 17663 19852 17672
rect 19800 17629 19809 17663
rect 19809 17629 19843 17663
rect 19843 17629 19852 17663
rect 19800 17620 19852 17629
rect 20720 17620 20772 17672
rect 20996 17620 21048 17672
rect 22652 17688 22704 17740
rect 23572 17756 23624 17808
rect 22928 17688 22980 17740
rect 16212 17484 16264 17536
rect 17684 17484 17736 17536
rect 17960 17484 18012 17536
rect 18236 17484 18288 17536
rect 19524 17484 19576 17536
rect 20168 17552 20220 17604
rect 20812 17552 20864 17604
rect 19708 17484 19760 17536
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 20720 17484 20772 17536
rect 22652 17484 22704 17536
rect 25228 17663 25280 17672
rect 24584 17527 24636 17536
rect 24584 17493 24593 17527
rect 24593 17493 24627 17527
rect 24627 17493 24636 17527
rect 24584 17484 24636 17493
rect 25228 17629 25237 17663
rect 25237 17629 25271 17663
rect 25271 17629 25280 17663
rect 25228 17620 25280 17629
rect 25596 17756 25648 17808
rect 28172 17833 28181 17867
rect 28181 17833 28215 17867
rect 28215 17833 28224 17867
rect 28172 17824 28224 17833
rect 30472 17824 30524 17876
rect 28356 17756 28408 17808
rect 30748 17756 30800 17808
rect 25504 17688 25556 17740
rect 25780 17688 25832 17740
rect 26148 17688 26200 17740
rect 26516 17688 26568 17740
rect 26056 17663 26108 17672
rect 26056 17629 26065 17663
rect 26065 17629 26099 17663
rect 26099 17629 26108 17663
rect 26056 17620 26108 17629
rect 27620 17688 27672 17740
rect 27712 17731 27764 17740
rect 27712 17697 27721 17731
rect 27721 17697 27755 17731
rect 27755 17697 27764 17731
rect 27712 17688 27764 17697
rect 29552 17688 29604 17740
rect 29736 17688 29788 17740
rect 31300 17688 31352 17740
rect 27436 17620 27488 17672
rect 28080 17663 28132 17672
rect 28080 17629 28089 17663
rect 28089 17629 28123 17663
rect 28123 17629 28132 17663
rect 28080 17620 28132 17629
rect 29092 17620 29144 17672
rect 30472 17620 30524 17672
rect 30748 17620 30800 17672
rect 25780 17552 25832 17604
rect 26148 17552 26200 17604
rect 26240 17595 26292 17604
rect 26240 17561 26249 17595
rect 26249 17561 26283 17595
rect 26283 17561 26292 17595
rect 26240 17552 26292 17561
rect 26792 17552 26844 17604
rect 26976 17595 27028 17604
rect 26976 17561 26985 17595
rect 26985 17561 27019 17595
rect 27019 17561 27028 17595
rect 26976 17552 27028 17561
rect 25964 17527 26016 17536
rect 25964 17493 25973 17527
rect 25973 17493 26007 17527
rect 26007 17493 26016 17527
rect 25964 17484 26016 17493
rect 26700 17527 26752 17536
rect 26700 17493 26709 17527
rect 26709 17493 26743 17527
rect 26743 17493 26752 17527
rect 26700 17484 26752 17493
rect 27528 17552 27580 17604
rect 29368 17552 29420 17604
rect 29736 17552 29788 17604
rect 31576 17552 31628 17604
rect 28264 17484 28316 17536
rect 28540 17484 28592 17536
rect 29276 17484 29328 17536
rect 30012 17484 30064 17536
rect 31300 17484 31352 17536
rect 31668 17484 31720 17536
rect 8632 17382 8684 17434
rect 8696 17382 8748 17434
rect 8760 17382 8812 17434
rect 8824 17382 8876 17434
rect 8888 17382 8940 17434
rect 16314 17382 16366 17434
rect 16378 17382 16430 17434
rect 16442 17382 16494 17434
rect 16506 17382 16558 17434
rect 16570 17382 16622 17434
rect 23996 17382 24048 17434
rect 24060 17382 24112 17434
rect 24124 17382 24176 17434
rect 24188 17382 24240 17434
rect 24252 17382 24304 17434
rect 31678 17382 31730 17434
rect 31742 17382 31794 17434
rect 31806 17382 31858 17434
rect 31870 17382 31922 17434
rect 31934 17382 31986 17434
rect 10968 17280 11020 17332
rect 13636 17280 13688 17332
rect 12900 17212 12952 17264
rect 13176 17212 13228 17264
rect 13268 17255 13320 17264
rect 13268 17221 13293 17255
rect 13293 17221 13320 17255
rect 13268 17212 13320 17221
rect 14096 17323 14148 17332
rect 14096 17289 14121 17323
rect 14121 17289 14148 17323
rect 14096 17280 14148 17289
rect 15200 17280 15252 17332
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 11336 17144 11388 17196
rect 12348 17187 12400 17196
rect 12348 17153 12357 17187
rect 12357 17153 12391 17187
rect 12391 17153 12400 17187
rect 12348 17144 12400 17153
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 15476 17212 15528 17264
rect 16948 17280 17000 17332
rect 17500 17280 17552 17332
rect 18972 17280 19024 17332
rect 19432 17280 19484 17332
rect 14648 17144 14700 17196
rect 14924 17144 14976 17196
rect 15016 17144 15068 17196
rect 15384 17144 15436 17196
rect 11520 17076 11572 17128
rect 9680 17008 9732 17060
rect 12256 17008 12308 17060
rect 13176 17008 13228 17060
rect 15292 17076 15344 17128
rect 16672 17144 16724 17196
rect 17408 17212 17460 17264
rect 17776 17212 17828 17264
rect 18328 17212 18380 17264
rect 20628 17212 20680 17264
rect 20812 17212 20864 17264
rect 23940 17280 23992 17332
rect 24492 17280 24544 17332
rect 21732 17212 21784 17264
rect 22928 17212 22980 17264
rect 24676 17212 24728 17264
rect 25044 17212 25096 17264
rect 26516 17212 26568 17264
rect 26700 17212 26752 17264
rect 16488 17076 16540 17128
rect 16580 17076 16632 17128
rect 15844 17008 15896 17060
rect 17408 17076 17460 17128
rect 17868 17076 17920 17128
rect 17960 17076 18012 17128
rect 17040 17051 17092 17060
rect 17040 17017 17049 17051
rect 17049 17017 17083 17051
rect 17083 17017 17092 17051
rect 17040 17008 17092 17017
rect 18420 17076 18472 17128
rect 18512 17076 18564 17128
rect 21088 17144 21140 17196
rect 24032 17144 24084 17196
rect 28172 17280 28224 17332
rect 28540 17280 28592 17332
rect 28908 17280 28960 17332
rect 29184 17280 29236 17332
rect 22836 17076 22888 17128
rect 23020 17076 23072 17128
rect 10508 16983 10560 16992
rect 10508 16949 10517 16983
rect 10517 16949 10551 16983
rect 10551 16949 10560 16983
rect 10508 16940 10560 16949
rect 12164 16940 12216 16992
rect 13728 16940 13780 16992
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 14280 16983 14332 16992
rect 14280 16949 14289 16983
rect 14289 16949 14323 16983
rect 14323 16949 14332 16983
rect 14280 16940 14332 16949
rect 15108 16940 15160 16992
rect 15200 16983 15252 16992
rect 15200 16949 15209 16983
rect 15209 16949 15243 16983
rect 15243 16949 15252 16983
rect 15200 16940 15252 16949
rect 15660 16940 15712 16992
rect 16028 16940 16080 16992
rect 20812 17008 20864 17060
rect 21180 17008 21232 17060
rect 21640 17008 21692 17060
rect 17684 16940 17736 16992
rect 18144 16940 18196 16992
rect 18328 16940 18380 16992
rect 19064 16940 19116 16992
rect 21456 16940 21508 16992
rect 22008 16940 22060 16992
rect 22468 16940 22520 16992
rect 25320 17076 25372 17128
rect 26056 17119 26108 17128
rect 26056 17085 26065 17119
rect 26065 17085 26099 17119
rect 26099 17085 26108 17119
rect 26056 17076 26108 17085
rect 26700 17076 26752 17128
rect 27436 17212 27488 17264
rect 27712 17212 27764 17264
rect 28356 17144 28408 17196
rect 29184 17144 29236 17196
rect 30012 17255 30064 17264
rect 29368 17144 29420 17196
rect 25596 17008 25648 17060
rect 26516 17051 26568 17060
rect 26516 17017 26525 17051
rect 26525 17017 26559 17051
rect 26559 17017 26568 17051
rect 29460 17076 29512 17128
rect 30012 17221 30021 17255
rect 30021 17221 30055 17255
rect 30055 17221 30064 17255
rect 30012 17212 30064 17221
rect 30472 17280 30524 17332
rect 29828 17144 29880 17196
rect 30472 17144 30524 17196
rect 32128 17076 32180 17128
rect 26516 17008 26568 17017
rect 27528 17008 27580 17060
rect 28264 17051 28316 17060
rect 28264 17017 28273 17051
rect 28273 17017 28307 17051
rect 28307 17017 28316 17051
rect 28264 17008 28316 17017
rect 29000 17008 29052 17060
rect 29184 17051 29236 17060
rect 29184 17017 29193 17051
rect 29193 17017 29227 17051
rect 29227 17017 29236 17051
rect 29184 17008 29236 17017
rect 30472 16940 30524 16992
rect 31668 16940 31720 16992
rect 4791 16838 4843 16890
rect 4855 16838 4907 16890
rect 4919 16838 4971 16890
rect 4983 16838 5035 16890
rect 5047 16838 5099 16890
rect 12473 16838 12525 16890
rect 12537 16838 12589 16890
rect 12601 16838 12653 16890
rect 12665 16838 12717 16890
rect 12729 16838 12781 16890
rect 20155 16838 20207 16890
rect 20219 16838 20271 16890
rect 20283 16838 20335 16890
rect 20347 16838 20399 16890
rect 20411 16838 20463 16890
rect 27837 16838 27889 16890
rect 27901 16838 27953 16890
rect 27965 16838 28017 16890
rect 28029 16838 28081 16890
rect 28093 16838 28145 16890
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 11612 16736 11664 16788
rect 13452 16736 13504 16788
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 15844 16736 15896 16788
rect 16212 16736 16264 16788
rect 9864 16668 9916 16720
rect 10416 16711 10468 16720
rect 10416 16677 10425 16711
rect 10425 16677 10459 16711
rect 10459 16677 10468 16711
rect 10416 16668 10468 16677
rect 12992 16711 13044 16720
rect 12992 16677 13001 16711
rect 13001 16677 13035 16711
rect 13035 16677 13044 16711
rect 12992 16668 13044 16677
rect 13728 16711 13780 16720
rect 13728 16677 13737 16711
rect 13737 16677 13771 16711
rect 13771 16677 13780 16711
rect 13728 16668 13780 16677
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 10968 16600 11020 16652
rect 11612 16643 11664 16652
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 11244 16532 11296 16584
rect 12164 16600 12216 16652
rect 12624 16464 12676 16516
rect 12716 16464 12768 16516
rect 12992 16396 13044 16448
rect 13360 16532 13412 16584
rect 14188 16532 14240 16584
rect 14464 16532 14516 16584
rect 15200 16668 15252 16720
rect 18880 16711 18932 16720
rect 15108 16600 15160 16652
rect 18880 16677 18889 16711
rect 18889 16677 18923 16711
rect 18923 16677 18932 16711
rect 18880 16668 18932 16677
rect 19800 16736 19852 16788
rect 21456 16736 21508 16788
rect 21548 16736 21600 16788
rect 23480 16736 23532 16788
rect 23940 16779 23992 16788
rect 23940 16745 23949 16779
rect 23949 16745 23983 16779
rect 23983 16745 23992 16779
rect 23940 16736 23992 16745
rect 24032 16736 24084 16788
rect 26424 16736 26476 16788
rect 26884 16736 26936 16788
rect 28448 16736 28500 16788
rect 14832 16532 14884 16584
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15200 16532 15252 16584
rect 13360 16396 13412 16448
rect 14648 16464 14700 16516
rect 15936 16532 15988 16584
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16212 16575 16264 16584
rect 16028 16532 16080 16541
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 17960 16600 18012 16652
rect 22008 16668 22060 16720
rect 25596 16668 25648 16720
rect 26332 16668 26384 16720
rect 23480 16600 23532 16652
rect 16580 16532 16632 16584
rect 16672 16532 16724 16584
rect 16948 16532 17000 16584
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 19248 16532 19300 16584
rect 21364 16532 21416 16584
rect 14372 16396 14424 16448
rect 14464 16396 14516 16448
rect 15476 16396 15528 16448
rect 15660 16396 15712 16448
rect 16028 16396 16080 16448
rect 17684 16464 17736 16516
rect 17960 16464 18012 16516
rect 19340 16464 19392 16516
rect 19800 16464 19852 16516
rect 16488 16396 16540 16448
rect 21456 16464 21508 16516
rect 21364 16396 21416 16448
rect 23664 16532 23716 16584
rect 21824 16464 21876 16516
rect 22836 16464 22888 16516
rect 25320 16600 25372 16652
rect 25780 16600 25832 16652
rect 26056 16643 26108 16652
rect 26056 16609 26065 16643
rect 26065 16609 26099 16643
rect 26099 16609 26108 16643
rect 26056 16600 26108 16609
rect 26148 16643 26200 16652
rect 26148 16609 26157 16643
rect 26157 16609 26191 16643
rect 26191 16609 26200 16643
rect 26148 16600 26200 16609
rect 26976 16600 27028 16652
rect 28264 16668 28316 16720
rect 31300 16736 31352 16788
rect 27436 16600 27488 16652
rect 24860 16575 24912 16584
rect 24492 16464 24544 16516
rect 24860 16541 24869 16575
rect 24869 16541 24903 16575
rect 24903 16541 24912 16575
rect 24860 16532 24912 16541
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25964 16575 26016 16584
rect 25228 16532 25280 16541
rect 25964 16541 25973 16575
rect 25973 16541 26007 16575
rect 26007 16541 26016 16575
rect 25964 16532 26016 16541
rect 26608 16532 26660 16584
rect 27712 16532 27764 16584
rect 29000 16575 29052 16584
rect 24032 16396 24084 16448
rect 25320 16464 25372 16516
rect 26884 16396 26936 16448
rect 27068 16439 27120 16448
rect 27068 16405 27077 16439
rect 27077 16405 27111 16439
rect 27111 16405 27120 16439
rect 27068 16396 27120 16405
rect 27436 16396 27488 16448
rect 29000 16541 29009 16575
rect 29009 16541 29043 16575
rect 29043 16541 29052 16575
rect 29000 16532 29052 16541
rect 29184 16532 29236 16584
rect 28816 16464 28868 16516
rect 30656 16532 30708 16584
rect 31300 16464 31352 16516
rect 28448 16396 28500 16448
rect 29644 16396 29696 16448
rect 29736 16439 29788 16448
rect 29736 16405 29745 16439
rect 29745 16405 29779 16439
rect 29779 16405 29788 16439
rect 29736 16396 29788 16405
rect 30380 16396 30432 16448
rect 30656 16439 30708 16448
rect 30656 16405 30665 16439
rect 30665 16405 30699 16439
rect 30699 16405 30708 16439
rect 30656 16396 30708 16405
rect 8632 16294 8684 16346
rect 8696 16294 8748 16346
rect 8760 16294 8812 16346
rect 8824 16294 8876 16346
rect 8888 16294 8940 16346
rect 16314 16294 16366 16346
rect 16378 16294 16430 16346
rect 16442 16294 16494 16346
rect 16506 16294 16558 16346
rect 16570 16294 16622 16346
rect 23996 16294 24048 16346
rect 24060 16294 24112 16346
rect 24124 16294 24176 16346
rect 24188 16294 24240 16346
rect 24252 16294 24304 16346
rect 31678 16294 31730 16346
rect 31742 16294 31794 16346
rect 31806 16294 31858 16346
rect 31870 16294 31922 16346
rect 31934 16294 31986 16346
rect 10876 16192 10928 16244
rect 12348 16192 12400 16244
rect 14188 16192 14240 16244
rect 14740 16192 14792 16244
rect 15016 16192 15068 16244
rect 16396 16192 16448 16244
rect 16856 16192 16908 16244
rect 11244 16124 11296 16176
rect 16764 16124 16816 16176
rect 17868 16192 17920 16244
rect 18144 16192 18196 16244
rect 18880 16192 18932 16244
rect 19156 16192 19208 16244
rect 20536 16235 20588 16244
rect 11336 16056 11388 16108
rect 12992 16056 13044 16108
rect 13360 16056 13412 16108
rect 13820 16056 13872 16108
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 14556 16056 14608 16108
rect 15200 16056 15252 16108
rect 15752 16056 15804 16108
rect 19064 16124 19116 16176
rect 17776 16099 17828 16108
rect 15292 15988 15344 16040
rect 15476 15988 15528 16040
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 15844 15988 15896 16040
rect 16672 15988 16724 16040
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 18052 16056 18104 16108
rect 18328 16056 18380 16108
rect 20536 16201 20545 16235
rect 20545 16201 20579 16235
rect 20579 16201 20588 16235
rect 20536 16192 20588 16201
rect 23296 16192 23348 16244
rect 20628 16124 20680 16176
rect 22284 16167 22336 16176
rect 22284 16133 22293 16167
rect 22293 16133 22327 16167
rect 22327 16133 22336 16167
rect 22284 16124 22336 16133
rect 22560 16124 22612 16176
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 18696 15988 18748 16040
rect 19064 16031 19116 16040
rect 19064 15997 19073 16031
rect 19073 15997 19107 16031
rect 19107 15997 19116 16031
rect 19064 15988 19116 15997
rect 19156 15988 19208 16040
rect 20260 15988 20312 16040
rect 21180 16056 21232 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 24032 16192 24084 16244
rect 24860 16192 24912 16244
rect 26056 16192 26108 16244
rect 28356 16192 28408 16244
rect 29920 16192 29972 16244
rect 30104 16192 30156 16244
rect 31300 16192 31352 16244
rect 31668 16192 31720 16244
rect 23940 16124 23992 16176
rect 25044 16124 25096 16176
rect 26148 16124 26200 16176
rect 14096 15963 14148 15972
rect 14096 15929 14105 15963
rect 14105 15929 14139 15963
rect 14139 15929 14148 15963
rect 14096 15920 14148 15929
rect 14188 15963 14240 15972
rect 14188 15929 14197 15963
rect 14197 15929 14231 15963
rect 14231 15929 14240 15963
rect 14188 15920 14240 15929
rect 15384 15920 15436 15972
rect 16212 15920 16264 15972
rect 16580 15920 16632 15972
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 15476 15852 15528 15904
rect 15844 15852 15896 15904
rect 16120 15852 16172 15904
rect 16672 15852 16724 15904
rect 16856 15852 16908 15904
rect 17224 15852 17276 15904
rect 17500 15920 17552 15972
rect 18328 15920 18380 15972
rect 21548 15988 21600 16040
rect 22376 15988 22428 16040
rect 23756 15988 23808 16040
rect 26516 16056 26568 16108
rect 27436 16056 27488 16108
rect 27896 16124 27948 16176
rect 17684 15852 17736 15904
rect 18512 15852 18564 15904
rect 23388 15920 23440 15972
rect 23572 15920 23624 15972
rect 23664 15920 23716 15972
rect 26608 15988 26660 16040
rect 20260 15852 20312 15904
rect 27068 15920 27120 15972
rect 27896 15920 27948 15972
rect 25596 15852 25648 15904
rect 26240 15852 26292 15904
rect 28080 15920 28132 15972
rect 29644 16124 29696 16176
rect 30748 16124 30800 16176
rect 29184 16056 29236 16108
rect 29276 16056 29328 16108
rect 29368 15988 29420 16040
rect 29920 16056 29972 16108
rect 30196 15988 30248 16040
rect 29644 15920 29696 15972
rect 30748 15963 30800 15972
rect 30748 15929 30757 15963
rect 30757 15929 30791 15963
rect 30791 15929 30800 15963
rect 30748 15920 30800 15929
rect 29092 15852 29144 15904
rect 29368 15852 29420 15904
rect 4791 15750 4843 15802
rect 4855 15750 4907 15802
rect 4919 15750 4971 15802
rect 4983 15750 5035 15802
rect 5047 15750 5099 15802
rect 12473 15750 12525 15802
rect 12537 15750 12589 15802
rect 12601 15750 12653 15802
rect 12665 15750 12717 15802
rect 12729 15750 12781 15802
rect 20155 15750 20207 15802
rect 20219 15750 20271 15802
rect 20283 15750 20335 15802
rect 20347 15750 20399 15802
rect 20411 15750 20463 15802
rect 27837 15750 27889 15802
rect 27901 15750 27953 15802
rect 27965 15750 28017 15802
rect 28029 15750 28081 15802
rect 28093 15750 28145 15802
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 11796 15691 11848 15700
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 14924 15648 14976 15700
rect 15108 15648 15160 15700
rect 15844 15648 15896 15700
rect 15936 15648 15988 15700
rect 16304 15648 16356 15700
rect 16488 15691 16540 15700
rect 16488 15657 16497 15691
rect 16497 15657 16531 15691
rect 16531 15657 16540 15691
rect 16488 15648 16540 15657
rect 11244 15580 11296 15632
rect 15568 15580 15620 15632
rect 13084 15512 13136 15564
rect 16120 15580 16172 15632
rect 17040 15648 17092 15700
rect 17592 15580 17644 15632
rect 18972 15648 19024 15700
rect 19156 15580 19208 15632
rect 19432 15580 19484 15632
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 11796 15444 11848 15496
rect 13268 15444 13320 15496
rect 15936 15512 15988 15564
rect 16948 15512 17000 15564
rect 19064 15512 19116 15564
rect 20076 15512 20128 15564
rect 20904 15648 20956 15700
rect 21456 15648 21508 15700
rect 24676 15648 24728 15700
rect 25964 15648 26016 15700
rect 27068 15648 27120 15700
rect 27896 15691 27948 15700
rect 27896 15657 27905 15691
rect 27905 15657 27939 15691
rect 27939 15657 27948 15691
rect 27896 15648 27948 15657
rect 23112 15580 23164 15632
rect 23572 15580 23624 15632
rect 27436 15580 27488 15632
rect 28816 15648 28868 15700
rect 29000 15648 29052 15700
rect 28264 15580 28316 15632
rect 29092 15580 29144 15632
rect 30196 15580 30248 15632
rect 10876 15376 10928 15428
rect 13084 15376 13136 15428
rect 15016 15444 15068 15496
rect 16212 15444 16264 15496
rect 16580 15444 16632 15496
rect 15660 15419 15712 15428
rect 12992 15351 13044 15360
rect 12992 15317 13001 15351
rect 13001 15317 13035 15351
rect 13035 15317 13044 15351
rect 12992 15308 13044 15317
rect 15660 15385 15669 15419
rect 15669 15385 15703 15419
rect 15703 15385 15712 15419
rect 15660 15376 15712 15385
rect 16488 15376 16540 15428
rect 15568 15308 15620 15360
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 17592 15376 17644 15428
rect 17868 15308 17920 15360
rect 18696 15376 18748 15428
rect 19616 15376 19668 15428
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 20720 15376 20772 15428
rect 23756 15444 23808 15496
rect 24492 15444 24544 15496
rect 26792 15512 26844 15564
rect 26884 15444 26936 15496
rect 27528 15512 27580 15564
rect 28264 15444 28316 15496
rect 28632 15512 28684 15564
rect 29460 15444 29512 15496
rect 22008 15376 22060 15428
rect 22192 15376 22244 15428
rect 18880 15308 18932 15360
rect 19432 15308 19484 15360
rect 27804 15376 27856 15428
rect 28356 15376 28408 15428
rect 30472 15376 30524 15428
rect 30656 15419 30708 15428
rect 30656 15385 30665 15419
rect 30665 15385 30699 15419
rect 30699 15385 30708 15419
rect 30656 15376 30708 15385
rect 26148 15308 26200 15360
rect 26332 15351 26384 15360
rect 26332 15317 26341 15351
rect 26341 15317 26375 15351
rect 26375 15317 26384 15351
rect 26332 15308 26384 15317
rect 26792 15351 26844 15360
rect 26792 15317 26801 15351
rect 26801 15317 26835 15351
rect 26835 15317 26844 15351
rect 26792 15308 26844 15317
rect 28448 15308 28500 15360
rect 28632 15308 28684 15360
rect 29184 15308 29236 15360
rect 29920 15308 29972 15360
rect 31668 15308 31720 15360
rect 8632 15206 8684 15258
rect 8696 15206 8748 15258
rect 8760 15206 8812 15258
rect 8824 15206 8876 15258
rect 8888 15206 8940 15258
rect 16314 15206 16366 15258
rect 16378 15206 16430 15258
rect 16442 15206 16494 15258
rect 16506 15206 16558 15258
rect 16570 15206 16622 15258
rect 23996 15206 24048 15258
rect 24060 15206 24112 15258
rect 24124 15206 24176 15258
rect 24188 15206 24240 15258
rect 24252 15206 24304 15258
rect 31678 15206 31730 15258
rect 31742 15206 31794 15258
rect 31806 15206 31858 15258
rect 31870 15206 31922 15258
rect 31934 15206 31986 15258
rect 11336 15104 11388 15156
rect 12164 15104 12216 15156
rect 12348 15036 12400 15088
rect 13912 15036 13964 15088
rect 14740 15104 14792 15156
rect 15200 15104 15252 15156
rect 15384 15104 15436 15156
rect 17500 15104 17552 15156
rect 18328 15104 18380 15156
rect 15108 15079 15160 15088
rect 15108 15045 15117 15079
rect 15117 15045 15151 15079
rect 15151 15045 15160 15079
rect 15108 15036 15160 15045
rect 15660 15036 15712 15088
rect 19800 15036 19852 15088
rect 15292 15011 15344 15020
rect 15292 14977 15301 15011
rect 15301 14977 15335 15011
rect 15335 14977 15344 15011
rect 15292 14968 15344 14977
rect 15384 15011 15436 15020
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 15568 14968 15620 15020
rect 17408 14968 17460 15020
rect 17868 14968 17920 15020
rect 18604 14968 18656 15020
rect 14924 14832 14976 14884
rect 15200 14832 15252 14884
rect 16120 14900 16172 14952
rect 16304 14943 16356 14952
rect 16304 14909 16313 14943
rect 16313 14909 16347 14943
rect 16347 14909 16356 14943
rect 16304 14900 16356 14909
rect 16488 14900 16540 14952
rect 17684 14943 17736 14952
rect 17316 14832 17368 14884
rect 17684 14909 17693 14943
rect 17693 14909 17727 14943
rect 17727 14909 17736 14943
rect 17684 14900 17736 14909
rect 18788 14832 18840 14884
rect 14004 14807 14056 14816
rect 14004 14773 14013 14807
rect 14013 14773 14047 14807
rect 14047 14773 14056 14807
rect 14004 14764 14056 14773
rect 14648 14764 14700 14816
rect 15844 14764 15896 14816
rect 16488 14764 16540 14816
rect 16672 14764 16724 14816
rect 17776 14764 17828 14816
rect 19524 14900 19576 14952
rect 21732 15104 21784 15156
rect 22836 15104 22888 15156
rect 24768 15104 24820 15156
rect 28632 15104 28684 15156
rect 28816 15104 28868 15156
rect 30012 15104 30064 15156
rect 30104 15104 30156 15156
rect 30564 15104 30616 15156
rect 23388 15036 23440 15088
rect 24584 15036 24636 15088
rect 25228 15036 25280 15088
rect 25964 15036 26016 15088
rect 26240 15036 26292 15088
rect 27804 15036 27856 15088
rect 30196 15036 30248 15088
rect 30472 15036 30524 15088
rect 21456 14943 21508 14952
rect 21456 14909 21465 14943
rect 21465 14909 21499 14943
rect 21499 14909 21508 14943
rect 21456 14900 21508 14909
rect 21548 14900 21600 14952
rect 22744 14900 22796 14952
rect 20812 14832 20864 14884
rect 22376 14832 22428 14884
rect 24584 14900 24636 14952
rect 25504 14900 25556 14952
rect 25688 14900 25740 14952
rect 25964 14900 26016 14952
rect 27712 14968 27764 15020
rect 27988 14968 28040 15020
rect 27896 14900 27948 14952
rect 28632 14968 28684 15020
rect 29644 15011 29696 15020
rect 29644 14977 29653 15011
rect 29653 14977 29687 15011
rect 29687 14977 29696 15011
rect 29644 14968 29696 14977
rect 29736 14968 29788 15020
rect 32404 14968 32456 15020
rect 28448 14900 28500 14952
rect 19708 14764 19760 14816
rect 20076 14764 20128 14816
rect 21732 14764 21784 14816
rect 22008 14764 22060 14816
rect 22284 14764 22336 14816
rect 23664 14764 23716 14816
rect 26884 14832 26936 14884
rect 28632 14832 28684 14884
rect 24492 14764 24544 14816
rect 26056 14764 26108 14816
rect 27620 14764 27672 14816
rect 28172 14764 28224 14816
rect 29184 14832 29236 14884
rect 30012 14900 30064 14952
rect 29092 14764 29144 14816
rect 29920 14764 29972 14816
rect 30012 14764 30064 14816
rect 4791 14662 4843 14714
rect 4855 14662 4907 14714
rect 4919 14662 4971 14714
rect 4983 14662 5035 14714
rect 5047 14662 5099 14714
rect 12473 14662 12525 14714
rect 12537 14662 12589 14714
rect 12601 14662 12653 14714
rect 12665 14662 12717 14714
rect 12729 14662 12781 14714
rect 20155 14662 20207 14714
rect 20219 14662 20271 14714
rect 20283 14662 20335 14714
rect 20347 14662 20399 14714
rect 20411 14662 20463 14714
rect 27837 14662 27889 14714
rect 27901 14662 27953 14714
rect 27965 14662 28017 14714
rect 28029 14662 28081 14714
rect 28093 14662 28145 14714
rect 10968 14560 11020 14612
rect 12164 14492 12216 14544
rect 14372 14492 14424 14544
rect 15476 14560 15528 14612
rect 17040 14560 17092 14612
rect 17316 14603 17368 14612
rect 17316 14569 17325 14603
rect 17325 14569 17359 14603
rect 17359 14569 17368 14603
rect 17316 14560 17368 14569
rect 16948 14492 17000 14544
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 13728 14424 13780 14476
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 16304 14424 16356 14476
rect 18052 14560 18104 14612
rect 18236 14560 18288 14612
rect 20444 14560 20496 14612
rect 18604 14492 18656 14544
rect 18880 14535 18932 14544
rect 18880 14501 18889 14535
rect 18889 14501 18923 14535
rect 18923 14501 18932 14535
rect 18880 14492 18932 14501
rect 19248 14492 19300 14544
rect 21180 14560 21232 14612
rect 21456 14560 21508 14612
rect 25412 14560 25464 14612
rect 26792 14603 26844 14612
rect 22376 14492 22428 14544
rect 25504 14492 25556 14544
rect 26792 14569 26801 14603
rect 26801 14569 26835 14603
rect 26835 14569 26844 14603
rect 26792 14560 26844 14569
rect 27160 14560 27212 14612
rect 30472 14603 30524 14612
rect 30472 14569 30481 14603
rect 30481 14569 30515 14603
rect 30515 14569 30524 14603
rect 30472 14560 30524 14569
rect 31392 14560 31444 14612
rect 26884 14492 26936 14544
rect 27804 14492 27856 14544
rect 27896 14492 27948 14544
rect 28448 14492 28500 14544
rect 14372 14288 14424 14340
rect 16120 14356 16172 14408
rect 17868 14424 17920 14476
rect 18052 14424 18104 14476
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 16764 14356 16816 14408
rect 16948 14356 17000 14408
rect 17040 14356 17092 14408
rect 17316 14356 17368 14408
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 18236 14356 18288 14408
rect 15568 14288 15620 14340
rect 15844 14288 15896 14340
rect 16304 14288 16356 14340
rect 17132 14288 17184 14340
rect 19616 14424 19668 14476
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 13360 14220 13412 14272
rect 16764 14220 16816 14272
rect 19156 14220 19208 14272
rect 19708 14220 19760 14272
rect 21364 14424 21416 14476
rect 23020 14424 23072 14476
rect 24768 14424 24820 14476
rect 26976 14424 27028 14476
rect 22744 14356 22796 14408
rect 21456 14288 21508 14340
rect 22836 14288 22888 14340
rect 26056 14356 26108 14408
rect 27436 14399 27488 14408
rect 27436 14365 27445 14399
rect 27445 14365 27479 14399
rect 27479 14365 27488 14399
rect 27436 14356 27488 14365
rect 28632 14424 28684 14476
rect 29000 14399 29052 14408
rect 20352 14220 20404 14272
rect 21088 14220 21140 14272
rect 21180 14220 21232 14272
rect 22008 14220 22060 14272
rect 23480 14220 23532 14272
rect 24124 14288 24176 14340
rect 25044 14288 25096 14340
rect 26792 14331 26844 14340
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 25688 14220 25740 14272
rect 26056 14220 26108 14272
rect 26792 14297 26819 14331
rect 26819 14297 26844 14331
rect 26792 14288 26844 14297
rect 26884 14288 26936 14340
rect 27988 14220 28040 14272
rect 28448 14288 28500 14340
rect 29000 14365 29009 14399
rect 29009 14365 29043 14399
rect 29043 14365 29052 14399
rect 29000 14356 29052 14365
rect 29644 14356 29696 14408
rect 29828 14356 29880 14408
rect 30564 14356 30616 14408
rect 31024 14356 31076 14408
rect 29276 14288 29328 14340
rect 28816 14220 28868 14272
rect 29828 14263 29880 14272
rect 29828 14229 29837 14263
rect 29837 14229 29871 14263
rect 29871 14229 29880 14263
rect 29828 14220 29880 14229
rect 8632 14118 8684 14170
rect 8696 14118 8748 14170
rect 8760 14118 8812 14170
rect 8824 14118 8876 14170
rect 8888 14118 8940 14170
rect 16314 14118 16366 14170
rect 16378 14118 16430 14170
rect 16442 14118 16494 14170
rect 16506 14118 16558 14170
rect 16570 14118 16622 14170
rect 23996 14118 24048 14170
rect 24060 14118 24112 14170
rect 24124 14118 24176 14170
rect 24188 14118 24240 14170
rect 24252 14118 24304 14170
rect 31678 14118 31730 14170
rect 31742 14118 31794 14170
rect 31806 14118 31858 14170
rect 31870 14118 31922 14170
rect 31934 14118 31986 14170
rect 13084 14016 13136 14068
rect 13360 14016 13412 14068
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 14096 14016 14148 14068
rect 14372 13991 14424 14000
rect 14372 13957 14381 13991
rect 14381 13957 14415 13991
rect 14415 13957 14424 13991
rect 14372 13948 14424 13957
rect 15200 13948 15252 14000
rect 14464 13880 14516 13932
rect 15660 13923 15712 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 14740 13812 14792 13864
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 16396 13880 16448 13932
rect 16764 14016 16816 14068
rect 18236 14016 18288 14068
rect 22008 14016 22060 14068
rect 23664 14016 23716 14068
rect 23848 14016 23900 14068
rect 27620 14016 27672 14068
rect 28632 14016 28684 14068
rect 28724 14016 28776 14068
rect 30012 14016 30064 14068
rect 17224 13991 17276 14000
rect 17224 13957 17233 13991
rect 17233 13957 17267 13991
rect 17267 13957 17276 13991
rect 17224 13948 17276 13957
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17408 13923 17460 13932
rect 17132 13880 17184 13889
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 17868 13880 17920 13932
rect 18052 13923 18104 13932
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 16672 13812 16724 13864
rect 16764 13812 16816 13864
rect 14004 13744 14056 13796
rect 18328 13812 18380 13864
rect 19432 13948 19484 14000
rect 19616 13948 19668 14000
rect 20536 13948 20588 14000
rect 21732 13948 21784 14000
rect 18696 13880 18748 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 20444 13812 20496 13864
rect 21732 13812 21784 13864
rect 23848 13880 23900 13932
rect 24400 13880 24452 13932
rect 24768 13880 24820 13932
rect 23664 13812 23716 13864
rect 26424 13948 26476 14000
rect 25412 13880 25464 13932
rect 25504 13880 25556 13932
rect 26148 13880 26200 13932
rect 26700 13880 26752 13932
rect 29000 13948 29052 14000
rect 26884 13880 26936 13932
rect 27804 13923 27856 13932
rect 27252 13855 27304 13864
rect 20812 13744 20864 13796
rect 20996 13744 21048 13796
rect 23388 13744 23440 13796
rect 24768 13744 24820 13796
rect 25044 13744 25096 13796
rect 15384 13676 15436 13728
rect 18420 13676 18472 13728
rect 19156 13676 19208 13728
rect 21364 13676 21416 13728
rect 24216 13676 24268 13728
rect 25412 13719 25464 13728
rect 25412 13685 25421 13719
rect 25421 13685 25455 13719
rect 25455 13685 25464 13719
rect 25412 13676 25464 13685
rect 27252 13821 27261 13855
rect 27261 13821 27295 13855
rect 27295 13821 27304 13855
rect 27252 13812 27304 13821
rect 26240 13744 26292 13796
rect 26792 13744 26844 13796
rect 27804 13889 27813 13923
rect 27813 13889 27847 13923
rect 27847 13889 27856 13923
rect 27804 13880 27856 13889
rect 28080 13880 28132 13932
rect 28448 13923 28500 13932
rect 28448 13889 28457 13923
rect 28457 13889 28491 13923
rect 28491 13889 28500 13923
rect 28448 13880 28500 13889
rect 27988 13744 28040 13796
rect 28908 13880 28960 13932
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 29736 13880 29788 13932
rect 30840 13880 30892 13932
rect 31484 13880 31536 13932
rect 25688 13676 25740 13728
rect 25964 13676 26016 13728
rect 27896 13676 27948 13728
rect 29000 13676 29052 13728
rect 29184 13719 29236 13728
rect 29184 13685 29193 13719
rect 29193 13685 29227 13719
rect 29227 13685 29236 13719
rect 29184 13676 29236 13685
rect 4791 13574 4843 13626
rect 4855 13574 4907 13626
rect 4919 13574 4971 13626
rect 4983 13574 5035 13626
rect 5047 13574 5099 13626
rect 12473 13574 12525 13626
rect 12537 13574 12589 13626
rect 12601 13574 12653 13626
rect 12665 13574 12717 13626
rect 12729 13574 12781 13626
rect 20155 13574 20207 13626
rect 20219 13574 20271 13626
rect 20283 13574 20335 13626
rect 20347 13574 20399 13626
rect 20411 13574 20463 13626
rect 27837 13574 27889 13626
rect 27901 13574 27953 13626
rect 27965 13574 28017 13626
rect 28029 13574 28081 13626
rect 28093 13574 28145 13626
rect 15200 13515 15252 13524
rect 15200 13481 15209 13515
rect 15209 13481 15243 13515
rect 15243 13481 15252 13515
rect 15200 13472 15252 13481
rect 15292 13472 15344 13524
rect 16304 13472 16356 13524
rect 14832 13404 14884 13456
rect 16948 13404 17000 13456
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 16028 13336 16080 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 19248 13472 19300 13524
rect 19340 13472 19392 13524
rect 18788 13404 18840 13456
rect 19616 13404 19668 13456
rect 26976 13472 27028 13524
rect 27344 13515 27396 13524
rect 27344 13481 27353 13515
rect 27353 13481 27387 13515
rect 27387 13481 27396 13515
rect 27344 13472 27396 13481
rect 28172 13472 28224 13524
rect 28540 13515 28592 13524
rect 28540 13481 28549 13515
rect 28549 13481 28583 13515
rect 28583 13481 28592 13515
rect 28540 13472 28592 13481
rect 30012 13515 30064 13524
rect 30012 13481 30021 13515
rect 30021 13481 30055 13515
rect 30055 13481 30064 13515
rect 30012 13472 30064 13481
rect 30656 13472 30708 13524
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 16212 13268 16264 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 18512 13311 18564 13320
rect 16948 13200 17000 13252
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18696 13268 18748 13320
rect 21364 13336 21416 13388
rect 22008 13336 22060 13388
rect 24216 13336 24268 13388
rect 24860 13336 24912 13388
rect 27712 13404 27764 13456
rect 19800 13268 19852 13320
rect 24032 13311 24084 13320
rect 14280 13132 14332 13184
rect 18880 13132 18932 13184
rect 19616 13132 19668 13184
rect 20996 13200 21048 13252
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 25964 13311 26016 13320
rect 21364 13200 21416 13252
rect 22652 13200 22704 13252
rect 25504 13200 25556 13252
rect 25964 13277 25973 13311
rect 25973 13277 26007 13311
rect 26007 13277 26016 13311
rect 25964 13268 26016 13277
rect 30748 13336 30800 13388
rect 27436 13268 27488 13320
rect 27528 13268 27580 13320
rect 29276 13268 29328 13320
rect 31208 13268 31260 13320
rect 26148 13200 26200 13252
rect 27620 13200 27672 13252
rect 22284 13132 22336 13184
rect 25412 13132 25464 13184
rect 28264 13132 28316 13184
rect 28908 13132 28960 13184
rect 8632 13030 8684 13082
rect 8696 13030 8748 13082
rect 8760 13030 8812 13082
rect 8824 13030 8876 13082
rect 8888 13030 8940 13082
rect 16314 13030 16366 13082
rect 16378 13030 16430 13082
rect 16442 13030 16494 13082
rect 16506 13030 16558 13082
rect 16570 13030 16622 13082
rect 23996 13030 24048 13082
rect 24060 13030 24112 13082
rect 24124 13030 24176 13082
rect 24188 13030 24240 13082
rect 24252 13030 24304 13082
rect 31678 13030 31730 13082
rect 31742 13030 31794 13082
rect 31806 13030 31858 13082
rect 31870 13030 31922 13082
rect 31934 13030 31986 13082
rect 15844 12928 15896 12980
rect 16212 12903 16264 12912
rect 16212 12869 16221 12903
rect 16221 12869 16255 12903
rect 16255 12869 16264 12903
rect 16212 12860 16264 12869
rect 18144 12860 18196 12912
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 18236 12835 18288 12844
rect 18236 12801 18245 12835
rect 18245 12801 18279 12835
rect 18279 12801 18288 12835
rect 18236 12792 18288 12801
rect 18420 12860 18472 12912
rect 19156 12860 19208 12912
rect 19248 12903 19300 12912
rect 19248 12869 19257 12903
rect 19257 12869 19291 12903
rect 19291 12869 19300 12903
rect 19248 12860 19300 12869
rect 18512 12792 18564 12844
rect 18788 12724 18840 12776
rect 16672 12656 16724 12708
rect 17960 12588 18012 12640
rect 19524 12656 19576 12708
rect 19064 12631 19116 12640
rect 19064 12597 19073 12631
rect 19073 12597 19107 12631
rect 19107 12597 19116 12631
rect 19064 12588 19116 12597
rect 19340 12588 19392 12640
rect 20996 12860 21048 12912
rect 23848 12928 23900 12980
rect 25688 12928 25740 12980
rect 25872 12928 25924 12980
rect 27160 12928 27212 12980
rect 27344 12928 27396 12980
rect 29828 12860 29880 12912
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 24860 12792 24912 12844
rect 25044 12835 25096 12844
rect 25044 12801 25053 12835
rect 25053 12801 25087 12835
rect 25087 12801 25096 12835
rect 25044 12792 25096 12801
rect 25412 12792 25464 12844
rect 26240 12792 26292 12844
rect 26792 12792 26844 12844
rect 26976 12792 27028 12844
rect 27528 12792 27580 12844
rect 31300 12835 31352 12844
rect 31300 12801 31309 12835
rect 31309 12801 31343 12835
rect 31343 12801 31352 12835
rect 31300 12792 31352 12801
rect 20628 12724 20680 12776
rect 20720 12724 20772 12776
rect 23020 12724 23072 12776
rect 24768 12724 24820 12776
rect 24400 12656 24452 12708
rect 26608 12724 26660 12776
rect 27068 12724 27120 12776
rect 28356 12656 28408 12708
rect 28540 12656 28592 12708
rect 29736 12656 29788 12708
rect 19984 12588 20036 12640
rect 24768 12588 24820 12640
rect 25320 12588 25372 12640
rect 28632 12588 28684 12640
rect 29368 12588 29420 12640
rect 4791 12486 4843 12538
rect 4855 12486 4907 12538
rect 4919 12486 4971 12538
rect 4983 12486 5035 12538
rect 5047 12486 5099 12538
rect 12473 12486 12525 12538
rect 12537 12486 12589 12538
rect 12601 12486 12653 12538
rect 12665 12486 12717 12538
rect 12729 12486 12781 12538
rect 20155 12486 20207 12538
rect 20219 12486 20271 12538
rect 20283 12486 20335 12538
rect 20347 12486 20399 12538
rect 20411 12486 20463 12538
rect 27837 12486 27889 12538
rect 27901 12486 27953 12538
rect 27965 12486 28017 12538
rect 28029 12486 28081 12538
rect 28093 12486 28145 12538
rect 16212 12384 16264 12436
rect 17040 12384 17092 12436
rect 17684 12384 17736 12436
rect 19892 12384 19944 12436
rect 13728 12316 13780 12368
rect 18880 12316 18932 12368
rect 23572 12384 23624 12436
rect 24400 12384 24452 12436
rect 24676 12427 24728 12436
rect 24676 12393 24685 12427
rect 24685 12393 24719 12427
rect 24719 12393 24728 12427
rect 24676 12384 24728 12393
rect 24860 12384 24912 12436
rect 22284 12316 22336 12368
rect 22744 12316 22796 12368
rect 24952 12316 25004 12368
rect 25136 12384 25188 12436
rect 26976 12384 27028 12436
rect 28172 12384 28224 12436
rect 28448 12384 28500 12436
rect 31300 12427 31352 12436
rect 31300 12393 31309 12427
rect 31309 12393 31343 12427
rect 31343 12393 31352 12427
rect 31300 12384 31352 12393
rect 25320 12316 25372 12368
rect 25872 12316 25924 12368
rect 26700 12316 26752 12368
rect 28080 12316 28132 12368
rect 28816 12316 28868 12368
rect 13544 12248 13596 12300
rect 17408 12248 17460 12300
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 14924 12112 14976 12164
rect 18972 12248 19024 12300
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 18328 12180 18380 12232
rect 18420 12180 18472 12232
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 20076 12180 20128 12232
rect 20628 12223 20680 12232
rect 20628 12189 20637 12223
rect 20637 12189 20671 12223
rect 20671 12189 20680 12223
rect 20628 12180 20680 12189
rect 22744 12180 22796 12232
rect 23020 12180 23072 12232
rect 23388 12180 23440 12232
rect 22468 12112 22520 12164
rect 23664 12180 23716 12232
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 24860 12180 24912 12232
rect 27252 12248 27304 12300
rect 28356 12248 28408 12300
rect 29276 12248 29328 12300
rect 26056 12180 26108 12232
rect 26332 12180 26384 12232
rect 26884 12180 26936 12232
rect 28724 12180 28776 12232
rect 30472 12180 30524 12232
rect 17316 12044 17368 12096
rect 17684 12044 17736 12096
rect 18236 12044 18288 12096
rect 19892 12044 19944 12096
rect 21732 12044 21784 12096
rect 22376 12087 22428 12096
rect 22376 12053 22385 12087
rect 22385 12053 22419 12087
rect 22419 12053 22428 12087
rect 22376 12044 22428 12053
rect 24584 12044 24636 12096
rect 24952 12044 25004 12096
rect 25504 12112 25556 12164
rect 29368 12112 29420 12164
rect 27160 12087 27212 12096
rect 27160 12053 27169 12087
rect 27169 12053 27203 12087
rect 27203 12053 27212 12087
rect 27160 12044 27212 12053
rect 27988 12044 28040 12096
rect 28816 12087 28868 12096
rect 28816 12053 28825 12087
rect 28825 12053 28859 12087
rect 28859 12053 28868 12087
rect 28816 12044 28868 12053
rect 30196 12044 30248 12096
rect 30656 12044 30708 12096
rect 8632 11942 8684 11994
rect 8696 11942 8748 11994
rect 8760 11942 8812 11994
rect 8824 11942 8876 11994
rect 8888 11942 8940 11994
rect 16314 11942 16366 11994
rect 16378 11942 16430 11994
rect 16442 11942 16494 11994
rect 16506 11942 16558 11994
rect 16570 11942 16622 11994
rect 23996 11942 24048 11994
rect 24060 11942 24112 11994
rect 24124 11942 24176 11994
rect 24188 11942 24240 11994
rect 24252 11942 24304 11994
rect 31678 11942 31730 11994
rect 31742 11942 31794 11994
rect 31806 11942 31858 11994
rect 31870 11942 31922 11994
rect 31934 11942 31986 11994
rect 9588 11840 9640 11892
rect 17776 11840 17828 11892
rect 17040 11772 17092 11824
rect 18328 11840 18380 11892
rect 19524 11883 19576 11892
rect 19524 11849 19533 11883
rect 19533 11849 19567 11883
rect 19567 11849 19576 11883
rect 19524 11840 19576 11849
rect 22008 11883 22060 11892
rect 17960 11772 18012 11824
rect 15936 11704 15988 11756
rect 18236 11704 18288 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 17592 11636 17644 11688
rect 19892 11636 19944 11688
rect 16948 11568 17000 11620
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 22744 11840 22796 11892
rect 22928 11883 22980 11892
rect 22928 11849 22937 11883
rect 22937 11849 22971 11883
rect 22971 11849 22980 11883
rect 22928 11840 22980 11849
rect 23572 11883 23624 11892
rect 23572 11849 23581 11883
rect 23581 11849 23615 11883
rect 23615 11849 23624 11883
rect 23572 11840 23624 11849
rect 23848 11840 23900 11892
rect 25136 11840 25188 11892
rect 26148 11840 26200 11892
rect 22376 11815 22428 11824
rect 20904 11704 20956 11756
rect 20720 11636 20772 11688
rect 21272 11704 21324 11756
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 22376 11781 22385 11815
rect 22385 11781 22419 11815
rect 22419 11781 22428 11815
rect 22376 11772 22428 11781
rect 28080 11840 28132 11892
rect 28264 11840 28316 11892
rect 21916 11704 21968 11756
rect 23572 11704 23624 11756
rect 23848 11704 23900 11756
rect 24768 11704 24820 11756
rect 24860 11704 24912 11756
rect 25044 11704 25096 11756
rect 25872 11704 25924 11756
rect 26332 11747 26384 11756
rect 26332 11713 26341 11747
rect 26341 11713 26375 11747
rect 26375 11713 26384 11747
rect 27528 11772 27580 11824
rect 27620 11772 27672 11824
rect 30472 11772 30524 11824
rect 31300 11747 31352 11756
rect 26332 11704 26384 11713
rect 31300 11713 31309 11747
rect 31309 11713 31343 11747
rect 31343 11713 31352 11747
rect 31300 11704 31352 11713
rect 21180 11636 21232 11645
rect 22100 11568 22152 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 15108 11500 15160 11552
rect 17316 11500 17368 11552
rect 17408 11500 17460 11552
rect 20720 11500 20772 11552
rect 21088 11500 21140 11552
rect 24584 11568 24636 11620
rect 29460 11636 29512 11688
rect 26792 11568 26844 11620
rect 27988 11568 28040 11620
rect 23388 11500 23440 11552
rect 27712 11543 27764 11552
rect 27712 11509 27721 11543
rect 27721 11509 27755 11543
rect 27755 11509 27764 11543
rect 27712 11500 27764 11509
rect 29368 11543 29420 11552
rect 29368 11509 29377 11543
rect 29377 11509 29411 11543
rect 29411 11509 29420 11543
rect 29368 11500 29420 11509
rect 30380 11500 30432 11552
rect 4791 11398 4843 11450
rect 4855 11398 4907 11450
rect 4919 11398 4971 11450
rect 4983 11398 5035 11450
rect 5047 11398 5099 11450
rect 12473 11398 12525 11450
rect 12537 11398 12589 11450
rect 12601 11398 12653 11450
rect 12665 11398 12717 11450
rect 12729 11398 12781 11450
rect 20155 11398 20207 11450
rect 20219 11398 20271 11450
rect 20283 11398 20335 11450
rect 20347 11398 20399 11450
rect 20411 11398 20463 11450
rect 27837 11398 27889 11450
rect 27901 11398 27953 11450
rect 27965 11398 28017 11450
rect 28029 11398 28081 11450
rect 28093 11398 28145 11450
rect 16120 11296 16172 11348
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 22192 11339 22244 11348
rect 22192 11305 22201 11339
rect 22201 11305 22235 11339
rect 22235 11305 22244 11339
rect 22192 11296 22244 11305
rect 23296 11296 23348 11348
rect 23480 11339 23532 11348
rect 23480 11305 23489 11339
rect 23489 11305 23523 11339
rect 23523 11305 23532 11339
rect 23480 11296 23532 11305
rect 26608 11296 26660 11348
rect 26884 11296 26936 11348
rect 27988 11296 28040 11348
rect 29644 11296 29696 11348
rect 31300 11339 31352 11348
rect 31300 11305 31309 11339
rect 31309 11305 31343 11339
rect 31343 11305 31352 11339
rect 31300 11296 31352 11305
rect 21824 11228 21876 11280
rect 22008 11228 22060 11280
rect 28172 11228 28224 11280
rect 17316 11160 17368 11212
rect 19248 11160 19300 11212
rect 19892 11092 19944 11144
rect 20904 11160 20956 11212
rect 24584 11160 24636 11212
rect 27620 11160 27672 11212
rect 20812 11135 20864 11144
rect 20812 11101 20821 11135
rect 20821 11101 20855 11135
rect 20855 11101 20864 11135
rect 21456 11135 21508 11144
rect 20812 11092 20864 11101
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 22008 11092 22060 11144
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 28264 11092 28316 11144
rect 13452 11024 13504 11076
rect 20904 11024 20956 11076
rect 4160 10956 4212 11008
rect 9496 10956 9548 11008
rect 19156 10956 19208 11008
rect 20076 10956 20128 11008
rect 22836 11024 22888 11076
rect 24676 11067 24728 11076
rect 24676 11033 24685 11067
rect 24685 11033 24719 11067
rect 24719 11033 24728 11067
rect 24676 11024 24728 11033
rect 27528 11024 27580 11076
rect 27988 11024 28040 11076
rect 21088 10956 21140 11008
rect 25504 10956 25556 11008
rect 25780 10956 25832 11008
rect 26332 10999 26384 11008
rect 26332 10965 26341 10999
rect 26341 10965 26375 10999
rect 26375 10965 26384 10999
rect 26332 10956 26384 10965
rect 27068 10956 27120 11008
rect 27252 10956 27304 11008
rect 27712 10956 27764 11008
rect 28816 10956 28868 11008
rect 29736 10999 29788 11008
rect 29736 10965 29745 10999
rect 29745 10965 29779 10999
rect 29779 10965 29788 10999
rect 29736 10956 29788 10965
rect 8632 10854 8684 10906
rect 8696 10854 8748 10906
rect 8760 10854 8812 10906
rect 8824 10854 8876 10906
rect 8888 10854 8940 10906
rect 16314 10854 16366 10906
rect 16378 10854 16430 10906
rect 16442 10854 16494 10906
rect 16506 10854 16558 10906
rect 16570 10854 16622 10906
rect 23996 10854 24048 10906
rect 24060 10854 24112 10906
rect 24124 10854 24176 10906
rect 24188 10854 24240 10906
rect 24252 10854 24304 10906
rect 31678 10854 31730 10906
rect 31742 10854 31794 10906
rect 31806 10854 31858 10906
rect 31870 10854 31922 10906
rect 31934 10854 31986 10906
rect 19892 10752 19944 10804
rect 20536 10752 20588 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 22560 10752 22612 10804
rect 22652 10752 22704 10804
rect 23204 10752 23256 10804
rect 11520 10684 11572 10736
rect 22468 10684 22520 10736
rect 24676 10752 24728 10804
rect 31024 10795 31076 10804
rect 31024 10761 31033 10795
rect 31033 10761 31067 10795
rect 31067 10761 31076 10795
rect 31024 10752 31076 10761
rect 32588 10684 32640 10736
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 20720 10659 20772 10668
rect 1584 10591 1636 10600
rect 1584 10557 1593 10591
rect 1593 10557 1627 10591
rect 1627 10557 1636 10591
rect 1584 10548 1636 10557
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 20904 10659 20956 10668
rect 20904 10625 20913 10659
rect 20913 10625 20947 10659
rect 20947 10625 20956 10659
rect 20904 10616 20956 10625
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 23664 10616 23716 10668
rect 24584 10659 24636 10668
rect 24584 10625 24593 10659
rect 24593 10625 24627 10659
rect 24627 10625 24636 10659
rect 24584 10616 24636 10625
rect 25136 10616 25188 10668
rect 26332 10616 26384 10668
rect 29000 10548 29052 10600
rect 29920 10591 29972 10600
rect 29920 10557 29929 10591
rect 29929 10557 29963 10591
rect 29963 10557 29972 10591
rect 29920 10548 29972 10557
rect 5264 10480 5316 10532
rect 10324 10480 10376 10532
rect 20720 10480 20772 10532
rect 22192 10480 22244 10532
rect 22284 10480 22336 10532
rect 23204 10480 23256 10532
rect 17684 10412 17736 10464
rect 20812 10412 20864 10464
rect 21088 10412 21140 10464
rect 21548 10412 21600 10464
rect 24308 10412 24360 10464
rect 25136 10412 25188 10464
rect 26608 10412 26660 10464
rect 28356 10480 28408 10532
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 31392 10480 31444 10532
rect 27712 10412 27764 10421
rect 4791 10310 4843 10362
rect 4855 10310 4907 10362
rect 4919 10310 4971 10362
rect 4983 10310 5035 10362
rect 5047 10310 5099 10362
rect 12473 10310 12525 10362
rect 12537 10310 12589 10362
rect 12601 10310 12653 10362
rect 12665 10310 12717 10362
rect 12729 10310 12781 10362
rect 20155 10310 20207 10362
rect 20219 10310 20271 10362
rect 20283 10310 20335 10362
rect 20347 10310 20399 10362
rect 20411 10310 20463 10362
rect 27837 10310 27889 10362
rect 27901 10310 27953 10362
rect 27965 10310 28017 10362
rect 28029 10310 28081 10362
rect 28093 10310 28145 10362
rect 8116 10208 8168 10260
rect 20720 10208 20772 10260
rect 20996 10251 21048 10260
rect 20996 10217 21005 10251
rect 21005 10217 21039 10251
rect 21039 10217 21048 10251
rect 20996 10208 21048 10217
rect 22008 10208 22060 10260
rect 22652 10208 22704 10260
rect 23756 10251 23808 10260
rect 23756 10217 23765 10251
rect 23765 10217 23799 10251
rect 23799 10217 23808 10251
rect 23756 10208 23808 10217
rect 24400 10208 24452 10260
rect 25504 10251 25556 10260
rect 25504 10217 25513 10251
rect 25513 10217 25547 10251
rect 25547 10217 25556 10251
rect 25504 10208 25556 10217
rect 28264 10208 28316 10260
rect 30288 10251 30340 10260
rect 30288 10217 30297 10251
rect 30297 10217 30331 10251
rect 30331 10217 30340 10251
rect 30288 10208 30340 10217
rect 9312 10140 9364 10192
rect 22192 10140 22244 10192
rect 25228 10140 25280 10192
rect 20904 10072 20956 10124
rect 23112 10072 23164 10124
rect 23204 10072 23256 10124
rect 26792 10072 26844 10124
rect 13268 10004 13320 10056
rect 22100 10004 22152 10056
rect 23664 10004 23716 10056
rect 26976 10004 27028 10056
rect 31024 10004 31076 10056
rect 31300 10047 31352 10056
rect 31300 10013 31309 10047
rect 31309 10013 31343 10047
rect 31343 10013 31352 10047
rect 31300 10004 31352 10013
rect 4436 9936 4488 9988
rect 26424 9868 26476 9920
rect 26884 9936 26936 9988
rect 28448 9868 28500 9920
rect 29184 9868 29236 9920
rect 8632 9766 8684 9818
rect 8696 9766 8748 9818
rect 8760 9766 8812 9818
rect 8824 9766 8876 9818
rect 8888 9766 8940 9818
rect 16314 9766 16366 9818
rect 16378 9766 16430 9818
rect 16442 9766 16494 9818
rect 16506 9766 16558 9818
rect 16570 9766 16622 9818
rect 23996 9766 24048 9818
rect 24060 9766 24112 9818
rect 24124 9766 24176 9818
rect 24188 9766 24240 9818
rect 24252 9766 24304 9818
rect 31678 9766 31730 9818
rect 31742 9766 31794 9818
rect 31806 9766 31858 9818
rect 31870 9766 31922 9818
rect 31934 9766 31986 9818
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 21916 9664 21968 9716
rect 22100 9707 22152 9716
rect 22100 9673 22109 9707
rect 22109 9673 22143 9707
rect 22143 9673 22152 9707
rect 22652 9707 22704 9716
rect 22100 9664 22152 9673
rect 22652 9673 22661 9707
rect 22661 9673 22695 9707
rect 22695 9673 22704 9707
rect 23112 9707 23164 9716
rect 22652 9664 22704 9673
rect 23112 9673 23121 9707
rect 23121 9673 23155 9707
rect 23155 9673 23164 9707
rect 23112 9664 23164 9673
rect 25504 9664 25556 9716
rect 29644 9707 29696 9716
rect 29644 9673 29653 9707
rect 29653 9673 29687 9707
rect 29687 9673 29696 9707
rect 29644 9664 29696 9673
rect 12348 9596 12400 9648
rect 20628 9596 20680 9648
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 28908 9596 28960 9648
rect 6920 9528 6972 9580
rect 26608 9528 26660 9580
rect 28816 9528 28868 9580
rect 9128 9460 9180 9512
rect 24952 9460 25004 9512
rect 25228 9460 25280 9512
rect 26056 9460 26108 9512
rect 30196 9460 30248 9512
rect 10416 9392 10468 9444
rect 23756 9392 23808 9444
rect 7932 9324 7984 9376
rect 25596 9392 25648 9444
rect 32864 9392 32916 9444
rect 26424 9367 26476 9376
rect 26424 9333 26433 9367
rect 26433 9333 26467 9367
rect 26467 9333 26476 9367
rect 26424 9324 26476 9333
rect 30104 9367 30156 9376
rect 30104 9333 30113 9367
rect 30113 9333 30147 9367
rect 30147 9333 30156 9367
rect 30104 9324 30156 9333
rect 31300 9367 31352 9376
rect 31300 9333 31309 9367
rect 31309 9333 31343 9367
rect 31343 9333 31352 9367
rect 31300 9324 31352 9333
rect 4791 9222 4843 9274
rect 4855 9222 4907 9274
rect 4919 9222 4971 9274
rect 4983 9222 5035 9274
rect 5047 9222 5099 9274
rect 12473 9222 12525 9274
rect 12537 9222 12589 9274
rect 12601 9222 12653 9274
rect 12665 9222 12717 9274
rect 12729 9222 12781 9274
rect 20155 9222 20207 9274
rect 20219 9222 20271 9274
rect 20283 9222 20335 9274
rect 20347 9222 20399 9274
rect 20411 9222 20463 9274
rect 27837 9222 27889 9274
rect 27901 9222 27953 9274
rect 27965 9222 28017 9274
rect 28029 9222 28081 9274
rect 28093 9222 28145 9274
rect 6828 9120 6880 9172
rect 22928 9120 22980 9172
rect 23112 9163 23164 9172
rect 23112 9129 23121 9163
rect 23121 9129 23155 9163
rect 23155 9129 23164 9163
rect 23112 9120 23164 9129
rect 30196 9163 30248 9172
rect 30196 9129 30205 9163
rect 30205 9129 30239 9163
rect 30239 9129 30248 9163
rect 30196 9120 30248 9129
rect 25320 9052 25372 9104
rect 26148 9052 26200 9104
rect 27436 9052 27488 9104
rect 28172 9052 28224 9104
rect 9588 8984 9640 9036
rect 23848 8984 23900 9036
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 5448 8916 5500 8968
rect 20628 8916 20680 8968
rect 27712 8984 27764 9036
rect 28540 9027 28592 9036
rect 28540 8993 28549 9027
rect 28549 8993 28583 9027
rect 28583 8993 28592 9027
rect 28540 8984 28592 8993
rect 28356 8916 28408 8968
rect 29644 8916 29696 8968
rect 21916 8823 21968 8832
rect 21916 8789 21925 8823
rect 21925 8789 21959 8823
rect 21959 8789 21968 8823
rect 22560 8823 22612 8832
rect 21916 8780 21968 8789
rect 22560 8789 22569 8823
rect 22569 8789 22603 8823
rect 22603 8789 22612 8823
rect 22560 8780 22612 8789
rect 25228 8780 25280 8832
rect 29092 8823 29144 8832
rect 29092 8789 29101 8823
rect 29101 8789 29135 8823
rect 29135 8789 29144 8823
rect 29092 8780 29144 8789
rect 8632 8678 8684 8730
rect 8696 8678 8748 8730
rect 8760 8678 8812 8730
rect 8824 8678 8876 8730
rect 8888 8678 8940 8730
rect 16314 8678 16366 8730
rect 16378 8678 16430 8730
rect 16442 8678 16494 8730
rect 16506 8678 16558 8730
rect 16570 8678 16622 8730
rect 23996 8678 24048 8730
rect 24060 8678 24112 8730
rect 24124 8678 24176 8730
rect 24188 8678 24240 8730
rect 24252 8678 24304 8730
rect 31678 8678 31730 8730
rect 31742 8678 31794 8730
rect 31806 8678 31858 8730
rect 31870 8678 31922 8730
rect 31934 8678 31986 8730
rect 23112 8576 23164 8628
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 26240 8576 26292 8628
rect 27068 8576 27120 8628
rect 29184 8619 29236 8628
rect 29184 8585 29193 8619
rect 29193 8585 29227 8619
rect 29227 8585 29236 8619
rect 29184 8576 29236 8585
rect 29736 8619 29788 8628
rect 29736 8585 29745 8619
rect 29745 8585 29779 8619
rect 29779 8585 29788 8619
rect 29736 8576 29788 8585
rect 32036 8508 32088 8560
rect 22928 8440 22980 8492
rect 30748 8440 30800 8492
rect 14280 8372 14332 8424
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 1584 8304 1636 8313
rect 9496 8236 9548 8288
rect 21364 8236 21416 8288
rect 22560 8415 22612 8424
rect 22560 8381 22569 8415
rect 22569 8381 22603 8415
rect 22603 8381 22612 8415
rect 22560 8372 22612 8381
rect 28448 8372 28500 8424
rect 26240 8304 26292 8356
rect 28816 8304 28868 8356
rect 30380 8347 30432 8356
rect 30380 8313 30389 8347
rect 30389 8313 30423 8347
rect 30423 8313 30432 8347
rect 30380 8304 30432 8313
rect 31300 8347 31352 8356
rect 31300 8313 31309 8347
rect 31309 8313 31343 8347
rect 31343 8313 31352 8347
rect 31300 8304 31352 8313
rect 26056 8236 26108 8288
rect 4791 8134 4843 8186
rect 4855 8134 4907 8186
rect 4919 8134 4971 8186
rect 4983 8134 5035 8186
rect 5047 8134 5099 8186
rect 12473 8134 12525 8186
rect 12537 8134 12589 8186
rect 12601 8134 12653 8186
rect 12665 8134 12717 8186
rect 12729 8134 12781 8186
rect 20155 8134 20207 8186
rect 20219 8134 20271 8186
rect 20283 8134 20335 8186
rect 20347 8134 20399 8186
rect 20411 8134 20463 8186
rect 27837 8134 27889 8186
rect 27901 8134 27953 8186
rect 27965 8134 28017 8186
rect 28029 8134 28081 8186
rect 28093 8134 28145 8186
rect 10324 8032 10376 8084
rect 25228 8032 25280 8084
rect 25872 8075 25924 8084
rect 25872 8041 25881 8075
rect 25881 8041 25915 8075
rect 25915 8041 25924 8075
rect 25872 8032 25924 8041
rect 26792 8032 26844 8084
rect 27436 8032 27488 8084
rect 28356 8075 28408 8084
rect 28356 8041 28365 8075
rect 28365 8041 28399 8075
rect 28399 8041 28408 8075
rect 28356 8032 28408 8041
rect 28816 8075 28868 8084
rect 28816 8041 28825 8075
rect 28825 8041 28859 8075
rect 28859 8041 28868 8075
rect 29736 8075 29788 8084
rect 28816 8032 28868 8041
rect 29736 8041 29745 8075
rect 29745 8041 29779 8075
rect 29779 8041 29788 8075
rect 29736 8032 29788 8041
rect 30748 8032 30800 8084
rect 31392 8032 31444 8084
rect 32312 7964 32364 8016
rect 21364 7896 21416 7948
rect 7656 7828 7708 7880
rect 27252 7828 27304 7880
rect 27620 7896 27672 7948
rect 29184 7896 29236 7948
rect 30196 7896 30248 7948
rect 32772 7828 32824 7880
rect 9220 7692 9272 7744
rect 24860 7735 24912 7744
rect 24860 7701 24869 7735
rect 24869 7701 24903 7735
rect 24903 7701 24912 7735
rect 24860 7692 24912 7701
rect 28356 7760 28408 7812
rect 29092 7760 29144 7812
rect 26332 7692 26384 7744
rect 26700 7692 26752 7744
rect 8632 7590 8684 7642
rect 8696 7590 8748 7642
rect 8760 7590 8812 7642
rect 8824 7590 8876 7642
rect 8888 7590 8940 7642
rect 16314 7590 16366 7642
rect 16378 7590 16430 7642
rect 16442 7590 16494 7642
rect 16506 7590 16558 7642
rect 16570 7590 16622 7642
rect 23996 7590 24048 7642
rect 24060 7590 24112 7642
rect 24124 7590 24176 7642
rect 24188 7590 24240 7642
rect 24252 7590 24304 7642
rect 31678 7590 31730 7642
rect 31742 7590 31794 7642
rect 31806 7590 31858 7642
rect 31870 7590 31922 7642
rect 31934 7590 31986 7642
rect 25688 7488 25740 7540
rect 32128 7488 32180 7540
rect 26056 7463 26108 7472
rect 26056 7429 26065 7463
rect 26065 7429 26099 7463
rect 26099 7429 26108 7463
rect 26056 7420 26108 7429
rect 26608 7463 26660 7472
rect 26608 7429 26617 7463
rect 26617 7429 26651 7463
rect 26651 7429 26660 7463
rect 26608 7420 26660 7429
rect 27528 7420 27580 7472
rect 28540 7420 28592 7472
rect 30472 7463 30524 7472
rect 30472 7429 30481 7463
rect 30481 7429 30515 7463
rect 30515 7429 30524 7463
rect 30472 7420 30524 7429
rect 24860 7352 24912 7404
rect 26792 7352 26844 7404
rect 29920 7327 29972 7336
rect 29920 7293 29929 7327
rect 29929 7293 29963 7327
rect 29963 7293 29972 7327
rect 29920 7284 29972 7293
rect 30288 7284 30340 7336
rect 31300 7259 31352 7268
rect 31300 7225 31309 7259
rect 31309 7225 31343 7259
rect 31343 7225 31352 7259
rect 31300 7216 31352 7225
rect 24952 7191 25004 7200
rect 24952 7157 24961 7191
rect 24961 7157 24995 7191
rect 24995 7157 25004 7191
rect 24952 7148 25004 7157
rect 25688 7148 25740 7200
rect 4791 7046 4843 7098
rect 4855 7046 4907 7098
rect 4919 7046 4971 7098
rect 4983 7046 5035 7098
rect 5047 7046 5099 7098
rect 12473 7046 12525 7098
rect 12537 7046 12589 7098
rect 12601 7046 12653 7098
rect 12665 7046 12717 7098
rect 12729 7046 12781 7098
rect 20155 7046 20207 7098
rect 20219 7046 20271 7098
rect 20283 7046 20335 7098
rect 20347 7046 20399 7098
rect 20411 7046 20463 7098
rect 27837 7046 27889 7098
rect 27901 7046 27953 7098
rect 27965 7046 28017 7098
rect 28029 7046 28081 7098
rect 28093 7046 28145 7098
rect 25872 6876 25924 6928
rect 4252 6808 4304 6860
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 29460 6808 29512 6860
rect 31116 6808 31168 6860
rect 26424 6740 26476 6792
rect 29368 6740 29420 6792
rect 31024 6783 31076 6792
rect 31024 6749 31033 6783
rect 31033 6749 31067 6783
rect 31067 6749 31076 6783
rect 31024 6740 31076 6749
rect 27620 6672 27672 6724
rect 30472 6715 30524 6724
rect 30472 6681 30481 6715
rect 30481 6681 30515 6715
rect 30515 6681 30524 6715
rect 30472 6672 30524 6681
rect 25688 6647 25740 6656
rect 25688 6613 25697 6647
rect 25697 6613 25731 6647
rect 25731 6613 25740 6647
rect 25688 6604 25740 6613
rect 26240 6647 26292 6656
rect 26240 6613 26249 6647
rect 26249 6613 26283 6647
rect 26283 6613 26292 6647
rect 26240 6604 26292 6613
rect 26792 6647 26844 6656
rect 26792 6613 26801 6647
rect 26801 6613 26835 6647
rect 26835 6613 26844 6647
rect 26792 6604 26844 6613
rect 8632 6502 8684 6554
rect 8696 6502 8748 6554
rect 8760 6502 8812 6554
rect 8824 6502 8876 6554
rect 8888 6502 8940 6554
rect 16314 6502 16366 6554
rect 16378 6502 16430 6554
rect 16442 6502 16494 6554
rect 16506 6502 16558 6554
rect 16570 6502 16622 6554
rect 23996 6502 24048 6554
rect 24060 6502 24112 6554
rect 24124 6502 24176 6554
rect 24188 6502 24240 6554
rect 24252 6502 24304 6554
rect 31678 6502 31730 6554
rect 31742 6502 31794 6554
rect 31806 6502 31858 6554
rect 31870 6502 31922 6554
rect 31934 6502 31986 6554
rect 29736 6443 29788 6452
rect 29736 6409 29745 6443
rect 29745 6409 29779 6443
rect 29779 6409 29788 6443
rect 29736 6400 29788 6409
rect 25688 6196 25740 6248
rect 27620 6196 27672 6248
rect 28724 6239 28776 6248
rect 28724 6205 28733 6239
rect 28733 6205 28767 6239
rect 28767 6205 28776 6239
rect 28724 6196 28776 6205
rect 4528 6060 4580 6112
rect 29092 6128 29144 6180
rect 27712 6103 27764 6112
rect 27712 6069 27721 6103
rect 27721 6069 27755 6103
rect 27755 6069 27764 6103
rect 27712 6060 27764 6069
rect 31300 6103 31352 6112
rect 31300 6069 31309 6103
rect 31309 6069 31343 6103
rect 31343 6069 31352 6103
rect 31300 6060 31352 6069
rect 4791 5958 4843 6010
rect 4855 5958 4907 6010
rect 4919 5958 4971 6010
rect 4983 5958 5035 6010
rect 5047 5958 5099 6010
rect 12473 5958 12525 6010
rect 12537 5958 12589 6010
rect 12601 5958 12653 6010
rect 12665 5958 12717 6010
rect 12729 5958 12781 6010
rect 20155 5958 20207 6010
rect 20219 5958 20271 6010
rect 20283 5958 20335 6010
rect 20347 5958 20399 6010
rect 20411 5958 20463 6010
rect 27837 5958 27889 6010
rect 27901 5958 27953 6010
rect 27965 5958 28017 6010
rect 28029 5958 28081 6010
rect 28093 5958 28145 6010
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 8484 5652 8536 5704
rect 29000 5856 29052 5908
rect 29184 5899 29236 5908
rect 29184 5865 29193 5899
rect 29193 5865 29227 5899
rect 29227 5865 29236 5899
rect 29184 5856 29236 5865
rect 27712 5788 27764 5840
rect 28264 5788 28316 5840
rect 26608 5720 26660 5772
rect 31300 5695 31352 5704
rect 31300 5661 31309 5695
rect 31309 5661 31343 5695
rect 31343 5661 31352 5695
rect 31300 5652 31352 5661
rect 27620 5516 27672 5568
rect 28356 5516 28408 5568
rect 8632 5414 8684 5466
rect 8696 5414 8748 5466
rect 8760 5414 8812 5466
rect 8824 5414 8876 5466
rect 8888 5414 8940 5466
rect 16314 5414 16366 5466
rect 16378 5414 16430 5466
rect 16442 5414 16494 5466
rect 16506 5414 16558 5466
rect 16570 5414 16622 5466
rect 23996 5414 24048 5466
rect 24060 5414 24112 5466
rect 24124 5414 24176 5466
rect 24188 5414 24240 5466
rect 24252 5414 24304 5466
rect 31678 5414 31730 5466
rect 31742 5414 31794 5466
rect 31806 5414 31858 5466
rect 31870 5414 31922 5466
rect 31934 5414 31986 5466
rect 8208 5312 8260 5364
rect 12164 5244 12216 5296
rect 27160 5244 27212 5296
rect 31208 5312 31260 5364
rect 30656 5244 30708 5296
rect 24400 5176 24452 5228
rect 26240 5108 26292 5160
rect 29368 5151 29420 5160
rect 29368 5117 29377 5151
rect 29377 5117 29411 5151
rect 29411 5117 29420 5151
rect 29368 5108 29420 5117
rect 28356 5015 28408 5024
rect 28356 4981 28365 5015
rect 28365 4981 28399 5015
rect 28399 4981 28408 5015
rect 28356 4972 28408 4981
rect 28448 4972 28500 5024
rect 28908 5015 28960 5024
rect 28908 4981 28917 5015
rect 28917 4981 28951 5015
rect 28951 4981 28960 5015
rect 28908 4972 28960 4981
rect 4791 4870 4843 4922
rect 4855 4870 4907 4922
rect 4919 4870 4971 4922
rect 4983 4870 5035 4922
rect 5047 4870 5099 4922
rect 12473 4870 12525 4922
rect 12537 4870 12589 4922
rect 12601 4870 12653 4922
rect 12665 4870 12717 4922
rect 12729 4870 12781 4922
rect 20155 4870 20207 4922
rect 20219 4870 20271 4922
rect 20283 4870 20335 4922
rect 20347 4870 20399 4922
rect 20411 4870 20463 4922
rect 27837 4870 27889 4922
rect 27901 4870 27953 4922
rect 27965 4870 28017 4922
rect 28029 4870 28081 4922
rect 28093 4870 28145 4922
rect 28908 4768 28960 4820
rect 26148 4700 26200 4752
rect 27252 4632 27304 4684
rect 26792 4564 26844 4616
rect 8632 4326 8684 4378
rect 8696 4326 8748 4378
rect 8760 4326 8812 4378
rect 8824 4326 8876 4378
rect 8888 4326 8940 4378
rect 16314 4326 16366 4378
rect 16378 4326 16430 4378
rect 16442 4326 16494 4378
rect 16506 4326 16558 4378
rect 16570 4326 16622 4378
rect 23996 4326 24048 4378
rect 24060 4326 24112 4378
rect 24124 4326 24176 4378
rect 24188 4326 24240 4378
rect 24252 4326 24304 4378
rect 31678 4326 31730 4378
rect 31742 4326 31794 4378
rect 31806 4326 31858 4378
rect 31870 4326 31922 4378
rect 31934 4326 31986 4378
rect 30564 4088 30616 4140
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 28356 3884 28408 3936
rect 30472 3927 30524 3936
rect 30472 3893 30481 3927
rect 30481 3893 30515 3927
rect 30515 3893 30524 3927
rect 30472 3884 30524 3893
rect 31300 3927 31352 3936
rect 31300 3893 31309 3927
rect 31309 3893 31343 3927
rect 31343 3893 31352 3927
rect 31300 3884 31352 3893
rect 4791 3782 4843 3834
rect 4855 3782 4907 3834
rect 4919 3782 4971 3834
rect 4983 3782 5035 3834
rect 5047 3782 5099 3834
rect 12473 3782 12525 3834
rect 12537 3782 12589 3834
rect 12601 3782 12653 3834
rect 12665 3782 12717 3834
rect 12729 3782 12781 3834
rect 20155 3782 20207 3834
rect 20219 3782 20271 3834
rect 20283 3782 20335 3834
rect 20347 3782 20399 3834
rect 20411 3782 20463 3834
rect 27837 3782 27889 3834
rect 27901 3782 27953 3834
rect 27965 3782 28017 3834
rect 28029 3782 28081 3834
rect 28093 3782 28145 3834
rect 30472 3680 30524 3732
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 31300 3519 31352 3528
rect 31300 3485 31309 3519
rect 31309 3485 31343 3519
rect 31343 3485 31352 3519
rect 31300 3476 31352 3485
rect 8632 3238 8684 3290
rect 8696 3238 8748 3290
rect 8760 3238 8812 3290
rect 8824 3238 8876 3290
rect 8888 3238 8940 3290
rect 16314 3238 16366 3290
rect 16378 3238 16430 3290
rect 16442 3238 16494 3290
rect 16506 3238 16558 3290
rect 16570 3238 16622 3290
rect 23996 3238 24048 3290
rect 24060 3238 24112 3290
rect 24124 3238 24176 3290
rect 24188 3238 24240 3290
rect 24252 3238 24304 3290
rect 31678 3238 31730 3290
rect 31742 3238 31794 3290
rect 31806 3238 31858 3290
rect 31870 3238 31922 3290
rect 31934 3238 31986 3290
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 4791 2694 4843 2746
rect 4855 2694 4907 2746
rect 4919 2694 4971 2746
rect 4983 2694 5035 2746
rect 5047 2694 5099 2746
rect 12473 2694 12525 2746
rect 12537 2694 12589 2746
rect 12601 2694 12653 2746
rect 12665 2694 12717 2746
rect 12729 2694 12781 2746
rect 20155 2694 20207 2746
rect 20219 2694 20271 2746
rect 20283 2694 20335 2746
rect 20347 2694 20399 2746
rect 20411 2694 20463 2746
rect 27837 2694 27889 2746
rect 27901 2694 27953 2746
rect 27965 2694 28017 2746
rect 28029 2694 28081 2746
rect 28093 2694 28145 2746
rect 1400 2388 1452 2440
rect 8632 2150 8684 2202
rect 8696 2150 8748 2202
rect 8760 2150 8812 2202
rect 8824 2150 8876 2202
rect 8888 2150 8940 2202
rect 16314 2150 16366 2202
rect 16378 2150 16430 2202
rect 16442 2150 16494 2202
rect 16506 2150 16558 2202
rect 16570 2150 16622 2202
rect 23996 2150 24048 2202
rect 24060 2150 24112 2202
rect 24124 2150 24176 2202
rect 24188 2150 24240 2202
rect 24252 2150 24304 2202
rect 31678 2150 31730 2202
rect 31742 2150 31794 2202
rect 31806 2150 31858 2202
rect 31870 2150 31922 2202
rect 31934 2150 31986 2202
<< metal2 >>
rect 938 34350 994 35150
rect 2134 34490 2190 35150
rect 2134 34462 2268 34490
rect 2134 34350 2190 34462
rect 952 32434 980 34350
rect 1582 32600 1638 32609
rect 1582 32535 1638 32544
rect 940 32428 992 32434
rect 940 32370 992 32376
rect 1596 32026 1624 32535
rect 2240 32434 2268 34462
rect 3330 34350 3386 35150
rect 3974 34776 4030 34785
rect 3974 34711 4030 34720
rect 2870 33416 2926 33425
rect 2870 33351 2926 33360
rect 2884 32434 2912 33351
rect 2228 32428 2280 32434
rect 2228 32370 2280 32376
rect 2872 32428 2924 32434
rect 2872 32370 2924 32376
rect 1584 32020 1636 32026
rect 1584 31962 1636 31968
rect 1584 31136 1636 31142
rect 1584 31078 1636 31084
rect 1596 30977 1624 31078
rect 1582 30968 1638 30977
rect 1582 30903 1638 30912
rect 2688 30388 2740 30394
rect 2688 30330 2740 30336
rect 1584 30184 1636 30190
rect 1582 30152 1584 30161
rect 1636 30152 1638 30161
rect 1582 30087 1638 30096
rect 1584 28552 1636 28558
rect 1582 28520 1584 28529
rect 1636 28520 1638 28529
rect 1582 28455 1638 28464
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1596 27713 1624 27814
rect 1582 27704 1638 27713
rect 1582 27639 1638 27648
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 26081 1624 26318
rect 1582 26072 1638 26081
rect 1582 26007 1638 26016
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1584 23656 1636 23662
rect 1582 23624 1584 23633
rect 1636 23624 1638 23633
rect 1582 23559 1638 23568
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 1596 22817 1624 23054
rect 1582 22808 1638 22817
rect 1582 22743 1638 22752
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21185 1624 21286
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1584 20392 1636 20398
rect 1582 20360 1584 20369
rect 1636 20360 1638 20369
rect 1582 20295 1638 20304
rect 1584 18760 1636 18766
rect 1582 18728 1584 18737
rect 1636 18728 1638 18737
rect 1582 18663 1638 18672
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17921 1624 18022
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16289 1624 16594
rect 1582 16280 1638 16289
rect 1582 16215 1638 16224
rect 1584 15496 1636 15502
rect 1582 15464 1584 15473
rect 1636 15464 1638 15473
rect 1582 15399 1638 15408
rect 1584 13864 1636 13870
rect 1582 13832 1584 13841
rect 1636 13832 1638 13841
rect 1582 13767 1638 13776
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 13025 1624 13262
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 11393 1624 11494
rect 1582 11384 1638 11393
rect 1582 11319 1638 11328
rect 1584 10600 1636 10606
rect 1582 10568 1584 10577
rect 1636 10568 1638 10577
rect 1582 10503 1638 10512
rect 1584 8968 1636 8974
rect 1582 8936 1584 8945
rect 1636 8936 1638 8945
rect 1582 8871 1638 8880
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 8129 1624 8298
rect 1582 8120 1638 8129
rect 1582 8055 1638 8064
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6497 1624 6734
rect 1582 6488 1638 6497
rect 1582 6423 1638 6432
rect 2700 6225 2728 30330
rect 3884 27396 3936 27402
rect 3884 27338 3936 27344
rect 3896 17785 3924 27338
rect 3988 20369 4016 34711
rect 4526 34490 4582 35150
rect 5722 34490 5778 35150
rect 6642 34912 6698 34921
rect 6642 34847 6698 34856
rect 4526 34462 4660 34490
rect 4526 34350 4582 34462
rect 4342 32464 4398 32473
rect 4632 32434 4660 34462
rect 5722 34462 5856 34490
rect 5722 34350 5778 34462
rect 5828 32434 5856 34462
rect 4342 32399 4398 32408
rect 4620 32428 4672 32434
rect 4356 31754 4384 32399
rect 4620 32370 4672 32376
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 4791 32124 5099 32133
rect 4791 32122 4797 32124
rect 4853 32122 4877 32124
rect 4933 32122 4957 32124
rect 5013 32122 5037 32124
rect 5093 32122 5099 32124
rect 4853 32070 4855 32122
rect 5035 32070 5037 32122
rect 4791 32068 4797 32070
rect 4853 32068 4877 32070
rect 4933 32068 4957 32070
rect 5013 32068 5037 32070
rect 5093 32068 5099 32070
rect 4791 32059 5099 32068
rect 4356 31726 5396 31754
rect 4791 31036 5099 31045
rect 4791 31034 4797 31036
rect 4853 31034 4877 31036
rect 4933 31034 4957 31036
rect 5013 31034 5037 31036
rect 5093 31034 5099 31036
rect 4853 30982 4855 31034
rect 5035 30982 5037 31034
rect 4791 30980 4797 30982
rect 4853 30980 4877 30982
rect 4933 30980 4957 30982
rect 5013 30980 5037 30982
rect 5093 30980 5099 30982
rect 4791 30971 5099 30980
rect 4068 30864 4120 30870
rect 4068 30806 4120 30812
rect 3974 20360 4030 20369
rect 3974 20295 4030 20304
rect 3882 17776 3938 17785
rect 3882 17711 3938 17720
rect 4080 12753 4108 30806
rect 4791 29948 5099 29957
rect 4791 29946 4797 29948
rect 4853 29946 4877 29948
rect 4933 29946 4957 29948
rect 5013 29946 5037 29948
rect 5093 29946 5099 29948
rect 4853 29894 4855 29946
rect 5035 29894 5037 29946
rect 4791 29892 4797 29894
rect 4853 29892 4877 29894
rect 4933 29892 4957 29894
rect 5013 29892 5037 29894
rect 5093 29892 5099 29894
rect 4791 29883 5099 29892
rect 4526 29744 4582 29753
rect 4526 29679 4582 29688
rect 4160 28416 4212 28422
rect 4160 28358 4212 28364
rect 4172 24410 4200 28358
rect 4252 24880 4304 24886
rect 4252 24822 4304 24828
rect 4160 24404 4212 24410
rect 4160 24346 4212 24352
rect 4264 23322 4292 24822
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4356 23866 4384 24686
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 4252 23316 4304 23322
rect 4252 23258 4304 23264
rect 4264 22094 4292 23258
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4172 22066 4292 22094
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4172 11014 4200 22066
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4264 6866 4292 21898
rect 4448 9994 4476 22646
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 2686 6216 2742 6225
rect 2686 6151 2742 6160
rect 4540 6118 4568 29679
rect 4791 28860 5099 28869
rect 4791 28858 4797 28860
rect 4853 28858 4877 28860
rect 4933 28858 4957 28860
rect 5013 28858 5037 28860
rect 5093 28858 5099 28860
rect 4853 28806 4855 28858
rect 5035 28806 5037 28858
rect 4791 28804 4797 28806
rect 4853 28804 4877 28806
rect 4933 28804 4957 28806
rect 5013 28804 5037 28806
rect 5093 28804 5099 28806
rect 4791 28795 5099 28804
rect 4791 27772 5099 27781
rect 4791 27770 4797 27772
rect 4853 27770 4877 27772
rect 4933 27770 4957 27772
rect 5013 27770 5037 27772
rect 5093 27770 5099 27772
rect 4853 27718 4855 27770
rect 5035 27718 5037 27770
rect 4791 27716 4797 27718
rect 4853 27716 4877 27718
rect 4933 27716 4957 27718
rect 5013 27716 5037 27718
rect 5093 27716 5099 27718
rect 4791 27707 5099 27716
rect 5262 26888 5318 26897
rect 5262 26823 5318 26832
rect 4791 26684 5099 26693
rect 4791 26682 4797 26684
rect 4853 26682 4877 26684
rect 4933 26682 4957 26684
rect 5013 26682 5037 26684
rect 5093 26682 5099 26684
rect 4853 26630 4855 26682
rect 5035 26630 5037 26682
rect 4791 26628 4797 26630
rect 4853 26628 4877 26630
rect 4933 26628 4957 26630
rect 5013 26628 5037 26630
rect 5093 26628 5099 26630
rect 4791 26619 5099 26628
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 4791 25596 5099 25605
rect 4791 25594 4797 25596
rect 4853 25594 4877 25596
rect 4933 25594 4957 25596
rect 5013 25594 5037 25596
rect 5093 25594 5099 25596
rect 4853 25542 4855 25594
rect 5035 25542 5037 25594
rect 4791 25540 4797 25542
rect 4853 25540 4877 25542
rect 4933 25540 4957 25542
rect 5013 25540 5037 25542
rect 5093 25540 5099 25542
rect 4791 25531 5099 25540
rect 5184 24818 5212 26386
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 4791 24508 5099 24517
rect 4791 24506 4797 24508
rect 4853 24506 4877 24508
rect 4933 24506 4957 24508
rect 5013 24506 5037 24508
rect 5093 24506 5099 24508
rect 4853 24454 4855 24506
rect 5035 24454 5037 24506
rect 4791 24452 4797 24454
rect 4853 24452 4877 24454
rect 4933 24452 4957 24454
rect 5013 24452 5037 24454
rect 5093 24452 5099 24454
rect 4791 24443 5099 24452
rect 4791 23420 5099 23429
rect 4791 23418 4797 23420
rect 4853 23418 4877 23420
rect 4933 23418 4957 23420
rect 5013 23418 5037 23420
rect 5093 23418 5099 23420
rect 4853 23366 4855 23418
rect 5035 23366 5037 23418
rect 4791 23364 4797 23366
rect 4853 23364 4877 23366
rect 4933 23364 4957 23366
rect 5013 23364 5037 23366
rect 5093 23364 5099 23366
rect 4791 23355 5099 23364
rect 5080 23112 5132 23118
rect 5080 23054 5132 23060
rect 5092 22556 5120 23054
rect 5184 22710 5212 24754
rect 5172 22704 5224 22710
rect 5172 22646 5224 22652
rect 5092 22528 5212 22556
rect 4791 22332 5099 22341
rect 4791 22330 4797 22332
rect 4853 22330 4877 22332
rect 4933 22330 4957 22332
rect 5013 22330 5037 22332
rect 5093 22330 5099 22332
rect 4853 22278 4855 22330
rect 5035 22278 5037 22330
rect 4791 22276 4797 22278
rect 4853 22276 4877 22278
rect 4933 22276 4957 22278
rect 5013 22276 5037 22278
rect 5093 22276 5099 22278
rect 4791 22267 5099 22276
rect 4712 22024 4764 22030
rect 4710 21992 4712 22001
rect 4764 21992 4766 22001
rect 4710 21927 4766 21936
rect 4791 21244 5099 21253
rect 4791 21242 4797 21244
rect 4853 21242 4877 21244
rect 4933 21242 4957 21244
rect 5013 21242 5037 21244
rect 5093 21242 5099 21244
rect 4853 21190 4855 21242
rect 5035 21190 5037 21242
rect 4791 21188 4797 21190
rect 4853 21188 4877 21190
rect 4933 21188 4957 21190
rect 5013 21188 5037 21190
rect 5093 21188 5099 21190
rect 4791 21179 5099 21188
rect 4791 20156 5099 20165
rect 4791 20154 4797 20156
rect 4853 20154 4877 20156
rect 4933 20154 4957 20156
rect 5013 20154 5037 20156
rect 5093 20154 5099 20156
rect 4853 20102 4855 20154
rect 5035 20102 5037 20154
rect 4791 20100 4797 20102
rect 4853 20100 4877 20102
rect 4933 20100 4957 20102
rect 5013 20100 5037 20102
rect 5093 20100 5099 20102
rect 4791 20091 5099 20100
rect 4791 19068 5099 19077
rect 4791 19066 4797 19068
rect 4853 19066 4877 19068
rect 4933 19066 4957 19068
rect 5013 19066 5037 19068
rect 5093 19066 5099 19068
rect 4853 19014 4855 19066
rect 5035 19014 5037 19066
rect 4791 19012 4797 19014
rect 4853 19012 4877 19014
rect 4933 19012 4957 19014
rect 5013 19012 5037 19014
rect 5093 19012 5099 19014
rect 4791 19003 5099 19012
rect 4791 17980 5099 17989
rect 4791 17978 4797 17980
rect 4853 17978 4877 17980
rect 4933 17978 4957 17980
rect 5013 17978 5037 17980
rect 5093 17978 5099 17980
rect 4853 17926 4855 17978
rect 5035 17926 5037 17978
rect 4791 17924 4797 17926
rect 4853 17924 4877 17926
rect 4933 17924 4957 17926
rect 5013 17924 5037 17926
rect 5093 17924 5099 17926
rect 4791 17915 5099 17924
rect 4791 16892 5099 16901
rect 4791 16890 4797 16892
rect 4853 16890 4877 16892
rect 4933 16890 4957 16892
rect 5013 16890 5037 16892
rect 5093 16890 5099 16892
rect 4853 16838 4855 16890
rect 5035 16838 5037 16890
rect 4791 16836 4797 16838
rect 4853 16836 4877 16838
rect 4933 16836 4957 16838
rect 5013 16836 5037 16838
rect 5093 16836 5099 16838
rect 4791 16827 5099 16836
rect 4791 15804 5099 15813
rect 4791 15802 4797 15804
rect 4853 15802 4877 15804
rect 4933 15802 4957 15804
rect 5013 15802 5037 15804
rect 5093 15802 5099 15804
rect 4853 15750 4855 15802
rect 5035 15750 5037 15802
rect 4791 15748 4797 15750
rect 4853 15748 4877 15750
rect 4933 15748 4957 15750
rect 5013 15748 5037 15750
rect 5093 15748 5099 15750
rect 4791 15739 5099 15748
rect 4791 14716 5099 14725
rect 4791 14714 4797 14716
rect 4853 14714 4877 14716
rect 4933 14714 4957 14716
rect 5013 14714 5037 14716
rect 5093 14714 5099 14716
rect 4853 14662 4855 14714
rect 5035 14662 5037 14714
rect 4791 14660 4797 14662
rect 4853 14660 4877 14662
rect 4933 14660 4957 14662
rect 5013 14660 5037 14662
rect 5093 14660 5099 14662
rect 4791 14651 5099 14660
rect 4791 13628 5099 13637
rect 4791 13626 4797 13628
rect 4853 13626 4877 13628
rect 4933 13626 4957 13628
rect 5013 13626 5037 13628
rect 5093 13626 5099 13628
rect 4853 13574 4855 13626
rect 5035 13574 5037 13626
rect 4791 13572 4797 13574
rect 4853 13572 4877 13574
rect 4933 13572 4957 13574
rect 5013 13572 5037 13574
rect 5093 13572 5099 13574
rect 4791 13563 5099 13572
rect 4791 12540 5099 12549
rect 4791 12538 4797 12540
rect 4853 12538 4877 12540
rect 4933 12538 4957 12540
rect 5013 12538 5037 12540
rect 5093 12538 5099 12540
rect 4853 12486 4855 12538
rect 5035 12486 5037 12538
rect 4791 12484 4797 12486
rect 4853 12484 4877 12486
rect 4933 12484 4957 12486
rect 5013 12484 5037 12486
rect 5093 12484 5099 12486
rect 4791 12475 5099 12484
rect 4791 11452 5099 11461
rect 4791 11450 4797 11452
rect 4853 11450 4877 11452
rect 4933 11450 4957 11452
rect 5013 11450 5037 11452
rect 5093 11450 5099 11452
rect 4853 11398 4855 11450
rect 5035 11398 5037 11450
rect 4791 11396 4797 11398
rect 4853 11396 4877 11398
rect 4933 11396 4957 11398
rect 5013 11396 5037 11398
rect 5093 11396 5099 11398
rect 4791 11387 5099 11396
rect 4791 10364 5099 10373
rect 4791 10362 4797 10364
rect 4853 10362 4877 10364
rect 4933 10362 4957 10364
rect 5013 10362 5037 10364
rect 5093 10362 5099 10364
rect 4853 10310 4855 10362
rect 5035 10310 5037 10362
rect 4791 10308 4797 10310
rect 4853 10308 4877 10310
rect 4933 10308 4957 10310
rect 5013 10308 5037 10310
rect 5093 10308 5099 10310
rect 4791 10299 5099 10308
rect 4791 9276 5099 9285
rect 4791 9274 4797 9276
rect 4853 9274 4877 9276
rect 4933 9274 4957 9276
rect 5013 9274 5037 9276
rect 5093 9274 5099 9276
rect 4853 9222 4855 9274
rect 5035 9222 5037 9274
rect 4791 9220 4797 9222
rect 4853 9220 4877 9222
rect 4933 9220 4957 9222
rect 5013 9220 5037 9222
rect 5093 9220 5099 9222
rect 4791 9211 5099 9220
rect 4791 8188 5099 8197
rect 4791 8186 4797 8188
rect 4853 8186 4877 8188
rect 4933 8186 4957 8188
rect 5013 8186 5037 8188
rect 5093 8186 5099 8188
rect 4853 8134 4855 8186
rect 5035 8134 5037 8186
rect 4791 8132 4797 8134
rect 4853 8132 4877 8134
rect 4933 8132 4957 8134
rect 5013 8132 5037 8134
rect 5093 8132 5099 8134
rect 4791 8123 5099 8132
rect 4791 7100 5099 7109
rect 4791 7098 4797 7100
rect 4853 7098 4877 7100
rect 4933 7098 4957 7100
rect 5013 7098 5037 7100
rect 5093 7098 5099 7100
rect 4853 7046 4855 7098
rect 5035 7046 5037 7098
rect 4791 7044 4797 7046
rect 4853 7044 4877 7046
rect 4933 7044 4957 7046
rect 5013 7044 5037 7046
rect 5093 7044 5099 7046
rect 4791 7035 5099 7044
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4791 6012 5099 6021
rect 4791 6010 4797 6012
rect 4853 6010 4877 6012
rect 4933 6010 4957 6012
rect 5013 6010 5037 6012
rect 5093 6010 5099 6012
rect 4853 5958 4855 6010
rect 5035 5958 5037 6010
rect 4791 5956 4797 5958
rect 4853 5956 4877 5958
rect 4933 5956 4957 5958
rect 5013 5956 5037 5958
rect 5093 5956 5099 5958
rect 4791 5947 5099 5956
rect 1584 5704 1636 5710
rect 1582 5672 1584 5681
rect 1636 5672 1638 5681
rect 1582 5607 1638 5616
rect 5184 5273 5212 22528
rect 5276 10538 5304 26823
rect 5368 23594 5396 31726
rect 6368 28688 6420 28694
rect 6368 28630 6420 28636
rect 6380 27334 6408 28630
rect 6368 27328 6420 27334
rect 6368 27270 6420 27276
rect 6276 27056 6328 27062
rect 6276 26998 6328 27004
rect 6288 25498 6316 26998
rect 6380 25498 6408 27270
rect 6276 25492 6328 25498
rect 6276 25434 6328 25440
rect 6368 25492 6420 25498
rect 6368 25434 6420 25440
rect 5816 25152 5868 25158
rect 5816 25094 5868 25100
rect 5828 24342 5856 25094
rect 5998 24712 6054 24721
rect 5998 24647 6000 24656
rect 6052 24647 6054 24656
rect 6000 24618 6052 24624
rect 5816 24336 5868 24342
rect 5816 24278 5868 24284
rect 5814 24168 5870 24177
rect 5814 24103 5870 24112
rect 5908 24132 5960 24138
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 5368 22098 5396 23530
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5460 21690 5488 23122
rect 5644 22778 5672 24006
rect 5828 23322 5856 24103
rect 5908 24074 5960 24080
rect 5920 23322 5948 24074
rect 5816 23316 5868 23322
rect 5736 23276 5816 23304
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5552 21622 5580 22170
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5446 9616 5502 9625
rect 5446 9551 5502 9560
rect 5460 8974 5488 9551
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5736 8401 5764 23276
rect 5816 23258 5868 23264
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 6656 23050 6684 34847
rect 6918 34350 6974 35150
rect 8114 34490 8170 35150
rect 9310 34490 9366 35150
rect 8114 34462 8248 34490
rect 8114 34350 8170 34462
rect 8220 32434 8248 34462
rect 9310 34462 9444 34490
rect 9310 34350 9366 34462
rect 9128 33516 9180 33522
rect 9128 33458 9180 33464
rect 8632 32668 8940 32677
rect 8632 32666 8638 32668
rect 8694 32666 8718 32668
rect 8774 32666 8798 32668
rect 8854 32666 8878 32668
rect 8934 32666 8940 32668
rect 8694 32614 8696 32666
rect 8876 32614 8878 32666
rect 8632 32612 8638 32614
rect 8694 32612 8718 32614
rect 8774 32612 8798 32614
rect 8854 32612 8878 32614
rect 8934 32612 8940 32614
rect 8632 32603 8940 32612
rect 8208 32428 8260 32434
rect 8208 32370 8260 32376
rect 8632 31580 8940 31589
rect 8632 31578 8638 31580
rect 8694 31578 8718 31580
rect 8774 31578 8798 31580
rect 8854 31578 8878 31580
rect 8934 31578 8940 31580
rect 8694 31526 8696 31578
rect 8876 31526 8878 31578
rect 8632 31524 8638 31526
rect 8694 31524 8718 31526
rect 8774 31524 8798 31526
rect 8854 31524 8878 31526
rect 8934 31524 8940 31526
rect 8632 31515 8940 31524
rect 8206 31376 8262 31385
rect 8206 31311 8262 31320
rect 7840 29504 7892 29510
rect 7840 29446 7892 29452
rect 7378 29200 7434 29209
rect 7378 29135 7434 29144
rect 7392 27402 7420 29135
rect 7380 27396 7432 27402
rect 7380 27338 7432 27344
rect 7288 27328 7340 27334
rect 7288 27270 7340 27276
rect 7300 26790 7328 27270
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 6828 26308 6880 26314
rect 6828 26250 6880 26256
rect 6840 26194 6868 26250
rect 7300 26228 7328 26726
rect 7472 26240 7524 26246
rect 7300 26200 7472 26228
rect 6840 26166 6960 26194
rect 7472 26182 7524 26188
rect 6828 25424 6880 25430
rect 6828 25366 6880 25372
rect 6840 24426 6868 25366
rect 6932 24834 6960 26166
rect 7484 25702 7512 26182
rect 7852 25922 7880 29446
rect 8116 27872 8168 27878
rect 8116 27814 8168 27820
rect 8022 27432 8078 27441
rect 8022 27367 8024 27376
rect 8076 27367 8078 27376
rect 8024 27338 8076 27344
rect 7932 26308 7984 26314
rect 7932 26250 7984 26256
rect 7944 26042 7972 26250
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 7852 25894 7972 25922
rect 7656 25764 7708 25770
rect 7656 25706 7708 25712
rect 7472 25696 7524 25702
rect 7472 25638 7524 25644
rect 7484 25430 7512 25638
rect 7472 25424 7524 25430
rect 7472 25366 7524 25372
rect 6932 24806 7052 24834
rect 6840 24410 6960 24426
rect 6840 24404 6972 24410
rect 6840 24398 6920 24404
rect 6920 24346 6972 24352
rect 6918 24304 6974 24313
rect 6918 24239 6974 24248
rect 6932 24138 6960 24239
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 6932 23610 6960 24074
rect 7024 23866 7052 24806
rect 7668 24138 7696 25706
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 6748 23582 6960 23610
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 6552 23044 6604 23050
rect 6552 22986 6604 22992
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 5816 22500 5868 22506
rect 5816 22442 5868 22448
rect 5828 21690 5856 22442
rect 5920 22234 5948 22510
rect 6104 22438 6132 22918
rect 6368 22500 6420 22506
rect 6368 22442 6420 22448
rect 6092 22432 6144 22438
rect 6092 22374 6144 22380
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 6000 20800 6052 20806
rect 6104 20788 6132 22374
rect 6380 22234 6408 22442
rect 6564 22234 6592 22986
rect 6368 22228 6420 22234
rect 6368 22170 6420 22176
rect 6552 22228 6604 22234
rect 6552 22170 6604 22176
rect 6564 21894 6592 22170
rect 6552 21888 6604 21894
rect 6748 21865 6776 23582
rect 6826 23488 6882 23497
rect 6826 23423 6882 23432
rect 6552 21830 6604 21836
rect 6734 21856 6790 21865
rect 6052 20760 6132 20788
rect 6000 20742 6052 20748
rect 6012 19174 6040 20742
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6564 9625 6592 21830
rect 6734 21791 6790 21800
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6656 18154 6684 19110
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6550 9616 6606 9625
rect 6550 9551 6606 9560
rect 6840 9178 6868 23423
rect 7116 22778 7144 23598
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6932 9586 6960 19654
rect 7300 11257 7328 23802
rect 7668 22982 7696 24074
rect 7760 24070 7788 24550
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7484 21146 7512 22918
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7576 21622 7604 21830
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7392 20398 7420 20742
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 19718 7420 20334
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7484 19854 7512 20266
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7576 12434 7604 21558
rect 7760 21185 7788 24006
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7852 22137 7880 23462
rect 7838 22128 7894 22137
rect 7838 22063 7894 22072
rect 7944 22094 7972 25894
rect 8036 23118 8064 27338
rect 8128 25702 8156 27814
rect 8116 25696 8168 25702
rect 8116 25638 8168 25644
rect 8024 23112 8076 23118
rect 8220 23089 8248 31311
rect 9036 30932 9088 30938
rect 9036 30874 9088 30880
rect 8632 30492 8940 30501
rect 8632 30490 8638 30492
rect 8694 30490 8718 30492
rect 8774 30490 8798 30492
rect 8854 30490 8878 30492
rect 8934 30490 8940 30492
rect 8694 30438 8696 30490
rect 8876 30438 8878 30490
rect 8632 30436 8638 30438
rect 8694 30436 8718 30438
rect 8774 30436 8798 30438
rect 8854 30436 8878 30438
rect 8934 30436 8940 30438
rect 8632 30427 8940 30436
rect 9048 30326 9076 30874
rect 9036 30320 9088 30326
rect 9036 30262 9088 30268
rect 8632 29404 8940 29413
rect 8632 29402 8638 29404
rect 8694 29402 8718 29404
rect 8774 29402 8798 29404
rect 8854 29402 8878 29404
rect 8934 29402 8940 29404
rect 8694 29350 8696 29402
rect 8876 29350 8878 29402
rect 8632 29348 8638 29350
rect 8694 29348 8718 29350
rect 8774 29348 8798 29350
rect 8854 29348 8878 29350
rect 8934 29348 8940 29350
rect 8632 29339 8940 29348
rect 9048 29238 9076 30262
rect 9036 29232 9088 29238
rect 9036 29174 9088 29180
rect 9036 28552 9088 28558
rect 9036 28494 9088 28500
rect 8632 28316 8940 28325
rect 8632 28314 8638 28316
rect 8694 28314 8718 28316
rect 8774 28314 8798 28316
rect 8854 28314 8878 28316
rect 8934 28314 8940 28316
rect 8694 28262 8696 28314
rect 8876 28262 8878 28314
rect 8632 28260 8638 28262
rect 8694 28260 8718 28262
rect 8774 28260 8798 28262
rect 8854 28260 8878 28262
rect 8934 28260 8940 28262
rect 8632 28251 8940 28260
rect 8300 27940 8352 27946
rect 8300 27882 8352 27888
rect 8206 23080 8262 23089
rect 8024 23054 8076 23060
rect 8128 23038 8206 23066
rect 8128 22710 8156 23038
rect 8206 23015 8262 23024
rect 8206 22808 8262 22817
rect 8206 22743 8208 22752
rect 8260 22743 8262 22752
rect 8208 22714 8260 22720
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 8220 22409 8248 22714
rect 8206 22400 8262 22409
rect 8206 22335 8262 22344
rect 7944 22066 8248 22094
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7746 21176 7802 21185
rect 7656 21140 7708 21146
rect 7746 21111 7802 21120
rect 7656 21082 7708 21088
rect 7668 20262 7696 21082
rect 7944 20262 7972 21286
rect 8024 20800 8076 20806
rect 8024 20742 8076 20748
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7668 19417 7696 20198
rect 7944 20058 7972 20198
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7654 19408 7710 19417
rect 7654 19343 7710 19352
rect 7668 19174 7696 19343
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7392 12406 7604 12434
rect 7286 11248 7342 11257
rect 7286 11183 7342 11192
rect 7392 11121 7420 12406
rect 7378 11112 7434 11121
rect 7378 11047 7434 11056
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 5722 8392 5778 8401
rect 5722 8327 5778 8336
rect 7668 7886 7696 19110
rect 7944 18630 7972 19790
rect 8036 19786 8064 20742
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 8036 19446 8064 19722
rect 8024 19440 8076 19446
rect 8024 19382 8076 19388
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7944 9382 7972 18566
rect 8128 10266 8156 20742
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 8220 5370 8248 22066
rect 8312 21146 8340 27882
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8404 27674 8432 27814
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 9048 27606 9076 28494
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 9140 27418 9168 33458
rect 9416 32434 9444 34462
rect 10506 34350 10562 35150
rect 11702 34490 11758 35150
rect 12898 34490 12954 35150
rect 11702 34462 11836 34490
rect 11702 34350 11758 34462
rect 10140 33380 10192 33386
rect 10140 33322 10192 33328
rect 9588 32768 9640 32774
rect 9588 32710 9640 32716
rect 9404 32428 9456 32434
rect 9404 32370 9456 32376
rect 9600 31754 9628 32710
rect 9048 27390 9168 27418
rect 9232 31726 9628 31754
rect 10046 31784 10102 31793
rect 9048 27334 9076 27390
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 8632 27228 8940 27237
rect 8632 27226 8638 27228
rect 8694 27226 8718 27228
rect 8774 27226 8798 27228
rect 8854 27226 8878 27228
rect 8934 27226 8940 27228
rect 8694 27174 8696 27226
rect 8876 27174 8878 27226
rect 8632 27172 8638 27174
rect 8694 27172 8718 27174
rect 8774 27172 8798 27174
rect 8854 27172 8878 27174
rect 8934 27172 8940 27174
rect 8632 27163 8940 27172
rect 8484 27124 8536 27130
rect 8484 27066 8536 27072
rect 8390 25800 8446 25809
rect 8390 25735 8446 25744
rect 8404 24818 8432 25735
rect 8496 25498 8524 27066
rect 8632 26140 8940 26149
rect 8632 26138 8638 26140
rect 8694 26138 8718 26140
rect 8774 26138 8798 26140
rect 8854 26138 8878 26140
rect 8934 26138 8940 26140
rect 8694 26086 8696 26138
rect 8876 26086 8878 26138
rect 8632 26084 8638 26086
rect 8694 26084 8718 26086
rect 8774 26084 8798 26086
rect 8854 26084 8878 26086
rect 8934 26084 8940 26086
rect 8632 26075 8940 26084
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8588 25140 8616 25774
rect 9048 25362 9076 27270
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9036 25356 9088 25362
rect 9036 25298 9088 25304
rect 8496 25112 8616 25140
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8496 24614 8524 25112
rect 8632 25052 8940 25061
rect 8632 25050 8638 25052
rect 8694 25050 8718 25052
rect 8774 25050 8798 25052
rect 8854 25050 8878 25052
rect 8934 25050 8940 25052
rect 8694 24998 8696 25050
rect 8876 24998 8878 25050
rect 8632 24996 8638 24998
rect 8694 24996 8718 24998
rect 8774 24996 8798 24998
rect 8854 24996 8878 24998
rect 8934 24996 8940 24998
rect 8632 24987 8940 24996
rect 8484 24608 8536 24614
rect 8404 24568 8484 24596
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8298 21040 8354 21049
rect 8298 20975 8300 20984
rect 8352 20975 8354 20984
rect 8300 20946 8352 20952
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8312 20602 8340 20810
rect 8404 20806 8432 24568
rect 8484 24550 8536 24556
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8496 24138 8524 24346
rect 8956 24274 8984 24550
rect 8944 24268 8996 24274
rect 8944 24210 8996 24216
rect 8484 24132 8536 24138
rect 8484 24074 8536 24080
rect 8632 23964 8940 23973
rect 8632 23962 8638 23964
rect 8694 23962 8718 23964
rect 8774 23962 8798 23964
rect 8854 23962 8878 23964
rect 8934 23962 8940 23964
rect 8694 23910 8696 23962
rect 8876 23910 8878 23962
rect 8632 23908 8638 23910
rect 8694 23908 8718 23910
rect 8774 23908 8798 23910
rect 8854 23908 8878 23910
rect 8934 23908 8940 23910
rect 8632 23899 8940 23908
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8482 23352 8538 23361
rect 8482 23287 8484 23296
rect 8536 23287 8538 23296
rect 8484 23258 8536 23264
rect 8864 23225 8892 23462
rect 8850 23216 8906 23225
rect 8850 23151 8906 23160
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 8632 22876 8940 22885
rect 8632 22874 8638 22876
rect 8694 22874 8718 22876
rect 8774 22874 8798 22876
rect 8854 22874 8878 22876
rect 8934 22874 8940 22876
rect 8694 22822 8696 22874
rect 8876 22822 8878 22874
rect 8632 22820 8638 22822
rect 8694 22820 8718 22822
rect 8774 22820 8798 22822
rect 8854 22820 8878 22822
rect 8934 22820 8940 22822
rect 8632 22811 8940 22820
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8772 22094 8800 22374
rect 8496 22066 8800 22094
rect 8496 21894 8524 22066
rect 8772 22001 8800 22066
rect 8758 21992 8814 22001
rect 8758 21927 8814 21936
rect 8484 21888 8536 21894
rect 9048 21865 9076 22918
rect 9140 22094 9168 26930
rect 9232 24857 9260 31726
rect 10046 31719 10102 31728
rect 10060 30394 10088 31719
rect 10048 30388 10100 30394
rect 10048 30330 10100 30336
rect 9864 30252 9916 30258
rect 9864 30194 9916 30200
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9404 29640 9456 29646
rect 9404 29582 9456 29588
rect 9416 28422 9444 29582
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 9416 27334 9444 28358
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9416 26382 9444 27270
rect 9508 26926 9536 29990
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9600 28218 9628 29514
rect 9876 28762 9904 30194
rect 9954 30152 10010 30161
rect 9954 30087 10010 30096
rect 9968 29782 9996 30087
rect 9956 29776 10008 29782
rect 9956 29718 10008 29724
rect 9954 29064 10010 29073
rect 10152 29050 10180 33322
rect 10508 32972 10560 32978
rect 10508 32914 10560 32920
rect 10520 31754 10548 32914
rect 11808 32434 11836 34462
rect 12898 34462 13032 34490
rect 12898 34350 12954 34462
rect 12070 33960 12126 33969
rect 12070 33895 12126 33904
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11612 32292 11664 32298
rect 11612 32234 11664 32240
rect 10324 31748 10376 31754
rect 10520 31726 10640 31754
rect 10324 31690 10376 31696
rect 10336 30938 10364 31690
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10324 30932 10376 30938
rect 10324 30874 10376 30880
rect 10416 30048 10468 30054
rect 10416 29990 10468 29996
rect 10428 29306 10456 29990
rect 10520 29782 10548 31078
rect 10508 29776 10560 29782
rect 10508 29718 10560 29724
rect 10520 29510 10548 29718
rect 10508 29504 10560 29510
rect 10508 29446 10560 29452
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 10010 29022 10180 29050
rect 9954 28999 9956 29008
rect 10008 28999 10010 29008
rect 9956 28970 10008 28976
rect 9864 28756 9916 28762
rect 9864 28698 9916 28704
rect 10428 28422 10456 29242
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 10508 28008 10560 28014
rect 10322 27976 10378 27985
rect 10508 27950 10560 27956
rect 10322 27911 10378 27920
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9692 27588 9720 27814
rect 9600 27560 9720 27588
rect 9600 27130 9628 27560
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 9496 26920 9548 26926
rect 9496 26862 9548 26868
rect 9588 26784 9640 26790
rect 9588 26726 9640 26732
rect 9312 26376 9364 26382
rect 9310 26344 9312 26353
rect 9404 26376 9456 26382
rect 9364 26344 9366 26353
rect 9404 26318 9456 26324
rect 9310 26279 9366 26288
rect 9312 25764 9364 25770
rect 9416 25752 9444 26318
rect 9364 25724 9444 25752
rect 9312 25706 9364 25712
rect 9218 24848 9274 24857
rect 9324 24818 9352 25706
rect 9494 25392 9550 25401
rect 9494 25327 9550 25336
rect 9218 24783 9274 24792
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9416 23866 9444 24006
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9416 23118 9444 23802
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9324 22098 9352 22442
rect 9140 22066 9260 22094
rect 9128 21956 9180 21962
rect 9128 21898 9180 21904
rect 8484 21830 8536 21836
rect 9034 21856 9090 21865
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8390 20632 8446 20641
rect 8300 20596 8352 20602
rect 8390 20567 8446 20576
rect 8300 20538 8352 20544
rect 8404 9489 8432 20567
rect 8390 9480 8446 9489
rect 8390 9415 8446 9424
rect 8496 5710 8524 21830
rect 8632 21788 8940 21797
rect 9034 21791 9090 21800
rect 8632 21786 8638 21788
rect 8694 21786 8718 21788
rect 8774 21786 8798 21788
rect 8854 21786 8878 21788
rect 8934 21786 8940 21788
rect 8694 21734 8696 21786
rect 8876 21734 8878 21786
rect 8632 21732 8638 21734
rect 8694 21732 8718 21734
rect 8774 21732 8798 21734
rect 8854 21732 8878 21734
rect 8934 21732 8940 21734
rect 8632 21723 8940 21732
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8956 20874 8984 21286
rect 9140 21146 9168 21898
rect 9232 21350 9260 22066
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 8632 20700 8940 20709
rect 8632 20698 8638 20700
rect 8694 20698 8718 20700
rect 8774 20698 8798 20700
rect 8854 20698 8878 20700
rect 8934 20698 8940 20700
rect 8694 20646 8696 20698
rect 8876 20646 8878 20698
rect 8632 20644 8638 20646
rect 8694 20644 8718 20646
rect 8774 20644 8798 20646
rect 8854 20644 8878 20646
rect 8934 20644 8940 20646
rect 8632 20635 8940 20644
rect 9048 20641 9076 20742
rect 9034 20632 9090 20641
rect 9034 20567 9090 20576
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 8632 19612 8940 19621
rect 8632 19610 8638 19612
rect 8694 19610 8718 19612
rect 8774 19610 8798 19612
rect 8854 19610 8878 19612
rect 8934 19610 8940 19612
rect 8694 19558 8696 19610
rect 8876 19558 8878 19610
rect 8632 19556 8638 19558
rect 8694 19556 8718 19558
rect 8774 19556 8798 19558
rect 8854 19556 8878 19558
rect 8934 19556 8940 19558
rect 8632 19547 8940 19556
rect 9048 19514 9076 20198
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 8632 18524 8940 18533
rect 8632 18522 8638 18524
rect 8694 18522 8718 18524
rect 8774 18522 8798 18524
rect 8854 18522 8878 18524
rect 8934 18522 8940 18524
rect 8694 18470 8696 18522
rect 8876 18470 8878 18522
rect 8632 18468 8638 18470
rect 8694 18468 8718 18470
rect 8774 18468 8798 18470
rect 8854 18468 8878 18470
rect 8934 18468 8940 18470
rect 8632 18459 8940 18468
rect 8632 17436 8940 17445
rect 8632 17434 8638 17436
rect 8694 17434 8718 17436
rect 8774 17434 8798 17436
rect 8854 17434 8878 17436
rect 8934 17434 8940 17436
rect 8694 17382 8696 17434
rect 8876 17382 8878 17434
rect 8632 17380 8638 17382
rect 8694 17380 8718 17382
rect 8774 17380 8798 17382
rect 8854 17380 8878 17382
rect 8934 17380 8940 17382
rect 8632 17371 8940 17380
rect 8632 16348 8940 16357
rect 8632 16346 8638 16348
rect 8694 16346 8718 16348
rect 8774 16346 8798 16348
rect 8854 16346 8878 16348
rect 8934 16346 8940 16348
rect 8694 16294 8696 16346
rect 8876 16294 8878 16346
rect 8632 16292 8638 16294
rect 8694 16292 8718 16294
rect 8774 16292 8798 16294
rect 8854 16292 8878 16294
rect 8934 16292 8940 16294
rect 8632 16283 8940 16292
rect 8632 15260 8940 15269
rect 8632 15258 8638 15260
rect 8694 15258 8718 15260
rect 8774 15258 8798 15260
rect 8854 15258 8878 15260
rect 8934 15258 8940 15260
rect 8694 15206 8696 15258
rect 8876 15206 8878 15258
rect 8632 15204 8638 15206
rect 8694 15204 8718 15206
rect 8774 15204 8798 15206
rect 8854 15204 8878 15206
rect 8934 15204 8940 15206
rect 8632 15195 8940 15204
rect 8632 14172 8940 14181
rect 8632 14170 8638 14172
rect 8694 14170 8718 14172
rect 8774 14170 8798 14172
rect 8854 14170 8878 14172
rect 8934 14170 8940 14172
rect 8694 14118 8696 14170
rect 8876 14118 8878 14170
rect 8632 14116 8638 14118
rect 8694 14116 8718 14118
rect 8774 14116 8798 14118
rect 8854 14116 8878 14118
rect 8934 14116 8940 14118
rect 8632 14107 8940 14116
rect 8632 13084 8940 13093
rect 8632 13082 8638 13084
rect 8694 13082 8718 13084
rect 8774 13082 8798 13084
rect 8854 13082 8878 13084
rect 8934 13082 8940 13084
rect 8694 13030 8696 13082
rect 8876 13030 8878 13082
rect 8632 13028 8638 13030
rect 8694 13028 8718 13030
rect 8774 13028 8798 13030
rect 8854 13028 8878 13030
rect 8934 13028 8940 13030
rect 8632 13019 8940 13028
rect 8632 11996 8940 12005
rect 8632 11994 8638 11996
rect 8694 11994 8718 11996
rect 8774 11994 8798 11996
rect 8854 11994 8878 11996
rect 8934 11994 8940 11996
rect 8694 11942 8696 11994
rect 8876 11942 8878 11994
rect 8632 11940 8638 11942
rect 8694 11940 8718 11942
rect 8774 11940 8798 11942
rect 8854 11940 8878 11942
rect 8934 11940 8940 11942
rect 8632 11931 8940 11940
rect 8632 10908 8940 10917
rect 8632 10906 8638 10908
rect 8694 10906 8718 10908
rect 8774 10906 8798 10908
rect 8854 10906 8878 10908
rect 8934 10906 8940 10908
rect 8694 10854 8696 10906
rect 8876 10854 8878 10906
rect 8632 10852 8638 10854
rect 8694 10852 8718 10854
rect 8774 10852 8798 10854
rect 8854 10852 8878 10854
rect 8934 10852 8940 10854
rect 8632 10843 8940 10852
rect 8632 9820 8940 9829
rect 8632 9818 8638 9820
rect 8694 9818 8718 9820
rect 8774 9818 8798 9820
rect 8854 9818 8878 9820
rect 8934 9818 8940 9820
rect 8694 9766 8696 9818
rect 8876 9766 8878 9818
rect 8632 9764 8638 9766
rect 8694 9764 8718 9766
rect 8774 9764 8798 9766
rect 8854 9764 8878 9766
rect 8934 9764 8940 9766
rect 8632 9755 8940 9764
rect 9140 9518 9168 21082
rect 9324 21010 9352 21354
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18630 9260 19110
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8632 8732 8940 8741
rect 8632 8730 8638 8732
rect 8694 8730 8718 8732
rect 8774 8730 8798 8732
rect 8854 8730 8878 8732
rect 8934 8730 8940 8732
rect 8694 8678 8696 8730
rect 8876 8678 8878 8730
rect 8632 8676 8638 8678
rect 8694 8676 8718 8678
rect 8774 8676 8798 8678
rect 8854 8676 8878 8678
rect 8934 8676 8940 8678
rect 8632 8667 8940 8676
rect 9232 7750 9260 18566
rect 9324 10198 9352 20946
rect 9508 20874 9536 25327
rect 9600 24818 9628 26726
rect 9692 26217 9720 27560
rect 10048 27600 10100 27606
rect 10048 27542 10100 27548
rect 10060 27130 10088 27542
rect 10336 27538 10364 27911
rect 10140 27532 10192 27538
rect 10140 27474 10192 27480
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 10416 27532 10468 27538
rect 10416 27474 10468 27480
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9678 26208 9734 26217
rect 9678 26143 9734 26152
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9600 24274 9628 24754
rect 9784 24682 9812 26250
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 9772 24676 9824 24682
rect 9772 24618 9824 24624
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9692 24274 9720 24550
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9600 23594 9628 24074
rect 9678 23760 9734 23769
rect 9678 23695 9734 23704
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9600 23322 9628 23530
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9692 23202 9720 23695
rect 9770 23624 9826 23633
rect 9770 23559 9826 23568
rect 9600 23186 9720 23202
rect 9588 23180 9720 23186
rect 9640 23174 9720 23180
rect 9588 23122 9640 23128
rect 9784 22234 9812 23559
rect 9876 22506 9904 25094
rect 10152 24206 10180 27474
rect 10324 27396 10376 27402
rect 10324 27338 10376 27344
rect 10336 27062 10364 27338
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 10230 25120 10286 25129
rect 10230 25055 10286 25064
rect 10244 24750 10272 25055
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10232 24608 10284 24614
rect 10232 24550 10284 24556
rect 10244 24410 10272 24550
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9600 22030 9628 22170
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9876 21690 9904 22442
rect 9968 21962 9996 23598
rect 10152 23254 10180 24142
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 10244 22094 10272 24210
rect 10336 22642 10364 26998
rect 10428 23730 10456 27474
rect 10520 26790 10548 27950
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10520 23798 10548 26726
rect 10612 26518 10640 31726
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11426 30832 11482 30841
rect 11426 30767 11428 30776
rect 11480 30767 11482 30776
rect 11428 30738 11480 30744
rect 11532 30734 11560 31622
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 11520 30728 11572 30734
rect 11520 30670 11572 30676
rect 11072 29322 11100 30670
rect 11244 30592 11296 30598
rect 11244 30534 11296 30540
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 11164 29714 11192 30330
rect 11256 29850 11284 30534
rect 11244 29844 11296 29850
rect 11244 29786 11296 29792
rect 11256 29714 11284 29786
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 10980 29294 11100 29322
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10888 26790 10916 28358
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10612 25838 10640 26454
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10600 25220 10652 25226
rect 10600 25162 10652 25168
rect 10508 23792 10560 23798
rect 10508 23734 10560 23740
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10428 22710 10456 23666
rect 10612 23526 10640 25162
rect 10888 23866 10916 26726
rect 10980 26586 11008 29294
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 11072 27130 11100 28494
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 11164 26058 11192 29106
rect 11336 29028 11388 29034
rect 11336 28970 11388 28976
rect 11348 27946 11376 28970
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11428 28144 11480 28150
rect 11428 28086 11480 28092
rect 11336 27940 11388 27946
rect 11336 27882 11388 27888
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11256 27470 11284 27814
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 11072 26030 11192 26058
rect 11072 24614 11100 26030
rect 11152 25968 11204 25974
rect 11152 25910 11204 25916
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10612 23322 10640 23462
rect 10600 23316 10652 23322
rect 10600 23258 10652 23264
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 10416 22704 10468 22710
rect 10520 22681 10548 23054
rect 10416 22646 10468 22652
rect 10506 22672 10562 22681
rect 10324 22636 10376 22642
rect 10506 22607 10508 22616
rect 10324 22578 10376 22584
rect 10560 22607 10562 22616
rect 10508 22578 10560 22584
rect 10612 22545 10640 23258
rect 10598 22536 10654 22545
rect 10598 22471 10654 22480
rect 10796 22438 10824 23462
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10244 22066 10732 22094
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9770 21584 9826 21593
rect 9770 21519 9772 21528
rect 9824 21519 9826 21528
rect 9772 21490 9824 21496
rect 9876 21486 9904 21626
rect 9680 21480 9732 21486
rect 9678 21448 9680 21457
rect 9864 21480 9916 21486
rect 9732 21448 9734 21457
rect 9864 21422 9916 21428
rect 9678 21383 9734 21392
rect 10244 20942 10272 21966
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 9496 20868 9548 20874
rect 9496 20810 9548 20816
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9600 20618 9628 20742
rect 9600 20590 9720 20618
rect 9692 20534 9720 20590
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9678 20360 9734 20369
rect 9678 20295 9680 20304
rect 9732 20295 9734 20304
rect 9680 20266 9732 20272
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9508 18086 9536 19382
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9600 18290 9628 19246
rect 9784 19242 9812 20742
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9876 19786 9904 20538
rect 9968 20466 9996 20878
rect 9956 20460 10008 20466
rect 10232 20460 10284 20466
rect 10008 20420 10088 20448
rect 9956 20402 10008 20408
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9692 19145 9720 19178
rect 9876 19174 9904 19722
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9864 19168 9916 19174
rect 9678 19136 9734 19145
rect 9864 19110 9916 19116
rect 9678 19071 9734 19080
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9508 11778 9536 18022
rect 9600 11898 9628 18226
rect 9692 17066 9720 19071
rect 9968 18834 9996 19654
rect 10060 19310 10088 20420
rect 10232 20402 10284 20408
rect 10244 19854 10272 20402
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9876 17542 9904 18090
rect 9968 17882 9996 18770
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 10060 18465 10088 18634
rect 10046 18456 10102 18465
rect 10046 18391 10048 18400
rect 10100 18391 10102 18400
rect 10048 18362 10100 18368
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9876 16726 9904 17478
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 10336 11801 10364 21966
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10520 20942 10548 21286
rect 10612 21078 10640 21490
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10428 20505 10456 20742
rect 10414 20496 10470 20505
rect 10414 20431 10470 20440
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10612 20097 10640 20402
rect 10598 20088 10654 20097
rect 10598 20023 10654 20032
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 18465 10640 19790
rect 10598 18456 10654 18465
rect 10598 18391 10654 18400
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10428 17105 10456 17478
rect 10414 17096 10470 17105
rect 10414 17031 10470 17040
rect 10508 16992 10560 16998
rect 10506 16960 10508 16969
rect 10560 16960 10562 16969
rect 10506 16895 10562 16904
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 10322 11792 10378 11801
rect 9508 11750 9628 11778
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9508 8294 9536 10950
rect 9600 9042 9628 11750
rect 10322 11727 10378 11736
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 10336 8090 10364 10474
rect 10428 9450 10456 16662
rect 10704 12345 10732 22066
rect 10784 22092 10836 22098
rect 10888 22080 10916 22918
rect 10836 22052 10916 22080
rect 10784 22034 10836 22040
rect 10888 21554 10916 22052
rect 10876 21548 10928 21554
rect 10980 21536 11008 24006
rect 11072 23730 11100 24550
rect 11164 23798 11192 25910
rect 11244 25492 11296 25498
rect 11244 25434 11296 25440
rect 11152 23792 11204 23798
rect 11152 23734 11204 23740
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 11058 23352 11114 23361
rect 11058 23287 11114 23296
rect 11072 23254 11100 23287
rect 11060 23248 11112 23254
rect 11060 23190 11112 23196
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22166 11100 22374
rect 11164 22234 11192 23598
rect 11256 23118 11284 25434
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11242 22808 11298 22817
rect 11242 22743 11298 22752
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 11150 22128 11206 22137
rect 11150 22063 11206 22072
rect 11164 22030 11192 22063
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11256 21690 11284 22743
rect 11348 21962 11376 27882
rect 11440 25974 11468 28086
rect 11532 27169 11560 28358
rect 11624 27334 11652 32234
rect 11888 31952 11940 31958
rect 11888 31894 11940 31900
rect 11900 31754 11928 31894
rect 12084 31754 12112 33895
rect 12900 33312 12952 33318
rect 12900 33254 12952 33260
rect 12808 33176 12860 33182
rect 12808 33118 12860 33124
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 11716 31726 11928 31754
rect 11992 31726 12112 31754
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11518 27160 11574 27169
rect 11518 27095 11574 27104
rect 11716 27010 11744 31726
rect 11796 31136 11848 31142
rect 11848 31084 11928 31090
rect 11796 31078 11928 31084
rect 11808 31062 11928 31078
rect 11900 30870 11928 31062
rect 11888 30864 11940 30870
rect 11888 30806 11940 30812
rect 11796 30796 11848 30802
rect 11796 30738 11848 30744
rect 11808 28762 11836 30738
rect 11900 29170 11928 30806
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11796 28756 11848 28762
rect 11796 28698 11848 28704
rect 11992 28150 12020 31726
rect 12360 31686 12388 32166
rect 12473 32124 12781 32133
rect 12473 32122 12479 32124
rect 12535 32122 12559 32124
rect 12615 32122 12639 32124
rect 12695 32122 12719 32124
rect 12775 32122 12781 32124
rect 12535 32070 12537 32122
rect 12717 32070 12719 32122
rect 12473 32068 12479 32070
rect 12535 32068 12559 32070
rect 12615 32068 12639 32070
rect 12695 32068 12719 32070
rect 12775 32068 12781 32070
rect 12473 32059 12781 32068
rect 12348 31680 12400 31686
rect 12348 31622 12400 31628
rect 12348 31204 12400 31210
rect 12348 31146 12400 31152
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 12084 30258 12112 30670
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12072 29504 12124 29510
rect 12072 29446 12124 29452
rect 12084 29238 12112 29446
rect 12072 29232 12124 29238
rect 12072 29174 12124 29180
rect 12084 28762 12112 29174
rect 12072 28756 12124 28762
rect 12072 28698 12124 28704
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 12176 27962 12204 31078
rect 12256 30728 12308 30734
rect 12256 30670 12308 30676
rect 12268 29306 12296 30670
rect 12360 30598 12388 31146
rect 12820 31142 12848 33118
rect 12808 31136 12860 31142
rect 12808 31078 12860 31084
rect 12473 31036 12781 31045
rect 12473 31034 12479 31036
rect 12535 31034 12559 31036
rect 12615 31034 12639 31036
rect 12695 31034 12719 31036
rect 12775 31034 12781 31036
rect 12535 30982 12537 31034
rect 12717 30982 12719 31034
rect 12473 30980 12479 30982
rect 12535 30980 12559 30982
rect 12615 30980 12639 30982
rect 12695 30980 12719 30982
rect 12775 30980 12781 30982
rect 12473 30971 12781 30980
rect 12348 30592 12400 30598
rect 12348 30534 12400 30540
rect 12360 30326 12388 30534
rect 12820 30433 12848 31078
rect 12806 30424 12862 30433
rect 12806 30359 12862 30368
rect 12348 30320 12400 30326
rect 12348 30262 12400 30268
rect 12360 29578 12388 30262
rect 12808 30048 12860 30054
rect 12912 30036 12940 33254
rect 13004 32434 13032 34462
rect 14094 34350 14150 35150
rect 14830 34504 14886 34513
rect 14830 34439 14886 34448
rect 15290 34490 15346 35150
rect 15290 34462 15424 34490
rect 13266 34232 13322 34241
rect 13266 34167 13322 34176
rect 13176 33244 13228 33250
rect 13176 33186 13228 33192
rect 12992 32428 13044 32434
rect 12992 32370 13044 32376
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 13096 30802 13124 32166
rect 13188 31249 13216 33186
rect 13174 31240 13230 31249
rect 13174 31175 13230 31184
rect 13084 30796 13136 30802
rect 13084 30738 13136 30744
rect 13280 30054 13308 34167
rect 13636 32836 13688 32842
rect 13636 32778 13688 32784
rect 13544 32360 13596 32366
rect 13544 32302 13596 32308
rect 13556 31754 13584 32302
rect 13464 31726 13584 31754
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 13372 30433 13400 30602
rect 13358 30424 13414 30433
rect 13358 30359 13414 30368
rect 13358 30288 13414 30297
rect 13358 30223 13414 30232
rect 12860 30008 12940 30036
rect 12992 30048 13044 30054
rect 12808 29990 12860 29996
rect 12992 29990 13044 29996
rect 13268 30048 13320 30054
rect 13268 29990 13320 29996
rect 12473 29948 12781 29957
rect 12473 29946 12479 29948
rect 12535 29946 12559 29948
rect 12615 29946 12639 29948
rect 12695 29946 12719 29948
rect 12775 29946 12781 29948
rect 12535 29894 12537 29946
rect 12717 29894 12719 29946
rect 12473 29892 12479 29894
rect 12535 29892 12559 29894
rect 12615 29892 12639 29894
rect 12695 29892 12719 29894
rect 12775 29892 12781 29894
rect 12473 29883 12781 29892
rect 12820 29753 12848 29990
rect 12806 29744 12862 29753
rect 12806 29679 12862 29688
rect 12348 29572 12400 29578
rect 12348 29514 12400 29520
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 11992 27946 12204 27962
rect 11796 27940 11848 27946
rect 11796 27882 11848 27888
rect 11980 27940 12204 27946
rect 12032 27934 12204 27940
rect 11980 27882 12032 27888
rect 11808 27606 11836 27882
rect 12072 27872 12124 27878
rect 12072 27814 12124 27820
rect 11796 27600 11848 27606
rect 11796 27542 11848 27548
rect 12084 27402 12112 27814
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 12072 27396 12124 27402
rect 12072 27338 12124 27344
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11532 26982 11744 27010
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 11428 25968 11480 25974
rect 11428 25910 11480 25916
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 11440 24954 11468 25094
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11440 24177 11468 24890
rect 11426 24168 11482 24177
rect 11426 24103 11482 24112
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11440 23254 11468 23666
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11440 23118 11468 23190
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11428 22704 11480 22710
rect 11426 22672 11428 22681
rect 11480 22672 11482 22681
rect 11426 22607 11482 22616
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 10980 21508 11192 21536
rect 10876 21490 10928 21496
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10888 20777 10916 20878
rect 10874 20768 10930 20777
rect 10874 20703 10930 20712
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10888 19922 10916 20402
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10782 19544 10838 19553
rect 10782 19479 10838 19488
rect 10796 19174 10824 19479
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10888 18222 10916 19314
rect 10980 19281 11008 21354
rect 11164 20874 11192 21508
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11072 19961 11100 20742
rect 11152 20256 11204 20262
rect 11256 20233 11284 20742
rect 11348 20466 11376 21626
rect 11440 21622 11468 21898
rect 11428 21616 11480 21622
rect 11428 21558 11480 21564
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11440 20777 11468 20946
rect 11426 20768 11482 20777
rect 11426 20703 11482 20712
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11152 20198 11204 20204
rect 11242 20224 11298 20233
rect 11058 19952 11114 19961
rect 11058 19887 11114 19896
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10966 19272 11022 19281
rect 10966 19207 11022 19216
rect 11072 18834 11100 19314
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10980 18714 11008 18770
rect 10980 18686 11100 18714
rect 11164 18698 11192 20198
rect 11242 20159 11298 20168
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10888 16250 10916 18022
rect 10980 17338 11008 18566
rect 11072 18154 11100 18686
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11256 18290 11284 19654
rect 11348 19446 11376 20402
rect 11532 20074 11560 26982
rect 11612 26852 11664 26858
rect 11612 26794 11664 26800
rect 11624 26518 11652 26794
rect 11612 26512 11664 26518
rect 11612 26454 11664 26460
rect 11624 25498 11652 26454
rect 11808 26450 11836 26998
rect 11796 26444 11848 26450
rect 11796 26386 11848 26392
rect 11900 26194 11928 27270
rect 11980 26852 12032 26858
rect 11980 26794 12032 26800
rect 11716 26166 11928 26194
rect 11612 25492 11664 25498
rect 11612 25434 11664 25440
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11624 23497 11652 25298
rect 11716 24206 11744 26166
rect 11888 26036 11940 26042
rect 11888 25978 11940 25984
rect 11796 25764 11848 25770
rect 11796 25706 11848 25712
rect 11808 25294 11836 25706
rect 11900 25498 11928 25978
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11808 24410 11836 25094
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11610 23488 11666 23497
rect 11610 23423 11666 23432
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11624 22642 11652 23054
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11716 22681 11744 22918
rect 11702 22672 11758 22681
rect 11612 22636 11664 22642
rect 11702 22607 11758 22616
rect 11612 22578 11664 22584
rect 11624 22114 11652 22578
rect 11624 22086 11744 22114
rect 11532 20046 11652 20074
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 11532 19854 11560 19926
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11348 18766 11376 19246
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11440 18630 11468 19450
rect 11520 19440 11572 19446
rect 11520 19382 11572 19388
rect 11532 19174 11560 19382
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11532 18358 11560 18702
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11624 18193 11652 20046
rect 11716 19446 11744 22086
rect 11808 21622 11836 24346
rect 11900 24274 11928 24550
rect 11888 24268 11940 24274
rect 11888 24210 11940 24216
rect 11886 23896 11942 23905
rect 11886 23831 11942 23840
rect 11900 23032 11928 23831
rect 11992 23526 12020 26794
rect 12072 26308 12124 26314
rect 12072 26250 12124 26256
rect 12084 23769 12112 26250
rect 12176 25838 12204 27406
rect 12268 27305 12296 29242
rect 12473 28860 12781 28869
rect 12473 28858 12479 28860
rect 12535 28858 12559 28860
rect 12615 28858 12639 28860
rect 12695 28858 12719 28860
rect 12775 28858 12781 28860
rect 12535 28806 12537 28858
rect 12717 28806 12719 28858
rect 12473 28804 12479 28806
rect 12535 28804 12559 28806
rect 12615 28804 12639 28806
rect 12695 28804 12719 28806
rect 12775 28804 12781 28806
rect 12473 28795 12781 28804
rect 12440 28688 12492 28694
rect 12440 28630 12492 28636
rect 12452 27860 12480 28630
rect 12820 28150 12848 29242
rect 12898 29200 12954 29209
rect 12898 29135 12954 29144
rect 12808 28144 12860 28150
rect 12808 28086 12860 28092
rect 12820 27878 12848 28086
rect 12360 27832 12480 27860
rect 12808 27872 12860 27878
rect 12360 27554 12388 27832
rect 12808 27814 12860 27820
rect 12473 27772 12781 27781
rect 12473 27770 12479 27772
rect 12535 27770 12559 27772
rect 12615 27770 12639 27772
rect 12695 27770 12719 27772
rect 12775 27770 12781 27772
rect 12535 27718 12537 27770
rect 12717 27718 12719 27770
rect 12473 27716 12479 27718
rect 12535 27716 12559 27718
rect 12615 27716 12639 27718
rect 12695 27716 12719 27718
rect 12775 27716 12781 27718
rect 12473 27707 12781 27716
rect 12912 27606 12940 29135
rect 13004 27674 13032 29990
rect 13372 29850 13400 30223
rect 13360 29844 13412 29850
rect 13360 29786 13412 29792
rect 13084 29708 13136 29714
rect 13084 29650 13136 29656
rect 12992 27668 13044 27674
rect 12992 27610 13044 27616
rect 12900 27600 12952 27606
rect 12360 27526 12480 27554
rect 12900 27542 12952 27548
rect 12254 27296 12310 27305
rect 12254 27231 12310 27240
rect 12268 26586 12296 27231
rect 12452 26772 12480 27526
rect 13004 27112 13032 27610
rect 12360 26744 12480 26772
rect 12820 27084 13032 27112
rect 12360 26586 12388 26744
rect 12473 26684 12781 26693
rect 12473 26682 12479 26684
rect 12535 26682 12559 26684
rect 12615 26682 12639 26684
rect 12695 26682 12719 26684
rect 12775 26682 12781 26684
rect 12535 26630 12537 26682
rect 12717 26630 12719 26682
rect 12473 26628 12479 26630
rect 12535 26628 12559 26630
rect 12615 26628 12639 26630
rect 12695 26628 12719 26630
rect 12775 26628 12781 26630
rect 12473 26619 12781 26628
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12348 26580 12400 26586
rect 12820 26568 12848 27084
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12400 26540 12480 26568
rect 12348 26522 12400 26528
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 12164 25832 12216 25838
rect 12164 25774 12216 25780
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 25265 12204 25638
rect 12162 25256 12218 25265
rect 12162 25191 12218 25200
rect 12176 24954 12204 25191
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 12268 24614 12296 26386
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12360 26081 12388 26182
rect 12346 26072 12402 26081
rect 12346 26007 12402 26016
rect 12452 25684 12480 26540
rect 12728 26540 12848 26568
rect 12728 26246 12756 26540
rect 12806 26480 12862 26489
rect 12806 26415 12862 26424
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12360 25656 12480 25684
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12162 24304 12218 24313
rect 12162 24239 12218 24248
rect 12176 23866 12204 24239
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 12070 23760 12126 23769
rect 12070 23695 12126 23704
rect 12162 23624 12218 23633
rect 12162 23559 12218 23568
rect 12176 23526 12204 23559
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12176 23118 12204 23462
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 11900 23004 12020 23032
rect 11886 22944 11942 22953
rect 11886 22879 11942 22888
rect 11796 21616 11848 21622
rect 11796 21558 11848 21564
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 11808 20942 11836 21082
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11808 20466 11836 20742
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11808 19553 11836 20402
rect 11794 19544 11850 19553
rect 11794 19479 11850 19488
rect 11704 19440 11756 19446
rect 11704 19382 11756 19388
rect 11808 18873 11836 19479
rect 11794 18864 11850 18873
rect 11794 18799 11850 18808
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11610 18184 11666 18193
rect 11060 18148 11112 18154
rect 11610 18119 11666 18128
rect 11060 18090 11112 18096
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10980 16658 11008 17138
rect 11072 16794 11100 18090
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10888 15434 10916 16186
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10980 14618 11008 16594
rect 11256 16590 11284 18022
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11244 16584 11296 16590
rect 11150 16552 11206 16561
rect 11244 16526 11296 16532
rect 11150 16487 11206 16496
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10690 12336 10746 12345
rect 10690 12271 10746 12280
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 11164 7993 11192 16487
rect 11256 16182 11284 16526
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11256 15638 11284 16118
rect 11348 16114 11376 17138
rect 11532 17134 11560 17614
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11348 15706 11376 16050
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11348 15162 11376 15642
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11532 10742 11560 17070
rect 11624 16794 11652 17478
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11624 16153 11652 16594
rect 11610 16144 11666 16153
rect 11610 16079 11666 16088
rect 11808 15706 11836 18294
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11808 15502 11836 15642
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11900 12434 11928 22879
rect 11992 22778 12020 23004
rect 12072 22976 12124 22982
rect 12164 22976 12216 22982
rect 12072 22918 12124 22924
rect 12162 22944 12164 22953
rect 12216 22944 12218 22953
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11978 22264 12034 22273
rect 11978 22199 11980 22208
rect 12032 22199 12034 22208
rect 11980 22170 12032 22176
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11992 21010 12020 21626
rect 12084 21049 12112 22918
rect 12162 22879 12218 22888
rect 12162 22400 12218 22409
rect 12162 22335 12218 22344
rect 12176 21554 12204 22335
rect 12268 21962 12296 24006
rect 12360 23848 12388 25656
rect 12473 25596 12781 25605
rect 12473 25594 12479 25596
rect 12535 25594 12559 25596
rect 12615 25594 12639 25596
rect 12695 25594 12719 25596
rect 12775 25594 12781 25596
rect 12535 25542 12537 25594
rect 12717 25542 12719 25594
rect 12473 25540 12479 25542
rect 12535 25540 12559 25542
rect 12615 25540 12639 25542
rect 12695 25540 12719 25542
rect 12775 25540 12781 25542
rect 12473 25531 12781 25540
rect 12820 25430 12848 26415
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12912 25537 12940 26318
rect 12898 25528 12954 25537
rect 12898 25463 12954 25472
rect 12808 25424 12860 25430
rect 12808 25366 12860 25372
rect 12820 25106 12848 25366
rect 12900 25220 12952 25226
rect 12900 25162 12952 25168
rect 12728 25078 12848 25106
rect 12728 24818 12756 25078
rect 12806 24984 12862 24993
rect 12806 24919 12862 24928
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12820 24732 12848 24919
rect 12912 24886 12940 25162
rect 12900 24880 12952 24886
rect 12900 24822 12952 24828
rect 13004 24750 13032 26726
rect 13096 26586 13124 29650
rect 13372 29073 13400 29786
rect 13358 29064 13414 29073
rect 13358 28999 13414 29008
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 13084 25832 13136 25838
rect 13084 25774 13136 25780
rect 12900 24744 12952 24750
rect 12820 24704 12900 24732
rect 12900 24686 12952 24692
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 12473 24508 12781 24517
rect 12473 24506 12479 24508
rect 12535 24506 12559 24508
rect 12615 24506 12639 24508
rect 12695 24506 12719 24508
rect 12775 24506 12781 24508
rect 12535 24454 12537 24506
rect 12717 24454 12719 24506
rect 12473 24452 12479 24454
rect 12535 24452 12559 24454
rect 12615 24452 12639 24454
rect 12695 24452 12719 24454
rect 12775 24452 12781 24454
rect 12473 24443 12781 24452
rect 12438 24304 12494 24313
rect 12438 24239 12494 24248
rect 12452 24206 12480 24239
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12360 23820 12480 23848
rect 12346 23760 12402 23769
rect 12346 23695 12348 23704
rect 12400 23695 12402 23704
rect 12348 23666 12400 23672
rect 12452 23526 12480 23820
rect 12440 23520 12492 23526
rect 12346 23488 12402 23497
rect 12440 23462 12492 23468
rect 12346 23423 12402 23432
rect 12360 22778 12388 23423
rect 12473 23420 12781 23429
rect 12473 23418 12479 23420
rect 12535 23418 12559 23420
rect 12615 23418 12639 23420
rect 12695 23418 12719 23420
rect 12775 23418 12781 23420
rect 12535 23366 12537 23418
rect 12717 23366 12719 23418
rect 12473 23364 12479 23366
rect 12535 23364 12559 23366
rect 12615 23364 12639 23366
rect 12695 23364 12719 23366
rect 12775 23364 12781 23366
rect 12473 23355 12781 23364
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12452 22574 12480 23258
rect 12714 23216 12770 23225
rect 12714 23151 12770 23160
rect 12622 22944 12678 22953
rect 12728 22930 12756 23151
rect 12808 23112 12860 23118
rect 12806 23080 12808 23089
rect 12860 23080 12862 23089
rect 12806 23015 12862 23024
rect 12728 22902 12848 22930
rect 12622 22879 12678 22888
rect 12646 22794 12674 22879
rect 12646 22778 12756 22794
rect 12646 22772 12768 22778
rect 12646 22766 12716 22772
rect 12716 22714 12768 22720
rect 12820 22642 12848 22902
rect 12912 22778 12940 24686
rect 12990 23624 13046 23633
rect 12990 23559 13046 23568
rect 13004 23526 13032 23559
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12440 22568 12492 22574
rect 12912 22522 12940 22578
rect 12440 22510 12492 22516
rect 12728 22494 12940 22522
rect 12728 22438 12756 22494
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12716 22432 12768 22438
rect 13004 22386 13032 23122
rect 13096 22642 13124 25774
rect 13188 25294 13216 28494
rect 13268 28144 13320 28150
rect 13268 28086 13320 28092
rect 13280 27130 13308 28086
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13268 27124 13320 27130
rect 13268 27066 13320 27072
rect 13268 26580 13320 26586
rect 13268 26522 13320 26528
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13188 22760 13216 25094
rect 13280 24993 13308 26522
rect 13266 24984 13322 24993
rect 13372 24954 13400 28018
rect 13464 26790 13492 31726
rect 13542 31376 13598 31385
rect 13542 31311 13544 31320
rect 13596 31311 13598 31320
rect 13544 31282 13596 31288
rect 13648 30326 13676 32778
rect 14370 32328 14426 32337
rect 14844 32298 14872 34439
rect 15290 34350 15346 34462
rect 15396 32434 15424 34462
rect 16486 34350 16542 35150
rect 17314 34368 17370 34377
rect 16500 32858 16528 34350
rect 17682 34350 17738 35150
rect 18878 34350 18934 35150
rect 20074 34350 20130 35150
rect 21270 34350 21326 35150
rect 22466 34350 22522 35150
rect 23662 34350 23718 35150
rect 24858 34350 24914 35150
rect 25318 34640 25374 34649
rect 25318 34575 25374 34584
rect 24950 34504 25006 34513
rect 24950 34439 25006 34448
rect 17314 34303 17370 34312
rect 16500 32830 16712 32858
rect 16314 32668 16622 32677
rect 16314 32666 16320 32668
rect 16376 32666 16400 32668
rect 16456 32666 16480 32668
rect 16536 32666 16560 32668
rect 16616 32666 16622 32668
rect 16376 32614 16378 32666
rect 16558 32614 16560 32666
rect 16314 32612 16320 32614
rect 16376 32612 16400 32614
rect 16456 32612 16480 32614
rect 16536 32612 16560 32614
rect 16616 32612 16622 32614
rect 16314 32603 16622 32612
rect 16684 32434 16712 32830
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 14370 32263 14426 32272
rect 14832 32292 14884 32298
rect 14384 31754 14412 32263
rect 14832 32234 14884 32240
rect 14924 32292 14976 32298
rect 14924 32234 14976 32240
rect 16948 32292 17000 32298
rect 16948 32234 17000 32240
rect 14844 32026 14872 32234
rect 14832 32020 14884 32026
rect 14832 31962 14884 31968
rect 14740 31816 14792 31822
rect 14740 31758 14792 31764
rect 14292 31726 14412 31754
rect 14464 31748 14516 31754
rect 14004 31136 14056 31142
rect 14004 31078 14056 31084
rect 14016 30938 14044 31078
rect 14004 30932 14056 30938
rect 14004 30874 14056 30880
rect 13636 30320 13688 30326
rect 13636 30262 13688 30268
rect 13648 29306 13676 30262
rect 14096 30184 14148 30190
rect 14096 30126 14148 30132
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 13636 29300 13688 29306
rect 13636 29242 13688 29248
rect 13728 29232 13780 29238
rect 13728 29174 13780 29180
rect 13636 28960 13688 28966
rect 13636 28902 13688 28908
rect 13648 27606 13676 28902
rect 13636 27600 13688 27606
rect 13636 27542 13688 27548
rect 13544 27532 13596 27538
rect 13544 27474 13596 27480
rect 13452 26784 13504 26790
rect 13452 26726 13504 26732
rect 13464 25702 13492 26726
rect 13556 25906 13584 27474
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13648 26586 13676 26726
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13648 26081 13676 26182
rect 13634 26072 13690 26081
rect 13740 26042 13768 29174
rect 13818 28792 13874 28801
rect 13818 28727 13820 28736
rect 13872 28727 13874 28736
rect 13820 28698 13872 28704
rect 13912 28008 13964 28014
rect 13912 27950 13964 27956
rect 13818 27024 13874 27033
rect 13818 26959 13874 26968
rect 13634 26007 13690 26016
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13728 25900 13780 25906
rect 13728 25842 13780 25848
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 13266 24919 13322 24928
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13280 24313 13308 24754
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13266 24304 13322 24313
rect 13266 24239 13322 24248
rect 13372 24206 13400 24686
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13372 23662 13400 24006
rect 13464 23730 13492 25638
rect 13556 25276 13584 25842
rect 13634 25800 13690 25809
rect 13634 25735 13690 25744
rect 13648 25498 13676 25735
rect 13740 25537 13768 25842
rect 13726 25528 13782 25537
rect 13636 25492 13688 25498
rect 13726 25463 13782 25472
rect 13636 25434 13688 25440
rect 13636 25288 13688 25294
rect 13556 25248 13636 25276
rect 13556 24342 13584 25248
rect 13636 25230 13688 25236
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13544 24336 13596 24342
rect 13544 24278 13596 24284
rect 13542 24168 13598 24177
rect 13542 24103 13598 24112
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13360 23656 13412 23662
rect 13360 23598 13412 23604
rect 13556 23526 13584 24103
rect 13648 23526 13676 25094
rect 13740 24818 13768 25463
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13544 23520 13596 23526
rect 13266 23488 13322 23497
rect 13544 23462 13596 23468
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13266 23423 13322 23432
rect 13280 22982 13308 23423
rect 13556 23361 13584 23462
rect 13358 23352 13414 23361
rect 13358 23287 13414 23296
rect 13542 23352 13598 23361
rect 13542 23287 13598 23296
rect 13636 23316 13688 23322
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13187 22732 13216 22760
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 12716 22374 12768 22380
rect 12360 22098 12388 22374
rect 12820 22358 13032 22386
rect 12473 22332 12781 22341
rect 12473 22330 12479 22332
rect 12535 22330 12559 22332
rect 12615 22330 12639 22332
rect 12695 22330 12719 22332
rect 12775 22330 12781 22332
rect 12535 22278 12537 22330
rect 12717 22278 12719 22330
rect 12473 22276 12479 22278
rect 12535 22276 12559 22278
rect 12615 22276 12639 22278
rect 12695 22276 12719 22278
rect 12775 22276 12781 22278
rect 12473 22267 12781 22276
rect 12820 22216 12848 22358
rect 12728 22188 12848 22216
rect 12898 22264 12954 22273
rect 12898 22199 12954 22208
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12636 21865 12664 21966
rect 12622 21856 12678 21865
rect 12622 21791 12678 21800
rect 12254 21720 12310 21729
rect 12254 21655 12310 21664
rect 12438 21720 12494 21729
rect 12438 21655 12494 21664
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12268 21418 12296 21655
rect 12346 21448 12402 21457
rect 12256 21412 12308 21418
rect 12452 21434 12480 21655
rect 12728 21554 12756 22188
rect 12806 22128 12862 22137
rect 12806 22063 12862 22072
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12402 21406 12480 21434
rect 12530 21448 12586 21457
rect 12346 21383 12402 21392
rect 12530 21383 12532 21392
rect 12256 21354 12308 21360
rect 12584 21383 12586 21392
rect 12532 21354 12584 21360
rect 12473 21244 12781 21253
rect 12473 21242 12479 21244
rect 12535 21242 12559 21244
rect 12615 21242 12639 21244
rect 12695 21242 12719 21244
rect 12775 21242 12781 21244
rect 12535 21190 12537 21242
rect 12717 21190 12719 21242
rect 12473 21188 12479 21190
rect 12535 21188 12559 21190
rect 12615 21188 12639 21190
rect 12695 21188 12719 21190
rect 12775 21188 12781 21190
rect 12346 21176 12402 21185
rect 12473 21179 12781 21188
rect 12440 21140 12492 21146
rect 12402 21120 12440 21128
rect 12346 21111 12440 21120
rect 12360 21100 12440 21111
rect 12440 21082 12492 21088
rect 12070 21040 12126 21049
rect 11980 21004 12032 21010
rect 12070 20975 12126 20984
rect 11980 20946 12032 20952
rect 12072 20936 12124 20942
rect 12532 20936 12584 20942
rect 12072 20878 12124 20884
rect 12530 20904 12532 20913
rect 12584 20904 12586 20913
rect 12084 20777 12112 20878
rect 12530 20839 12586 20848
rect 12624 20800 12676 20806
rect 12070 20768 12126 20777
rect 12346 20768 12402 20777
rect 12070 20703 12126 20712
rect 12268 20726 12346 20754
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 11992 14521 12020 19926
rect 12084 19854 12112 20198
rect 12176 20058 12204 20334
rect 12268 20097 12296 20726
rect 12624 20742 12676 20748
rect 12346 20703 12402 20712
rect 12346 20632 12402 20641
rect 12346 20567 12402 20576
rect 12254 20088 12310 20097
rect 12164 20052 12216 20058
rect 12254 20023 12310 20032
rect 12164 19994 12216 20000
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12070 19680 12126 19689
rect 12070 19615 12126 19624
rect 12084 19446 12112 19615
rect 12176 19514 12204 19994
rect 12360 19922 12388 20567
rect 12532 20256 12584 20262
rect 12636 20244 12664 20742
rect 12820 20448 12848 22063
rect 12912 21894 12940 22199
rect 13096 22166 13124 22578
rect 13187 22556 13215 22732
rect 13372 22642 13400 23287
rect 13636 23258 13688 23264
rect 13450 23216 13506 23225
rect 13648 23202 13676 23258
rect 13740 23254 13768 24210
rect 13450 23151 13506 23160
rect 13556 23174 13676 23202
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 13464 23118 13492 23151
rect 13556 23118 13584 23174
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 13544 23112 13596 23118
rect 13832 23100 13860 26959
rect 13924 26217 13952 27950
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 13910 26208 13966 26217
rect 13910 26143 13966 26152
rect 13924 26042 13952 26143
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 13924 25430 13952 25774
rect 13912 25424 13964 25430
rect 13912 25366 13964 25372
rect 13910 24848 13966 24857
rect 13910 24783 13966 24792
rect 13924 24342 13952 24783
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 13912 24200 13964 24206
rect 13910 24168 13912 24177
rect 13964 24168 13966 24177
rect 14016 24138 14044 27338
rect 14108 25129 14136 30126
rect 14200 29782 14228 30126
rect 14188 29776 14240 29782
rect 14188 29718 14240 29724
rect 14200 29510 14228 29718
rect 14188 29504 14240 29510
rect 14188 29446 14240 29452
rect 14200 28966 14228 29446
rect 14188 28960 14240 28966
rect 14188 28902 14240 28908
rect 14200 28490 14228 28902
rect 14188 28484 14240 28490
rect 14188 28426 14240 28432
rect 14188 27464 14240 27470
rect 14186 27432 14188 27441
rect 14240 27432 14242 27441
rect 14186 27367 14242 27376
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14200 26761 14228 26862
rect 14186 26752 14242 26761
rect 14186 26687 14242 26696
rect 14094 25120 14150 25129
rect 14094 25055 14150 25064
rect 14108 24313 14136 25055
rect 14094 24304 14150 24313
rect 14094 24239 14150 24248
rect 13910 24103 13966 24112
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 13912 24064 13964 24070
rect 14096 24064 14148 24070
rect 13912 24006 13964 24012
rect 14002 24032 14058 24041
rect 13924 23526 13952 24006
rect 14096 24006 14148 24012
rect 14002 23967 14058 23976
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13910 23352 13966 23361
rect 13910 23287 13966 23296
rect 13924 23118 13952 23287
rect 13544 23054 13596 23060
rect 13648 23072 13860 23100
rect 13912 23112 13964 23118
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13187 22528 13216 22556
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 13004 21350 13032 21558
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13096 20806 13124 21966
rect 13188 21010 13216 22528
rect 13450 22536 13506 22545
rect 13268 22500 13320 22506
rect 13450 22471 13506 22480
rect 13268 22442 13320 22448
rect 13280 22409 13308 22442
rect 13266 22400 13322 22409
rect 13266 22335 13322 22344
rect 13464 22030 13492 22471
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13268 21888 13320 21894
rect 13556 21842 13584 22714
rect 13648 22098 13676 23072
rect 13912 23054 13964 23060
rect 13726 22944 13782 22953
rect 13726 22879 13782 22888
rect 13740 22273 13768 22879
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13726 22264 13782 22273
rect 13726 22199 13782 22208
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 13268 21830 13320 21836
rect 13280 21690 13308 21830
rect 13372 21814 13584 21842
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13372 21593 13400 21814
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13358 21584 13414 21593
rect 13358 21519 13414 21528
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13372 21146 13400 21286
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13464 21010 13492 21626
rect 13648 21185 13676 21830
rect 13634 21176 13690 21185
rect 13634 21111 13690 21120
rect 13176 21004 13228 21010
rect 13452 21004 13504 21010
rect 13176 20946 13228 20952
rect 13372 20964 13452 20992
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13266 20768 13322 20777
rect 13266 20703 13322 20712
rect 12898 20632 12954 20641
rect 12898 20567 12900 20576
rect 12952 20567 12954 20576
rect 12900 20538 12952 20544
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 12728 20420 12848 20448
rect 12728 20330 12756 20420
rect 12716 20324 12768 20330
rect 12716 20266 12768 20272
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 12584 20216 12664 20244
rect 12532 20198 12584 20204
rect 12473 20156 12781 20165
rect 12473 20154 12479 20156
rect 12535 20154 12559 20156
rect 12615 20154 12639 20156
rect 12695 20154 12719 20156
rect 12775 20154 12781 20156
rect 12535 20102 12537 20154
rect 12717 20102 12719 20154
rect 12473 20100 12479 20102
rect 12535 20100 12559 20102
rect 12615 20100 12639 20102
rect 12695 20100 12719 20102
rect 12775 20100 12781 20102
rect 12473 20091 12781 20100
rect 12820 19938 12848 20266
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12544 19910 12848 19938
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12176 18850 12204 19450
rect 12268 18970 12296 19790
rect 12544 19718 12572 19910
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12806 19816 12862 19825
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12530 19544 12586 19553
rect 12530 19479 12586 19488
rect 12544 19446 12572 19479
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12636 19378 12664 19790
rect 12716 19780 12768 19786
rect 12806 19751 12862 19760
rect 12716 19722 12768 19728
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12360 19145 12388 19314
rect 12728 19156 12756 19722
rect 12820 19718 12848 19751
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12912 19446 12940 20198
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 13004 19553 13032 19722
rect 12990 19544 13046 19553
rect 12990 19479 13046 19488
rect 12900 19440 12952 19446
rect 12806 19408 12862 19417
rect 12900 19382 12952 19388
rect 12806 19343 12808 19352
rect 12860 19343 12862 19352
rect 12808 19314 12860 19320
rect 12912 19310 12940 19382
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12346 19136 12402 19145
rect 12728 19128 12940 19156
rect 12346 19071 12402 19080
rect 12473 19068 12781 19077
rect 12473 19066 12479 19068
rect 12535 19066 12559 19068
rect 12615 19066 12639 19068
rect 12695 19066 12719 19068
rect 12775 19066 12781 19068
rect 12535 19014 12537 19066
rect 12717 19014 12719 19066
rect 12473 19012 12479 19014
rect 12535 19012 12559 19014
rect 12615 19012 12639 19014
rect 12695 19012 12719 19014
rect 12775 19012 12781 19014
rect 12473 19003 12781 19012
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12624 18896 12676 18902
rect 12176 18822 12296 18850
rect 12624 18838 12676 18844
rect 12268 18766 12296 18822
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 14929 12112 18566
rect 12176 18170 12204 18702
rect 12636 18222 12664 18838
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 18290 12848 18566
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12624 18216 12676 18222
rect 12176 18154 12296 18170
rect 12624 18158 12676 18164
rect 12176 18148 12308 18154
rect 12176 18142 12256 18148
rect 12256 18090 12308 18096
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17678 12204 18022
rect 12473 17980 12781 17989
rect 12473 17978 12479 17980
rect 12535 17978 12559 17980
rect 12615 17978 12639 17980
rect 12695 17978 12719 17980
rect 12775 17978 12781 17980
rect 12535 17926 12537 17978
rect 12717 17926 12719 17978
rect 12473 17924 12479 17926
rect 12535 17924 12559 17926
rect 12615 17924 12639 17926
rect 12695 17924 12719 17926
rect 12775 17924 12781 17926
rect 12473 17915 12781 17924
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12912 17513 12940 19128
rect 13004 18766 13032 19479
rect 13096 19378 13124 20470
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13188 19446 13216 19926
rect 13280 19854 13308 20703
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13176 19440 13228 19446
rect 13280 19417 13308 19450
rect 13176 19382 13228 19388
rect 13266 19408 13322 19417
rect 13084 19372 13136 19378
rect 13266 19343 13322 19352
rect 13084 19314 13136 19320
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13188 18329 13216 19246
rect 13372 19174 13400 20964
rect 13452 20946 13504 20952
rect 13636 20800 13688 20806
rect 13450 20768 13506 20777
rect 13636 20742 13688 20748
rect 13450 20703 13506 20712
rect 13464 20534 13492 20703
rect 13542 20632 13598 20641
rect 13542 20567 13598 20576
rect 13648 20584 13676 20742
rect 13556 20534 13584 20567
rect 13648 20556 13768 20584
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13740 20398 13768 20556
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13464 19553 13492 19790
rect 13450 19544 13506 19553
rect 13450 19479 13506 19488
rect 13450 19272 13506 19281
rect 13450 19207 13506 19216
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13280 18834 13308 19110
rect 13464 18902 13492 19207
rect 13556 18902 13584 20334
rect 13832 20097 13860 22578
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 21486 13952 22510
rect 14016 21622 14044 23967
rect 14108 23798 14136 24006
rect 14096 23792 14148 23798
rect 14096 23734 14148 23740
rect 14200 23526 14228 26687
rect 14292 25702 14320 31726
rect 14464 31690 14516 31696
rect 14476 30054 14504 31690
rect 14648 31680 14700 31686
rect 14648 31622 14700 31628
rect 14660 30598 14688 31622
rect 14752 31414 14780 31758
rect 14740 31408 14792 31414
rect 14740 31350 14792 31356
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 14740 31136 14792 31142
rect 14738 31104 14740 31113
rect 14792 31104 14794 31113
rect 14738 31039 14794 31048
rect 14648 30592 14700 30598
rect 14648 30534 14700 30540
rect 14660 30394 14688 30534
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14372 30048 14424 30054
rect 14372 29990 14424 29996
rect 14464 30048 14516 30054
rect 14516 30008 14596 30036
rect 14464 29990 14516 29996
rect 14384 29850 14412 29990
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14384 29345 14412 29786
rect 14370 29336 14426 29345
rect 14370 29271 14426 29280
rect 14372 29096 14424 29102
rect 14372 29038 14424 29044
rect 14462 29064 14518 29073
rect 14384 28014 14412 29038
rect 14462 28999 14518 29008
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14372 27668 14424 27674
rect 14372 27610 14424 27616
rect 14384 25770 14412 27610
rect 14476 26314 14504 28999
rect 14568 28218 14596 30008
rect 14660 29714 14688 30330
rect 14648 29708 14700 29714
rect 14648 29650 14700 29656
rect 14556 28212 14608 28218
rect 14556 28154 14608 28160
rect 14568 28121 14596 28154
rect 14554 28112 14610 28121
rect 14554 28047 14610 28056
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14462 25936 14518 25945
rect 14462 25871 14518 25880
rect 14372 25764 14424 25770
rect 14372 25706 14424 25712
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14292 25537 14320 25638
rect 14278 25528 14334 25537
rect 14278 25463 14334 25472
rect 14280 25424 14332 25430
rect 14280 25366 14332 25372
rect 14292 24818 14320 25366
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14384 24138 14412 25706
rect 14476 25498 14504 25871
rect 14464 25492 14516 25498
rect 14464 25434 14516 25440
rect 14464 25288 14516 25294
rect 14462 25256 14464 25265
rect 14516 25256 14518 25265
rect 14462 25191 14518 25200
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14292 23798 14320 24074
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14280 23588 14332 23594
rect 14280 23530 14332 23536
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14108 23361 14136 23462
rect 14094 23352 14150 23361
rect 14094 23287 14150 23296
rect 14188 23248 14240 23254
rect 14188 23190 14240 23196
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22778 14136 22918
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 14108 22234 14136 22510
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 14200 21894 14228 23190
rect 14292 22234 14320 23530
rect 14384 23322 14412 23666
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14384 22137 14412 23054
rect 14476 22234 14504 24550
rect 14568 23905 14596 27950
rect 14660 26586 14688 29650
rect 14752 29034 14780 31039
rect 14844 29578 14872 31282
rect 14936 30977 14964 32234
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 16028 32224 16080 32230
rect 16028 32166 16080 32172
rect 14922 30968 14978 30977
rect 14922 30903 14978 30912
rect 14924 30388 14976 30394
rect 14924 30330 14976 30336
rect 14832 29572 14884 29578
rect 14832 29514 14884 29520
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14752 28218 14780 28970
rect 14740 28212 14792 28218
rect 14740 28154 14792 28160
rect 14648 26580 14700 26586
rect 14648 26522 14700 26528
rect 14648 25696 14700 25702
rect 14648 25638 14700 25644
rect 14660 24177 14688 25638
rect 14752 25537 14780 28154
rect 14844 27402 14872 29514
rect 14936 28150 14964 30330
rect 15120 30190 15148 32166
rect 15936 31884 15988 31890
rect 15936 31826 15988 31832
rect 15844 31816 15896 31822
rect 15844 31758 15896 31764
rect 15660 31748 15712 31754
rect 15660 31690 15712 31696
rect 15568 31136 15620 31142
rect 15568 31078 15620 31084
rect 15580 30734 15608 31078
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15108 30184 15160 30190
rect 15476 30184 15528 30190
rect 15108 30126 15160 30132
rect 15382 30152 15438 30161
rect 15476 30126 15528 30132
rect 15382 30087 15438 30096
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 14924 28144 14976 28150
rect 14924 28086 14976 28092
rect 14922 27432 14978 27441
rect 14832 27396 14884 27402
rect 14922 27367 14978 27376
rect 14832 27338 14884 27344
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14738 25528 14794 25537
rect 14738 25463 14794 25472
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14752 24954 14780 25298
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14844 24886 14872 25842
rect 14936 25106 14964 27367
rect 15028 25906 15056 29446
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15108 27872 15160 27878
rect 15108 27814 15160 27820
rect 15120 26790 15148 27814
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15106 26344 15162 26353
rect 15106 26279 15108 26288
rect 15160 26279 15162 26288
rect 15108 26250 15160 26256
rect 15212 26194 15240 28358
rect 15304 27946 15332 28358
rect 15396 28218 15424 30087
rect 15488 29306 15516 30126
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15580 29238 15608 30670
rect 15672 30598 15700 31690
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15752 30592 15804 30598
rect 15752 30534 15804 30540
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15568 29028 15620 29034
rect 15568 28970 15620 28976
rect 15474 28656 15530 28665
rect 15474 28591 15530 28600
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 15292 27940 15344 27946
rect 15292 27882 15344 27888
rect 15304 27130 15332 27882
rect 15396 27674 15424 28154
rect 15384 27668 15436 27674
rect 15384 27610 15436 27616
rect 15382 27568 15438 27577
rect 15382 27503 15438 27512
rect 15292 27124 15344 27130
rect 15292 27066 15344 27072
rect 15396 26858 15424 27503
rect 15384 26852 15436 26858
rect 15384 26794 15436 26800
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15304 26602 15332 26726
rect 15304 26574 15424 26602
rect 15292 26512 15344 26518
rect 15292 26454 15344 26460
rect 15120 26166 15240 26194
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 14936 25078 15056 25106
rect 14922 24984 14978 24993
rect 14922 24919 14978 24928
rect 14832 24880 14884 24886
rect 14738 24848 14794 24857
rect 14832 24822 14884 24828
rect 14738 24783 14794 24792
rect 14752 24682 14780 24783
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14830 24576 14886 24585
rect 14830 24511 14886 24520
rect 14738 24440 14794 24449
rect 14738 24375 14740 24384
rect 14792 24375 14794 24384
rect 14740 24346 14792 24352
rect 14646 24168 14702 24177
rect 14646 24103 14702 24112
rect 14554 23896 14610 23905
rect 14554 23831 14610 23840
rect 14568 23798 14596 23831
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14660 23338 14688 24103
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14568 23310 14688 23338
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14370 22128 14426 22137
rect 14370 22063 14426 22072
rect 14568 21962 14596 23310
rect 14648 23112 14700 23118
rect 14752 23100 14780 23598
rect 14844 23594 14872 24511
rect 14936 24052 14964 24919
rect 15028 24410 15056 25078
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 15016 24064 15068 24070
rect 14936 24024 15016 24052
rect 15016 24006 15068 24012
rect 14922 23760 14978 23769
rect 15120 23730 15148 26166
rect 15304 26081 15332 26454
rect 15290 26072 15346 26081
rect 15290 26007 15346 26016
rect 15290 25936 15346 25945
rect 15290 25871 15292 25880
rect 15344 25871 15346 25880
rect 15292 25842 15344 25848
rect 15200 25492 15252 25498
rect 15252 25452 15332 25480
rect 15200 25434 15252 25440
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 14922 23695 14978 23704
rect 15108 23724 15160 23730
rect 14832 23588 14884 23594
rect 14832 23530 14884 23536
rect 14936 23497 14964 23695
rect 15108 23666 15160 23672
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 14922 23488 14978 23497
rect 14922 23423 14978 23432
rect 14830 23352 14886 23361
rect 14830 23287 14832 23296
rect 14884 23287 14886 23296
rect 14924 23316 14976 23322
rect 14832 23258 14884 23264
rect 14924 23258 14976 23264
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 14700 23072 14780 23100
rect 14648 23054 14700 23060
rect 14646 22808 14702 22817
rect 14646 22743 14702 22752
rect 14660 22710 14688 22743
rect 14648 22704 14700 22710
rect 14648 22646 14700 22652
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14646 21856 14702 21865
rect 14646 21791 14702 21800
rect 14186 21720 14242 21729
rect 14186 21655 14242 21664
rect 14004 21616 14056 21622
rect 14004 21558 14056 21564
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13818 20088 13874 20097
rect 13728 20052 13780 20058
rect 13924 20058 13952 20198
rect 13818 20023 13874 20032
rect 13912 20052 13964 20058
rect 13728 19994 13780 20000
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13648 19718 13676 19858
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13740 19446 13768 19994
rect 13832 19922 13860 20023
rect 13912 19994 13964 20000
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 14016 19689 14044 20538
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14108 20262 14136 20402
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14002 19680 14058 19689
rect 14002 19615 14058 19624
rect 14108 19514 14136 20198
rect 14200 19718 14228 21655
rect 14462 21584 14518 21593
rect 14462 21519 14518 21528
rect 14476 21010 14504 21519
rect 14660 21486 14688 21791
rect 14648 21480 14700 21486
rect 14752 21457 14780 23072
rect 14648 21422 14700 21428
rect 14738 21448 14794 21457
rect 14738 21383 14794 21392
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14476 20806 14504 20946
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14292 19990 14320 20402
rect 14752 20398 14780 20742
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19718 14320 19790
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13450 18728 13506 18737
rect 13372 18686 13450 18714
rect 13174 18320 13230 18329
rect 13174 18255 13230 18264
rect 13266 17912 13322 17921
rect 13266 17847 13322 17856
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13004 17542 13032 17682
rect 13280 17542 13308 17847
rect 12992 17536 13044 17542
rect 12898 17504 12954 17513
rect 13268 17536 13320 17542
rect 12992 17478 13044 17484
rect 13188 17496 13268 17524
rect 12898 17439 12954 17448
rect 12622 17368 12678 17377
rect 12622 17303 12678 17312
rect 13082 17368 13138 17377
rect 13082 17303 13138 17312
rect 12636 17202 12664 17303
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16658 12204 16934
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12162 16552 12218 16561
rect 12162 16487 12218 16496
rect 12176 15314 12204 16487
rect 12268 15473 12296 17002
rect 12360 16250 12388 17138
rect 12473 16892 12781 16901
rect 12473 16890 12479 16892
rect 12535 16890 12559 16892
rect 12615 16890 12639 16892
rect 12695 16890 12719 16892
rect 12775 16890 12781 16892
rect 12535 16838 12537 16890
rect 12717 16838 12719 16890
rect 12473 16836 12479 16838
rect 12535 16836 12559 16838
rect 12615 16836 12639 16838
rect 12695 16836 12719 16838
rect 12775 16836 12781 16838
rect 12473 16827 12781 16836
rect 12714 16688 12770 16697
rect 12714 16623 12770 16632
rect 12728 16522 12756 16623
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12636 16425 12664 16458
rect 12622 16416 12678 16425
rect 12622 16351 12678 16360
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12254 15464 12310 15473
rect 12254 15399 12310 15408
rect 12176 15286 12296 15314
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12070 14920 12126 14929
rect 12070 14855 12126 14864
rect 12176 14550 12204 15098
rect 12164 14544 12216 14550
rect 11978 14512 12034 14521
rect 12164 14486 12216 14492
rect 11978 14447 12034 14456
rect 12268 12434 12296 15286
rect 12360 15094 12388 16186
rect 12473 15804 12781 15813
rect 12473 15802 12479 15804
rect 12535 15802 12559 15804
rect 12615 15802 12639 15804
rect 12695 15802 12719 15804
rect 12775 15802 12781 15804
rect 12535 15750 12537 15802
rect 12717 15750 12719 15802
rect 12473 15748 12479 15750
rect 12535 15748 12559 15750
rect 12615 15748 12639 15750
rect 12695 15748 12719 15750
rect 12775 15748 12781 15750
rect 12473 15739 12781 15748
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12473 14716 12781 14725
rect 12473 14714 12479 14716
rect 12535 14714 12559 14716
rect 12615 14714 12639 14716
rect 12695 14714 12719 14716
rect 12775 14714 12781 14716
rect 12535 14662 12537 14714
rect 12717 14662 12719 14714
rect 12473 14660 12479 14662
rect 12535 14660 12559 14662
rect 12615 14660 12639 14662
rect 12695 14660 12719 14662
rect 12775 14660 12781 14662
rect 12473 14651 12781 14660
rect 12473 13628 12781 13637
rect 12473 13626 12479 13628
rect 12535 13626 12559 13628
rect 12615 13626 12639 13628
rect 12695 13626 12719 13628
rect 12775 13626 12781 13628
rect 12535 13574 12537 13626
rect 12717 13574 12719 13626
rect 12473 13572 12479 13574
rect 12535 13572 12559 13574
rect 12615 13572 12639 13574
rect 12695 13572 12719 13574
rect 12775 13572 12781 13574
rect 12473 13563 12781 13572
rect 12912 12889 12940 17206
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13004 16561 13032 16662
rect 12990 16552 13046 16561
rect 12990 16487 13046 16496
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16114 13032 16390
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13096 15570 13124 17303
rect 13188 17270 13216 17496
rect 13268 17478 13320 17484
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13096 15434 13124 15506
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12898 12880 12954 12889
rect 12898 12815 12954 12824
rect 12473 12540 12781 12549
rect 12473 12538 12479 12540
rect 12535 12538 12559 12540
rect 12615 12538 12639 12540
rect 12695 12538 12719 12540
rect 12775 12538 12781 12540
rect 12535 12486 12537 12538
rect 12717 12486 12719 12538
rect 12473 12484 12479 12486
rect 12535 12484 12559 12486
rect 12615 12484 12639 12486
rect 12695 12484 12719 12486
rect 12775 12484 12781 12486
rect 12473 12475 12781 12484
rect 11900 12406 12112 12434
rect 12268 12406 12388 12434
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11150 7984 11206 7993
rect 11150 7919 11206 7928
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8632 7644 8940 7653
rect 8632 7642 8638 7644
rect 8694 7642 8718 7644
rect 8774 7642 8798 7644
rect 8854 7642 8878 7644
rect 8934 7642 8940 7644
rect 8694 7590 8696 7642
rect 8876 7590 8878 7642
rect 8632 7588 8638 7590
rect 8694 7588 8718 7590
rect 8774 7588 8798 7590
rect 8854 7588 8878 7590
rect 8934 7588 8940 7590
rect 8632 7579 8940 7588
rect 12084 6914 12112 12406
rect 12360 9654 12388 12406
rect 13004 11529 13032 15302
rect 13096 14482 13124 15370
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13096 14074 13124 14418
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13188 11665 13216 17002
rect 13280 15722 13308 17206
rect 13372 16590 13400 18686
rect 13450 18663 13506 18672
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13450 17640 13506 17649
rect 13450 17575 13452 17584
rect 13504 17575 13506 17584
rect 13452 17546 13504 17552
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16114 13400 16390
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13360 15904 13412 15910
rect 13358 15872 13360 15881
rect 13412 15872 13414 15881
rect 13358 15807 13414 15816
rect 13280 15694 13400 15722
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 13870 13308 15438
rect 13372 14278 13400 15694
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13174 11656 13230 11665
rect 13174 11591 13230 11600
rect 12990 11520 13046 11529
rect 12473 11452 12781 11461
rect 12990 11455 13046 11464
rect 12473 11450 12479 11452
rect 12535 11450 12559 11452
rect 12615 11450 12639 11452
rect 12695 11450 12719 11452
rect 12775 11450 12781 11452
rect 12535 11398 12537 11450
rect 12717 11398 12719 11450
rect 12473 11396 12479 11398
rect 12535 11396 12559 11398
rect 12615 11396 12639 11398
rect 12695 11396 12719 11398
rect 12775 11396 12781 11398
rect 12473 11387 12781 11396
rect 12473 10364 12781 10373
rect 12473 10362 12479 10364
rect 12535 10362 12559 10364
rect 12615 10362 12639 10364
rect 12695 10362 12719 10364
rect 12775 10362 12781 10364
rect 12535 10310 12537 10362
rect 12717 10310 12719 10362
rect 12473 10308 12479 10310
rect 12535 10308 12559 10310
rect 12615 10308 12639 10310
rect 12695 10308 12719 10310
rect 12775 10308 12781 10310
rect 12473 10299 12781 10308
rect 13280 10062 13308 13806
rect 13372 12434 13400 14010
rect 13464 13705 13492 16730
rect 13450 13696 13506 13705
rect 13450 13631 13506 13640
rect 13372 12406 13492 12434
rect 13464 11082 13492 12406
rect 13556 12306 13584 18566
rect 13648 18290 13676 19314
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13740 19145 13768 19178
rect 13726 19136 13782 19145
rect 13726 19071 13782 19080
rect 13728 18964 13780 18970
rect 13924 18952 13952 19246
rect 14292 18970 14320 19314
rect 14476 19009 14504 20198
rect 14660 19786 14688 20266
rect 14844 20262 14872 23122
rect 14936 21690 14964 23258
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 15028 22506 15056 22646
rect 15120 22642 15148 23530
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15016 22500 15068 22506
rect 15016 22442 15068 22448
rect 15120 22148 15148 22578
rect 15028 22120 15148 22148
rect 14924 21684 14976 21690
rect 14924 21626 14976 21632
rect 15028 21078 15056 22120
rect 15212 22080 15240 25094
rect 15304 23905 15332 25452
rect 15396 24886 15424 26574
rect 15384 24880 15436 24886
rect 15384 24822 15436 24828
rect 15384 24744 15436 24750
rect 15382 24712 15384 24721
rect 15436 24712 15438 24721
rect 15382 24647 15438 24656
rect 15382 24576 15438 24585
rect 15382 24511 15438 24520
rect 15290 23896 15346 23905
rect 15396 23866 15424 24511
rect 15488 24018 15516 28591
rect 15580 25945 15608 28970
rect 15672 27878 15700 30534
rect 15764 29209 15792 30534
rect 15856 30161 15884 31758
rect 15842 30152 15898 30161
rect 15842 30087 15898 30096
rect 15750 29200 15806 29209
rect 15750 29135 15806 29144
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 15752 28960 15804 28966
rect 15752 28902 15804 28908
rect 15764 28490 15792 28902
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15764 27946 15792 28426
rect 15752 27940 15804 27946
rect 15752 27882 15804 27888
rect 15660 27872 15712 27878
rect 15660 27814 15712 27820
rect 15752 27668 15804 27674
rect 15752 27610 15804 27616
rect 15764 27577 15792 27610
rect 15750 27568 15806 27577
rect 15750 27503 15806 27512
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15672 27305 15700 27338
rect 15658 27296 15714 27305
rect 15658 27231 15714 27240
rect 15672 27130 15700 27231
rect 15660 27124 15712 27130
rect 15712 27084 15792 27112
rect 15660 27066 15712 27072
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 15566 25936 15622 25945
rect 15566 25871 15622 25880
rect 15580 25294 15608 25871
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15672 25158 15700 26250
rect 15764 26194 15792 27084
rect 15856 26314 15884 29106
rect 15948 28257 15976 31826
rect 16040 30410 16068 32166
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16212 31680 16264 31686
rect 16212 31622 16264 31628
rect 16118 31240 16174 31249
rect 16224 31210 16252 31622
rect 16314 31580 16622 31589
rect 16314 31578 16320 31580
rect 16376 31578 16400 31580
rect 16456 31578 16480 31580
rect 16536 31578 16560 31580
rect 16616 31578 16622 31580
rect 16376 31526 16378 31578
rect 16558 31526 16560 31578
rect 16314 31524 16320 31526
rect 16376 31524 16400 31526
rect 16456 31524 16480 31526
rect 16536 31524 16560 31526
rect 16616 31524 16622 31526
rect 16314 31515 16622 31524
rect 16118 31175 16174 31184
rect 16212 31204 16264 31210
rect 16132 30938 16160 31175
rect 16212 31146 16264 31152
rect 16224 30977 16252 31146
rect 16210 30968 16266 30977
rect 16120 30932 16172 30938
rect 16210 30903 16266 30912
rect 16120 30874 16172 30880
rect 16132 30569 16160 30874
rect 16118 30560 16174 30569
rect 16118 30495 16174 30504
rect 16314 30492 16622 30501
rect 16314 30490 16320 30492
rect 16376 30490 16400 30492
rect 16456 30490 16480 30492
rect 16536 30490 16560 30492
rect 16616 30490 16622 30492
rect 16376 30438 16378 30490
rect 16558 30438 16560 30490
rect 16314 30436 16320 30438
rect 16376 30436 16400 30438
rect 16456 30436 16480 30438
rect 16536 30436 16560 30438
rect 16616 30436 16622 30438
rect 16314 30427 16622 30436
rect 16040 30382 16252 30410
rect 16120 30320 16172 30326
rect 16120 30262 16172 30268
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 16040 29510 16068 29990
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16040 29306 16068 29446
rect 16028 29300 16080 29306
rect 16028 29242 16080 29248
rect 16040 28762 16068 29242
rect 16028 28756 16080 28762
rect 16028 28698 16080 28704
rect 15934 28248 15990 28257
rect 15934 28183 15936 28192
rect 15988 28183 15990 28192
rect 15936 28154 15988 28160
rect 15948 28123 15976 28154
rect 15934 27568 15990 27577
rect 16132 27554 16160 30262
rect 16224 29782 16252 30382
rect 16212 29776 16264 29782
rect 16212 29718 16264 29724
rect 16314 29404 16622 29413
rect 16314 29402 16320 29404
rect 16376 29402 16400 29404
rect 16456 29402 16480 29404
rect 16536 29402 16560 29404
rect 16616 29402 16622 29404
rect 16376 29350 16378 29402
rect 16558 29350 16560 29402
rect 16314 29348 16320 29350
rect 16376 29348 16400 29350
rect 16456 29348 16480 29350
rect 16536 29348 16560 29350
rect 16616 29348 16622 29350
rect 16314 29339 16622 29348
rect 16210 29064 16266 29073
rect 16210 28999 16212 29008
rect 16264 28999 16266 29008
rect 16212 28970 16264 28976
rect 16684 28540 16712 31758
rect 16960 31482 16988 32234
rect 16764 31476 16816 31482
rect 16764 31418 16816 31424
rect 16948 31476 17000 31482
rect 16948 31418 17000 31424
rect 16776 29345 16804 31418
rect 17040 31408 17092 31414
rect 17040 31350 17092 31356
rect 16854 30560 16910 30569
rect 17052 30546 17080 31350
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17236 30938 17264 31078
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17236 30841 17264 30874
rect 17222 30832 17278 30841
rect 17222 30767 17278 30776
rect 17130 30696 17186 30705
rect 17130 30631 17132 30640
rect 17184 30631 17186 30640
rect 17132 30602 17184 30608
rect 17052 30518 17264 30546
rect 16854 30495 16910 30504
rect 16868 29850 16896 30495
rect 16856 29844 16908 29850
rect 16856 29786 16908 29792
rect 16948 29844 17000 29850
rect 16948 29786 17000 29792
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16762 29336 16818 29345
rect 16762 29271 16818 29280
rect 16776 29102 16804 29271
rect 16764 29096 16816 29102
rect 16764 29038 16816 29044
rect 16684 28512 16804 28540
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16314 28316 16622 28325
rect 16314 28314 16320 28316
rect 16376 28314 16400 28316
rect 16456 28314 16480 28316
rect 16536 28314 16560 28316
rect 16616 28314 16622 28316
rect 16376 28262 16378 28314
rect 16558 28262 16560 28314
rect 16314 28260 16320 28262
rect 16376 28260 16400 28262
rect 16456 28260 16480 28262
rect 16536 28260 16560 28262
rect 16616 28260 16622 28262
rect 16314 28251 16622 28260
rect 16580 28144 16632 28150
rect 16580 28086 16632 28092
rect 16592 27674 16620 28086
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 15934 27503 15990 27512
rect 16040 27526 16160 27554
rect 16210 27568 16266 27577
rect 15948 26382 15976 27503
rect 16040 27062 16068 27526
rect 16210 27503 16266 27512
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 16028 27056 16080 27062
rect 16028 26998 16080 27004
rect 16026 26616 16082 26625
rect 16026 26551 16082 26560
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 15934 26208 15990 26217
rect 15764 26166 15884 26194
rect 15750 26072 15806 26081
rect 15750 26007 15806 26016
rect 15660 25152 15712 25158
rect 15580 25112 15660 25140
rect 15580 24818 15608 25112
rect 15660 25094 15712 25100
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15566 24440 15622 24449
rect 15566 24375 15622 24384
rect 15580 24138 15608 24375
rect 15672 24138 15700 24890
rect 15764 24410 15792 26007
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15750 24304 15806 24313
rect 15750 24239 15806 24248
rect 15568 24132 15620 24138
rect 15568 24074 15620 24080
rect 15660 24132 15712 24138
rect 15660 24074 15712 24080
rect 15764 24018 15792 24239
rect 15488 23990 15608 24018
rect 15290 23831 15346 23840
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15304 23322 15332 23530
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 15384 23248 15436 23254
rect 15384 23190 15436 23196
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 15120 22052 15240 22080
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 15014 20904 15070 20913
rect 15014 20839 15070 20848
rect 15028 20262 15056 20839
rect 15120 20714 15148 22052
rect 15304 22001 15332 22986
rect 15290 21992 15346 22001
rect 15200 21956 15252 21962
rect 15396 21962 15424 23190
rect 15488 22710 15516 23802
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15580 22574 15608 23990
rect 15672 23990 15792 24018
rect 15672 23798 15700 23990
rect 15660 23792 15712 23798
rect 15660 23734 15712 23740
rect 15750 23760 15806 23769
rect 15672 23118 15700 23734
rect 15856 23730 15884 26166
rect 15934 26143 15990 26152
rect 15948 25537 15976 26143
rect 15934 25528 15990 25537
rect 15934 25463 15990 25472
rect 15936 25424 15988 25430
rect 15936 25366 15988 25372
rect 15948 25265 15976 25366
rect 15934 25256 15990 25265
rect 15934 25191 15990 25200
rect 15934 25120 15990 25129
rect 15934 25055 15990 25064
rect 15948 24886 15976 25055
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 15934 24712 15990 24721
rect 16040 24698 16068 26551
rect 16132 25276 16160 27406
rect 16224 26858 16252 27503
rect 16314 27228 16622 27237
rect 16314 27226 16320 27228
rect 16376 27226 16400 27228
rect 16456 27226 16480 27228
rect 16536 27226 16560 27228
rect 16616 27226 16622 27228
rect 16376 27174 16378 27226
rect 16558 27174 16560 27226
rect 16314 27172 16320 27174
rect 16376 27172 16400 27174
rect 16456 27172 16480 27174
rect 16536 27172 16560 27174
rect 16616 27172 16622 27174
rect 16314 27163 16622 27172
rect 16488 27056 16540 27062
rect 16488 26998 16540 27004
rect 16212 26852 16264 26858
rect 16212 26794 16264 26800
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 16224 26024 16252 26522
rect 16396 26376 16448 26382
rect 16394 26344 16396 26353
rect 16448 26344 16450 26353
rect 16500 26314 16528 26998
rect 16578 26888 16634 26897
rect 16578 26823 16634 26832
rect 16592 26790 16620 26823
rect 16580 26784 16632 26790
rect 16580 26726 16632 26732
rect 16580 26512 16632 26518
rect 16684 26500 16712 28358
rect 16776 27334 16804 28512
rect 16868 28490 16896 29446
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 16868 28393 16896 28426
rect 16854 28384 16910 28393
rect 16854 28319 16910 28328
rect 16960 27826 16988 29786
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 17040 29572 17092 29578
rect 17040 29514 17092 29520
rect 17052 29102 17080 29514
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17144 28762 17172 29582
rect 17236 29510 17264 30518
rect 17224 29504 17276 29510
rect 17222 29472 17224 29481
rect 17276 29472 17278 29481
rect 17222 29407 17278 29416
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17132 28756 17184 28762
rect 17132 28698 17184 28704
rect 17236 28150 17264 28970
rect 17224 28144 17276 28150
rect 17224 28086 17276 28092
rect 16960 27798 17080 27826
rect 16948 27668 17000 27674
rect 16948 27610 17000 27616
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16632 26472 16712 26500
rect 16580 26454 16632 26460
rect 16592 26382 16620 26454
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16394 26279 16450 26288
rect 16488 26308 16540 26314
rect 16488 26250 16540 26256
rect 16314 26140 16622 26149
rect 16314 26138 16320 26140
rect 16376 26138 16400 26140
rect 16456 26138 16480 26140
rect 16536 26138 16560 26140
rect 16616 26138 16622 26140
rect 16376 26086 16378 26138
rect 16558 26086 16560 26138
rect 16314 26084 16320 26086
rect 16376 26084 16400 26086
rect 16456 26084 16480 26086
rect 16536 26084 16560 26086
rect 16616 26084 16622 26086
rect 16314 26075 16622 26084
rect 16488 26036 16540 26042
rect 16224 25996 16344 26024
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16224 25362 16252 25842
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 16123 25248 16160 25276
rect 16123 24970 16151 25248
rect 16316 25140 16344 25996
rect 16488 25978 16540 25984
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 16408 25702 16436 25842
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 16500 25430 16528 25978
rect 16684 25898 16712 26318
rect 16592 25870 16712 25898
rect 16592 25430 16620 25870
rect 16776 25838 16804 26998
rect 16868 26586 16896 27270
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16960 26432 16988 27610
rect 17052 27538 17080 27798
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 17052 26994 17080 27474
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17144 27062 17172 27406
rect 17132 27056 17184 27062
rect 17132 26998 17184 27004
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 17040 26852 17092 26858
rect 17040 26794 17092 26800
rect 17052 26586 17080 26794
rect 17132 26784 17184 26790
rect 17132 26726 17184 26732
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 16868 26404 16988 26432
rect 16868 25906 16896 26404
rect 17040 26376 17092 26382
rect 16960 26336 17040 26364
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 16764 25832 16816 25838
rect 16764 25774 16816 25780
rect 16488 25424 16540 25430
rect 16488 25366 16540 25372
rect 16580 25424 16632 25430
rect 16580 25366 16632 25372
rect 16224 25112 16344 25140
rect 16123 24942 16160 24970
rect 16132 24886 16160 24942
rect 16120 24880 16172 24886
rect 16120 24822 16172 24828
rect 16224 24800 16252 25112
rect 16314 25052 16622 25061
rect 16314 25050 16320 25052
rect 16376 25050 16400 25052
rect 16456 25050 16480 25052
rect 16536 25050 16560 25052
rect 16616 25050 16622 25052
rect 16376 24998 16378 25050
rect 16558 24998 16560 25050
rect 16314 24996 16320 24998
rect 16376 24996 16400 24998
rect 16456 24996 16480 24998
rect 16536 24996 16560 24998
rect 16616 24996 16622 24998
rect 16314 24987 16622 24996
rect 16580 24880 16632 24886
rect 16580 24822 16632 24828
rect 16224 24772 16344 24800
rect 16040 24670 16252 24698
rect 15934 24647 15936 24656
rect 15988 24647 15990 24656
rect 15936 24618 15988 24624
rect 16028 24608 16080 24614
rect 16080 24568 16160 24596
rect 16028 24550 16080 24556
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 15750 23695 15806 23704
rect 15844 23724 15896 23730
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 15290 21927 15346 21936
rect 15384 21956 15436 21962
rect 15200 21898 15252 21904
rect 15384 21898 15436 21904
rect 15212 20874 15240 21898
rect 15290 21584 15346 21593
rect 15290 21519 15292 21528
rect 15344 21519 15346 21528
rect 15292 21490 15344 21496
rect 15396 21146 15424 21898
rect 15474 21856 15530 21865
rect 15474 21791 15530 21800
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15290 20904 15346 20913
rect 15200 20868 15252 20874
rect 15290 20839 15346 20848
rect 15200 20810 15252 20816
rect 15120 20686 15240 20714
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 15016 20256 15068 20262
rect 15212 20233 15240 20686
rect 15304 20398 15332 20839
rect 15488 20806 15516 21791
rect 15672 21672 15700 22034
rect 15580 21644 15700 21672
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15580 20618 15608 21644
rect 15764 20942 15792 23695
rect 15844 23666 15896 23672
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15856 23118 15884 23258
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15948 23050 15976 24346
rect 16132 24198 16160 24568
rect 16224 24342 16252 24670
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 16316 24206 16344 24772
rect 16394 24712 16450 24721
rect 16394 24647 16450 24656
rect 16488 24676 16540 24682
rect 16408 24274 16436 24647
rect 16488 24618 16540 24624
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16304 24200 16356 24206
rect 16132 24170 16252 24198
rect 16224 24052 16252 24170
rect 16304 24142 16356 24148
rect 16500 24052 16528 24618
rect 16592 24313 16620 24822
rect 16578 24304 16634 24313
rect 16578 24239 16634 24248
rect 16684 24154 16712 25774
rect 16762 25528 16818 25537
rect 16762 25463 16764 25472
rect 16816 25463 16818 25472
rect 16764 25434 16816 25440
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16776 24993 16804 25094
rect 16762 24984 16818 24993
rect 16762 24919 16818 24928
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16776 24274 16804 24754
rect 16868 24721 16896 25842
rect 16960 25838 16988 26336
rect 17144 26364 17172 26726
rect 17144 26336 17183 26364
rect 17040 26318 17092 26324
rect 17155 26246 17183 26336
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 17132 26240 17184 26246
rect 17236 26217 17264 28086
rect 17328 26994 17356 34303
rect 18236 32836 18288 32842
rect 18236 32778 18288 32784
rect 18248 32570 18276 32778
rect 18236 32564 18288 32570
rect 18236 32506 18288 32512
rect 18050 32464 18106 32473
rect 18892 32434 18920 34350
rect 19522 33144 19578 33153
rect 19522 33079 19578 33088
rect 19246 32872 19302 32881
rect 19246 32807 19302 32816
rect 18050 32399 18106 32408
rect 18880 32428 18932 32434
rect 17776 32224 17828 32230
rect 17776 32166 17828 32172
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 17420 30190 17448 31622
rect 17788 31521 17816 32166
rect 17774 31512 17830 31521
rect 17774 31447 17830 31456
rect 18064 31210 18092 32399
rect 18880 32370 18932 32376
rect 19064 32292 19116 32298
rect 19064 32234 19116 32240
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18800 32026 18828 32166
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18052 31204 18104 31210
rect 18052 31146 18104 31152
rect 18144 31204 18196 31210
rect 18144 31146 18196 31152
rect 17776 31136 17828 31142
rect 17776 31078 17828 31084
rect 17684 30932 17736 30938
rect 17684 30874 17736 30880
rect 17500 30796 17552 30802
rect 17500 30738 17552 30744
rect 17408 30184 17460 30190
rect 17408 30126 17460 30132
rect 17408 30048 17460 30054
rect 17408 29990 17460 29996
rect 17420 29306 17448 29990
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17408 28756 17460 28762
rect 17408 28698 17460 28704
rect 17420 27674 17448 28698
rect 17512 27674 17540 30738
rect 17696 30598 17724 30874
rect 17684 30592 17736 30598
rect 17684 30534 17736 30540
rect 17788 29850 17816 31078
rect 17868 30728 17920 30734
rect 17868 30670 17920 30676
rect 17776 29844 17828 29850
rect 17776 29786 17828 29792
rect 17684 29572 17736 29578
rect 17684 29514 17736 29520
rect 17592 29504 17644 29510
rect 17592 29446 17644 29452
rect 17604 28694 17632 29446
rect 17592 28688 17644 28694
rect 17592 28630 17644 28636
rect 17408 27668 17460 27674
rect 17408 27610 17460 27616
rect 17500 27668 17552 27674
rect 17500 27610 17552 27616
rect 17498 27568 17554 27577
rect 17604 27538 17632 28630
rect 17498 27503 17554 27512
rect 17592 27532 17644 27538
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17512 26926 17540 27503
rect 17592 27474 17644 27480
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17500 26920 17552 26926
rect 17406 26888 17462 26897
rect 17316 26852 17368 26858
rect 17500 26862 17552 26868
rect 17406 26823 17462 26832
rect 17316 26794 17368 26800
rect 17132 26182 17184 26188
rect 17222 26208 17278 26217
rect 16948 25832 17000 25838
rect 16948 25774 17000 25780
rect 16854 24712 16910 24721
rect 16854 24647 16910 24656
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16868 24313 16896 24550
rect 16854 24304 16910 24313
rect 16764 24268 16816 24274
rect 16854 24239 16910 24248
rect 16764 24210 16816 24216
rect 16856 24200 16908 24206
rect 16684 24126 16804 24154
rect 16856 24142 16908 24148
rect 16118 24032 16174 24041
rect 16224 24024 16528 24052
rect 16672 24064 16724 24070
rect 16776 24041 16804 24126
rect 16672 24006 16724 24012
rect 16762 24032 16818 24041
rect 16118 23967 16174 23976
rect 16132 23730 16160 23967
rect 16314 23964 16622 23973
rect 16314 23962 16320 23964
rect 16376 23962 16400 23964
rect 16456 23962 16480 23964
rect 16536 23962 16560 23964
rect 16616 23962 16622 23964
rect 16376 23910 16378 23962
rect 16558 23910 16560 23962
rect 16314 23908 16320 23910
rect 16376 23908 16400 23910
rect 16456 23908 16480 23910
rect 16536 23908 16560 23910
rect 16616 23908 16622 23910
rect 16314 23899 16622 23908
rect 16684 23798 16712 24006
rect 16762 23967 16818 23976
rect 16868 23882 16896 24142
rect 16960 24138 16988 25774
rect 16948 24132 17000 24138
rect 16948 24074 17000 24080
rect 16776 23854 16896 23882
rect 16672 23792 16724 23798
rect 16672 23734 16724 23740
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16212 23724 16264 23730
rect 16212 23666 16264 23672
rect 16120 23588 16172 23594
rect 16224 23576 16252 23666
rect 16776 23662 16804 23854
rect 16856 23792 16908 23798
rect 16856 23734 16908 23740
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16172 23548 16252 23576
rect 16580 23588 16632 23594
rect 16120 23530 16172 23536
rect 16580 23530 16632 23536
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16408 23361 16436 23462
rect 16210 23352 16266 23361
rect 16394 23352 16450 23361
rect 16266 23310 16344 23338
rect 16210 23287 16266 23296
rect 16120 23180 16172 23186
rect 16040 23140 16120 23168
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15842 22808 15898 22817
rect 15842 22743 15898 22752
rect 15856 22710 15884 22743
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 15842 22400 15898 22409
rect 15842 22335 15898 22344
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15856 20874 15884 22335
rect 15948 22030 15976 22986
rect 16040 22953 16068 23140
rect 16120 23122 16172 23128
rect 16212 23112 16264 23118
rect 16316 23100 16344 23310
rect 16592 23322 16620 23530
rect 16394 23287 16450 23296
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16396 23112 16448 23118
rect 16316 23072 16396 23100
rect 16212 23054 16264 23060
rect 16396 23054 16448 23060
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 16026 22944 16082 22953
rect 16026 22879 16082 22888
rect 16132 22778 16160 22986
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 16040 22574 16068 22714
rect 16028 22568 16080 22574
rect 16028 22510 16080 22516
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 16040 21962 16068 22510
rect 16224 22506 16252 23054
rect 16684 22982 16712 23258
rect 16868 23118 16896 23734
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16314 22876 16622 22885
rect 16314 22874 16320 22876
rect 16376 22874 16400 22876
rect 16456 22874 16480 22876
rect 16536 22874 16560 22876
rect 16616 22874 16622 22876
rect 16376 22822 16378 22874
rect 16558 22822 16560 22874
rect 16314 22820 16320 22822
rect 16376 22820 16400 22822
rect 16456 22820 16480 22822
rect 16536 22820 16560 22822
rect 16616 22820 16622 22822
rect 16314 22811 16622 22820
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16212 22500 16264 22506
rect 16212 22442 16264 22448
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16132 21865 16160 22034
rect 16316 21876 16344 22578
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16500 21962 16528 22442
rect 16592 22166 16620 22714
rect 16776 22642 16804 22918
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16670 22264 16726 22273
rect 16670 22199 16726 22208
rect 16580 22160 16632 22166
rect 16580 22102 16632 22108
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16118 21856 16174 21865
rect 16118 21791 16174 21800
rect 16224 21848 16344 21876
rect 16118 21720 16174 21729
rect 16028 21684 16080 21690
rect 16118 21655 16120 21664
rect 16028 21626 16080 21632
rect 16172 21655 16174 21664
rect 16120 21626 16172 21632
rect 16040 21554 16068 21626
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 15948 21418 15976 21490
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 16224 21298 16252 21848
rect 16314 21788 16622 21797
rect 16314 21786 16320 21788
rect 16376 21786 16400 21788
rect 16456 21786 16480 21788
rect 16536 21786 16560 21788
rect 16616 21786 16622 21788
rect 16376 21734 16378 21786
rect 16558 21734 16560 21786
rect 16314 21732 16320 21734
rect 16376 21732 16400 21734
rect 16456 21732 16480 21734
rect 16536 21732 16560 21734
rect 16616 21732 16622 21734
rect 16314 21723 16622 21732
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 16132 21270 16252 21298
rect 16026 21176 16082 21185
rect 16026 21111 16082 21120
rect 16040 20874 16068 21111
rect 16132 21078 16160 21270
rect 16316 21078 16344 21558
rect 16394 21176 16450 21185
rect 16394 21111 16450 21120
rect 16488 21140 16540 21146
rect 16120 21072 16172 21078
rect 16120 21014 16172 21020
rect 16304 21072 16356 21078
rect 16304 21014 16356 21020
rect 16408 21010 16436 21111
rect 16488 21082 16540 21088
rect 16500 21010 16528 21082
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16592 20942 16620 21626
rect 16684 21622 16712 22199
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 16776 21400 16804 22442
rect 16868 21842 16896 22646
rect 16960 22506 16988 23054
rect 17052 22506 17080 26182
rect 17222 26143 17278 26152
rect 17328 26081 17356 26794
rect 17420 26450 17448 26823
rect 17604 26586 17632 27338
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 17498 26480 17554 26489
rect 17408 26444 17460 26450
rect 17498 26415 17554 26424
rect 17592 26444 17644 26450
rect 17408 26386 17460 26392
rect 17408 26308 17460 26314
rect 17408 26250 17460 26256
rect 17314 26072 17370 26081
rect 17314 26007 17370 26016
rect 17420 25956 17448 26250
rect 17328 25928 17448 25956
rect 17224 25764 17276 25770
rect 17224 25706 17276 25712
rect 17236 25650 17264 25706
rect 17226 25622 17264 25650
rect 17130 25528 17186 25537
rect 17226 25498 17254 25622
rect 17130 25463 17132 25472
rect 17184 25463 17186 25472
rect 17224 25492 17276 25498
rect 17132 25434 17184 25440
rect 17224 25434 17276 25440
rect 17328 25430 17356 25928
rect 17512 25888 17540 26415
rect 17696 26432 17724 29514
rect 17774 29472 17830 29481
rect 17774 29407 17830 29416
rect 17788 29170 17816 29407
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17776 28688 17828 28694
rect 17776 28630 17828 28636
rect 17644 26404 17724 26432
rect 17592 26386 17644 26392
rect 17604 26353 17632 26386
rect 17590 26344 17646 26353
rect 17590 26279 17646 26288
rect 17592 25900 17644 25906
rect 17512 25860 17592 25888
rect 17592 25842 17644 25848
rect 17408 25696 17460 25702
rect 17684 25696 17736 25702
rect 17408 25638 17460 25644
rect 17682 25664 17684 25673
rect 17736 25664 17738 25673
rect 17316 25424 17368 25430
rect 17316 25366 17368 25372
rect 17316 25288 17368 25294
rect 17420 25276 17448 25638
rect 17682 25599 17738 25608
rect 17498 25528 17554 25537
rect 17498 25463 17500 25472
rect 17552 25463 17554 25472
rect 17500 25434 17552 25440
rect 17696 25412 17724 25599
rect 17788 25498 17816 28630
rect 17880 27674 17908 30670
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17972 28506 18000 29990
rect 18064 29170 18092 30602
rect 18156 30297 18184 31146
rect 18142 30288 18198 30297
rect 18142 30223 18198 30232
rect 18144 30116 18196 30122
rect 18144 30058 18196 30064
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18064 28762 18092 29106
rect 18052 28756 18104 28762
rect 18052 28698 18104 28704
rect 17972 28478 18092 28506
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 17972 27606 18000 28358
rect 17960 27600 18012 27606
rect 17866 27568 17922 27577
rect 18064 27577 18092 28478
rect 17960 27542 18012 27548
rect 18050 27568 18106 27577
rect 17866 27503 17922 27512
rect 17880 26625 17908 27503
rect 17972 27452 18000 27542
rect 18050 27503 18106 27512
rect 17972 27424 18092 27452
rect 18064 26994 18092 27424
rect 18156 27044 18184 30058
rect 18248 29850 18276 31962
rect 18328 31748 18380 31754
rect 18328 31690 18380 31696
rect 18340 30938 18368 31690
rect 18420 31340 18472 31346
rect 18420 31282 18472 31288
rect 18328 30932 18380 30938
rect 18328 30874 18380 30880
rect 18340 30258 18368 30874
rect 18328 30252 18380 30258
rect 18328 30194 18380 30200
rect 18236 29844 18288 29850
rect 18236 29786 18288 29792
rect 18340 29510 18368 30194
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18236 29164 18288 29170
rect 18236 29106 18288 29112
rect 18248 28937 18276 29106
rect 18234 28928 18290 28937
rect 18234 28863 18290 28872
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18248 27470 18276 28494
rect 18432 27849 18460 31282
rect 18972 31136 19024 31142
rect 18972 31078 19024 31084
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18616 30054 18644 30194
rect 18604 30048 18656 30054
rect 18604 29990 18656 29996
rect 18708 29617 18736 30874
rect 18984 30705 19012 31078
rect 18970 30696 19026 30705
rect 18970 30631 19026 30640
rect 18972 30592 19024 30598
rect 18972 30534 19024 30540
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18788 29776 18840 29782
rect 18786 29744 18788 29753
rect 18840 29744 18842 29753
rect 18786 29679 18842 29688
rect 18510 29608 18566 29617
rect 18510 29543 18566 29552
rect 18694 29608 18750 29617
rect 18694 29543 18750 29552
rect 18524 28937 18552 29543
rect 18602 29336 18658 29345
rect 18602 29271 18658 29280
rect 18696 29300 18748 29306
rect 18510 28928 18566 28937
rect 18510 28863 18566 28872
rect 18512 28756 18564 28762
rect 18512 28698 18564 28704
rect 18524 28064 18552 28698
rect 18616 28370 18644 29271
rect 18696 29242 18748 29248
rect 18708 28558 18736 29242
rect 18788 29028 18840 29034
rect 18788 28970 18840 28976
rect 18800 28665 18828 28970
rect 18786 28656 18842 28665
rect 18786 28591 18842 28600
rect 18696 28552 18748 28558
rect 18696 28494 18748 28500
rect 18616 28342 18736 28370
rect 18602 28248 18658 28257
rect 18708 28218 18736 28342
rect 18602 28183 18604 28192
rect 18656 28183 18658 28192
rect 18696 28212 18748 28218
rect 18604 28154 18656 28160
rect 18696 28154 18748 28160
rect 18788 28076 18840 28082
rect 18524 28036 18736 28064
rect 18418 27840 18474 27849
rect 18602 27840 18658 27849
rect 18418 27775 18474 27784
rect 18524 27798 18602 27826
rect 18432 27606 18460 27775
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 18420 27600 18472 27606
rect 18420 27542 18472 27548
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 18340 27169 18368 27542
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18326 27160 18382 27169
rect 18326 27095 18382 27104
rect 18236 27056 18288 27062
rect 18156 27016 18236 27044
rect 18236 26998 18288 27004
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17866 26616 17922 26625
rect 17866 26551 17868 26560
rect 17920 26551 17922 26560
rect 17868 26522 17920 26528
rect 17972 26489 18000 26726
rect 17958 26480 18014 26489
rect 17868 26444 17920 26450
rect 17958 26415 18014 26424
rect 17868 26386 17920 26392
rect 17880 25888 17908 26386
rect 17880 25860 18000 25888
rect 17868 25696 17920 25702
rect 17868 25638 17920 25644
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17604 25384 17724 25412
rect 17500 25288 17552 25294
rect 17420 25248 17500 25276
rect 17316 25230 17368 25236
rect 17604 25265 17632 25384
rect 17880 25344 17908 25638
rect 17696 25316 17908 25344
rect 17500 25230 17552 25236
rect 17590 25256 17646 25265
rect 17328 24857 17356 25230
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17130 24848 17186 24857
rect 17314 24848 17370 24857
rect 17130 24783 17186 24792
rect 17224 24812 17276 24818
rect 17144 23730 17172 24783
rect 17314 24783 17370 24792
rect 17224 24754 17276 24760
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17130 23352 17186 23361
rect 17130 23287 17186 23296
rect 17144 23186 17172 23287
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 16948 22500 17000 22506
rect 16948 22442 17000 22448
rect 17040 22500 17092 22506
rect 17040 22442 17092 22448
rect 16946 22264 17002 22273
rect 17144 22234 17172 22986
rect 17236 22681 17264 24754
rect 17328 24206 17356 24783
rect 17420 24682 17448 25094
rect 17512 24721 17540 25230
rect 17590 25191 17646 25200
rect 17498 24712 17554 24721
rect 17408 24676 17460 24682
rect 17498 24647 17554 24656
rect 17408 24618 17460 24624
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17406 24440 17462 24449
rect 17406 24375 17462 24384
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17420 24070 17448 24375
rect 17498 24304 17554 24313
rect 17498 24239 17554 24248
rect 17512 24206 17540 24239
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17604 23905 17632 24550
rect 17314 23896 17370 23905
rect 17314 23831 17370 23840
rect 17590 23896 17646 23905
rect 17590 23831 17646 23840
rect 17328 23730 17356 23831
rect 17696 23730 17724 25316
rect 17868 25220 17920 25226
rect 17788 25180 17868 25208
rect 17788 25129 17816 25180
rect 17868 25162 17920 25168
rect 17972 25129 18000 25860
rect 18064 25158 18092 26930
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18248 26518 18276 26862
rect 18328 26852 18380 26858
rect 18328 26794 18380 26800
rect 18340 26761 18368 26794
rect 18326 26752 18382 26761
rect 18326 26687 18382 26696
rect 18236 26512 18288 26518
rect 18142 26480 18198 26489
rect 18236 26454 18288 26460
rect 18142 26415 18198 26424
rect 18156 26246 18184 26415
rect 18432 26382 18460 27406
rect 18236 26376 18288 26382
rect 18420 26376 18472 26382
rect 18326 26344 18382 26353
rect 18288 26324 18326 26330
rect 18236 26318 18326 26324
rect 18248 26302 18326 26318
rect 18420 26318 18472 26324
rect 18326 26279 18382 26288
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18326 26208 18382 26217
rect 18052 25152 18104 25158
rect 17774 25120 17830 25129
rect 17774 25055 17830 25064
rect 17958 25120 18014 25129
rect 18052 25094 18104 25100
rect 17958 25055 18014 25064
rect 18156 24936 18184 26182
rect 18326 26143 18382 26152
rect 18234 26072 18290 26081
rect 18234 26007 18290 26016
rect 18248 25974 18276 26007
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 18236 25832 18288 25838
rect 18340 25786 18368 26143
rect 18432 26081 18460 26318
rect 18418 26072 18474 26081
rect 18418 26007 18474 26016
rect 18418 25936 18474 25945
rect 18418 25871 18420 25880
rect 18472 25871 18474 25880
rect 18420 25842 18472 25848
rect 18236 25774 18288 25780
rect 18248 25702 18276 25774
rect 18328 25758 18368 25786
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18328 25514 18356 25758
rect 18524 25650 18552 27798
rect 18708 27826 18736 28036
rect 18788 28018 18840 28024
rect 18602 27775 18658 27784
rect 18694 27798 18736 27826
rect 18694 27690 18722 27798
rect 18616 27662 18722 27690
rect 18616 26926 18644 27662
rect 18696 27464 18748 27470
rect 18800 27452 18828 28018
rect 18892 27713 18920 29990
rect 18984 28257 19012 30534
rect 19076 29578 19104 32234
rect 19156 31476 19208 31482
rect 19156 31418 19208 31424
rect 19064 29572 19116 29578
rect 19064 29514 19116 29520
rect 18970 28248 19026 28257
rect 18970 28183 19026 28192
rect 18984 28082 19012 28183
rect 18978 28076 19030 28082
rect 18978 28018 19030 28024
rect 18970 27976 19026 27985
rect 19076 27962 19104 29514
rect 19168 28218 19196 31418
rect 19260 30841 19288 32807
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 19246 30832 19302 30841
rect 19246 30767 19302 30776
rect 19352 30433 19380 30874
rect 19536 30598 19564 33079
rect 19892 32836 19944 32842
rect 19892 32778 19944 32784
rect 19904 32026 19932 32778
rect 20088 32434 20116 34350
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 21640 32768 21692 32774
rect 21640 32710 21692 32716
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 20155 32124 20463 32133
rect 20155 32122 20161 32124
rect 20217 32122 20241 32124
rect 20297 32122 20321 32124
rect 20377 32122 20401 32124
rect 20457 32122 20463 32124
rect 20217 32070 20219 32122
rect 20399 32070 20401 32122
rect 20155 32068 20161 32070
rect 20217 32068 20241 32070
rect 20297 32068 20321 32070
rect 20377 32068 20401 32070
rect 20457 32068 20463 32070
rect 20155 32059 20463 32068
rect 20534 32056 20590 32065
rect 19892 32020 19944 32026
rect 19720 31980 19892 32008
rect 19614 31648 19670 31657
rect 19614 31583 19670 31592
rect 19524 30592 19576 30598
rect 19524 30534 19576 30540
rect 19338 30424 19394 30433
rect 19248 30388 19300 30394
rect 19338 30359 19394 30368
rect 19432 30388 19484 30394
rect 19248 30330 19300 30336
rect 19432 30330 19484 30336
rect 19260 30122 19288 30330
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19248 30116 19300 30122
rect 19248 30058 19300 30064
rect 19248 29708 19300 29714
rect 19248 29650 19300 29656
rect 19260 29492 19288 29650
rect 19352 29617 19380 30262
rect 19444 30025 19472 30330
rect 19536 30297 19564 30534
rect 19522 30288 19578 30297
rect 19522 30223 19578 30232
rect 19430 30016 19486 30025
rect 19430 29951 19486 29960
rect 19432 29844 19484 29850
rect 19432 29786 19484 29792
rect 19338 29608 19394 29617
rect 19338 29543 19394 29552
rect 19260 29464 19380 29492
rect 19246 29200 19302 29209
rect 19246 29135 19248 29144
rect 19300 29135 19302 29144
rect 19248 29106 19300 29112
rect 19246 28928 19302 28937
rect 19246 28863 19302 28872
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19168 27985 19196 28018
rect 19026 27934 19104 27962
rect 19154 27976 19210 27985
rect 18970 27911 19026 27920
rect 19154 27911 19210 27920
rect 18878 27704 18934 27713
rect 18878 27639 18934 27648
rect 18748 27424 18828 27452
rect 18696 27406 18748 27412
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18708 26382 18736 27406
rect 18785 26784 18837 26790
rect 18785 26726 18837 26732
rect 18696 26376 18748 26382
rect 18602 26344 18658 26353
rect 18696 26318 18748 26324
rect 18602 26279 18658 26288
rect 18616 26246 18644 26279
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18602 26072 18658 26081
rect 18708 26042 18736 26318
rect 18602 26007 18658 26016
rect 18696 26036 18748 26042
rect 18616 25770 18644 26007
rect 18696 25978 18748 25984
rect 18604 25764 18656 25770
rect 18604 25706 18656 25712
rect 18524 25622 18736 25650
rect 18328 25486 18368 25514
rect 18340 25294 18368 25486
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 18236 25220 18288 25226
rect 18236 25162 18288 25168
rect 18064 24908 18184 24936
rect 17776 24880 17828 24886
rect 17828 24840 17908 24868
rect 17776 24822 17828 24828
rect 17880 24188 17908 24840
rect 18064 24818 18092 24908
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17958 24712 18014 24721
rect 17958 24647 18014 24656
rect 18052 24676 18104 24682
rect 17972 24614 18000 24647
rect 18052 24618 18104 24624
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 18064 24256 18092 24618
rect 18156 24313 18184 24754
rect 18063 24228 18092 24256
rect 18142 24304 18198 24313
rect 18142 24239 18198 24248
rect 17960 24200 18012 24206
rect 17880 24160 17960 24188
rect 17960 24142 18012 24148
rect 18063 24154 18091 24228
rect 18144 24200 18196 24206
rect 18063 24126 18092 24154
rect 18144 24142 18196 24148
rect 17868 24064 17920 24070
rect 17788 24024 17868 24052
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17788 23304 17816 24024
rect 17868 24006 17920 24012
rect 17958 24032 18014 24041
rect 17958 23967 18014 23976
rect 17972 23712 18000 23967
rect 17420 23276 17816 23304
rect 17880 23684 18000 23712
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17328 22817 17356 23054
rect 17420 22953 17448 23276
rect 17774 23216 17830 23225
rect 17880 23202 17908 23684
rect 18064 23610 18092 24126
rect 18156 24041 18184 24142
rect 18142 24032 18198 24041
rect 18142 23967 18198 23976
rect 18142 23896 18198 23905
rect 18142 23831 18198 23840
rect 18156 23798 18184 23831
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 17830 23186 17908 23202
rect 17972 23582 18092 23610
rect 18144 23588 18196 23594
rect 17830 23180 17920 23186
rect 17830 23174 17868 23180
rect 17774 23151 17830 23160
rect 17868 23122 17920 23128
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17406 22944 17462 22953
rect 17406 22879 17462 22888
rect 17314 22808 17370 22817
rect 17314 22743 17370 22752
rect 17408 22704 17460 22710
rect 17222 22672 17278 22681
rect 17408 22646 17460 22652
rect 17222 22607 17278 22616
rect 16946 22199 17002 22208
rect 17132 22228 17184 22234
rect 16960 22098 16988 22199
rect 17132 22170 17184 22176
rect 17236 22137 17264 22607
rect 17316 22500 17368 22506
rect 17316 22442 17368 22448
rect 17222 22128 17278 22137
rect 16948 22092 17000 22098
rect 17328 22098 17356 22442
rect 17420 22438 17448 22646
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 17222 22063 17278 22072
rect 17316 22092 17368 22098
rect 16948 22034 17000 22040
rect 17316 22034 17368 22040
rect 17420 22030 17448 22102
rect 17408 22024 17460 22030
rect 17130 21992 17186 22001
rect 17408 21966 17460 21972
rect 17130 21927 17186 21936
rect 16868 21814 16988 21842
rect 16844 21684 16896 21690
rect 16960 21672 16988 21814
rect 17040 21684 17092 21690
rect 16960 21644 17040 21672
rect 16844 21626 16896 21632
rect 17040 21626 17092 21632
rect 16868 21604 16896 21626
rect 16868 21576 16988 21604
rect 16960 21570 16988 21576
rect 17144 21570 17172 21927
rect 17316 21888 17368 21894
rect 17368 21836 17448 21842
rect 17316 21830 17448 21836
rect 17328 21814 17448 21830
rect 17420 21690 17448 21814
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17328 21593 17356 21626
rect 16960 21542 17172 21570
rect 17314 21584 17370 21593
rect 17314 21519 17370 21528
rect 16776 21372 16896 21400
rect 16868 21078 16896 21372
rect 16856 21072 16908 21078
rect 16670 21040 16726 21049
rect 16856 21014 16908 21020
rect 16670 20975 16726 20984
rect 16580 20936 16632 20942
rect 16302 20904 16358 20913
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 16028 20868 16080 20874
rect 16358 20862 16528 20890
rect 16580 20878 16632 20884
rect 16302 20839 16358 20848
rect 16028 20810 16080 20816
rect 15660 20800 15712 20806
rect 15658 20768 15660 20777
rect 15936 20800 15988 20806
rect 15712 20768 15714 20777
rect 15658 20703 15714 20712
rect 15856 20748 15936 20754
rect 16500 20788 16528 20862
rect 16684 20788 16712 20975
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16500 20760 16712 20788
rect 15856 20742 15988 20748
rect 15856 20726 15976 20742
rect 15580 20590 15792 20618
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15016 20198 15068 20204
rect 15198 20224 15254 20233
rect 15198 20159 15254 20168
rect 14830 20088 14886 20097
rect 14830 20023 14886 20032
rect 14844 19854 14872 20023
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14752 19700 14780 19790
rect 15028 19700 15056 19790
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 14752 19672 15056 19700
rect 14740 19372 14792 19378
rect 14792 19320 14872 19334
rect 14740 19314 14872 19320
rect 14752 19306 14872 19314
rect 14462 19000 14518 19009
rect 13728 18906 13780 18912
rect 13832 18924 13952 18952
rect 14280 18964 14332 18970
rect 13740 18766 13768 18906
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13648 17610 13676 18226
rect 13740 18086 13768 18566
rect 13832 18329 13860 18924
rect 14462 18935 14518 18944
rect 14280 18906 14332 18912
rect 13910 18864 13966 18873
rect 13910 18799 13966 18808
rect 14004 18828 14056 18834
rect 13818 18320 13874 18329
rect 13818 18255 13874 18264
rect 13924 18154 13952 18799
rect 14004 18770 14056 18776
rect 14016 18222 14044 18770
rect 14462 18728 14518 18737
rect 14462 18663 14518 18672
rect 14476 18358 14504 18663
rect 14096 18352 14148 18358
rect 14094 18320 14096 18329
rect 14280 18352 14332 18358
rect 14148 18320 14150 18329
rect 14464 18352 14516 18358
rect 14332 18312 14412 18340
rect 14280 18294 14332 18300
rect 14094 18255 14150 18264
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13648 12434 13676 17274
rect 13740 16998 13768 17478
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13740 14482 13768 16662
rect 13832 16114 13860 18022
rect 13924 16114 13952 18090
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13924 15994 13952 16050
rect 13832 15966 13952 15994
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13832 14074 13860 15966
rect 13912 15088 13964 15094
rect 13910 15056 13912 15065
rect 13964 15056 13966 15065
rect 13910 14991 13966 15000
rect 14016 14940 14044 18158
rect 14096 17332 14148 17338
rect 14200 17320 14228 18158
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 14148 17292 14228 17320
rect 14096 17274 14148 17280
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16833 14136 16934
rect 14094 16824 14150 16833
rect 14094 16759 14150 16768
rect 14200 16697 14228 17292
rect 14292 16998 14320 17546
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14186 16688 14242 16697
rect 14186 16623 14242 16632
rect 14200 16590 14228 16623
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14200 16250 14228 16526
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14186 16008 14242 16017
rect 14096 15972 14148 15978
rect 14186 15943 14188 15952
rect 14096 15914 14148 15920
rect 14240 15943 14242 15952
rect 14188 15914 14240 15920
rect 13924 14912 14044 14940
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13924 12434 13952 14912
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 13802 14044 14758
rect 14108 14074 14136 15914
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 14292 13190 14320 16934
rect 14384 16697 14412 18312
rect 14844 18340 14872 19306
rect 14924 19168 14976 19174
rect 14922 19136 14924 19145
rect 14976 19136 14978 19145
rect 14922 19071 14978 19080
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14936 18465 14964 18634
rect 14922 18456 14978 18465
rect 15028 18426 15056 18906
rect 15120 18698 15148 19722
rect 15212 19394 15240 20159
rect 15382 20088 15438 20097
rect 15382 20023 15438 20032
rect 15396 19530 15424 20023
rect 15488 19854 15516 20334
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15580 19666 15608 19790
rect 15672 19786 15700 20402
rect 15660 19780 15712 19786
rect 15660 19722 15712 19728
rect 15580 19638 15700 19666
rect 15396 19502 15608 19530
rect 15212 19366 15332 19394
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15212 19122 15240 19246
rect 15304 19242 15332 19366
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15384 19236 15436 19242
rect 15384 19178 15436 19184
rect 15212 19094 15332 19122
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 14922 18391 14978 18400
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 14924 18352 14976 18358
rect 14844 18312 14924 18340
rect 14464 18294 14516 18300
rect 14924 18294 14976 18300
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14464 18148 14516 18154
rect 14568 18136 14596 18226
rect 14516 18108 14596 18136
rect 14464 18090 14516 18096
rect 14832 18080 14884 18086
rect 14830 18048 14832 18057
rect 14884 18048 14886 18057
rect 14830 17983 14886 17992
rect 14554 17912 14610 17921
rect 14554 17847 14556 17856
rect 14608 17847 14610 17856
rect 14556 17818 14608 17824
rect 14936 17785 14964 18294
rect 15304 18086 15332 19094
rect 15396 18873 15424 19178
rect 15488 18970 15516 19246
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15382 18864 15438 18873
rect 15382 18799 15438 18808
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15154 18080 15206 18086
rect 15154 18022 15206 18028
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 14922 17776 14978 17785
rect 14922 17711 14978 17720
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14568 17320 14596 17546
rect 14936 17490 14964 17711
rect 15028 17678 15056 18022
rect 15166 17898 15194 18022
rect 15166 17870 15224 17898
rect 15196 17814 15224 17870
rect 15108 17808 15160 17814
rect 15106 17776 15108 17785
rect 15196 17808 15252 17814
rect 15160 17776 15162 17785
rect 15196 17768 15200 17808
rect 15200 17750 15252 17756
rect 15106 17711 15162 17720
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15200 17536 15252 17542
rect 14936 17462 15056 17490
rect 15200 17478 15252 17484
rect 14568 17292 14780 17320
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14554 17096 14610 17105
rect 14554 17031 14610 17040
rect 14462 16824 14518 16833
rect 14462 16759 14518 16768
rect 14370 16688 14426 16697
rect 14370 16623 14426 16632
rect 14384 16454 14412 16623
rect 14476 16590 14504 16759
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14372 16448 14424 16454
rect 14464 16448 14516 16454
rect 14372 16390 14424 16396
rect 14462 16416 14464 16425
rect 14516 16416 14518 16425
rect 14462 16351 14518 16360
rect 14568 16232 14596 17031
rect 14660 16522 14688 17138
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14752 16425 14780 17292
rect 15028 17202 15056 17462
rect 15212 17338 15240 17478
rect 15200 17332 15252 17338
rect 15396 17320 15424 18799
rect 15580 18698 15608 19502
rect 15672 18834 15700 19638
rect 15764 18873 15792 20590
rect 15856 19689 15884 20726
rect 16314 20700 16622 20709
rect 16314 20698 16320 20700
rect 16376 20698 16400 20700
rect 16456 20698 16480 20700
rect 16536 20698 16560 20700
rect 16616 20698 16622 20700
rect 16376 20646 16378 20698
rect 16558 20646 16560 20698
rect 16314 20644 16320 20646
rect 16376 20644 16400 20646
rect 16456 20644 16480 20646
rect 16536 20644 16560 20646
rect 16616 20644 16622 20646
rect 16118 20632 16174 20641
rect 16314 20635 16622 20644
rect 16776 20641 16804 20810
rect 16118 20567 16174 20576
rect 16762 20632 16818 20641
rect 16762 20567 16818 20576
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15948 19718 15976 20334
rect 16132 20262 16160 20567
rect 16868 20482 16896 21014
rect 17512 20992 17540 23054
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17604 21486 17632 22578
rect 17696 22273 17724 23054
rect 17868 23044 17920 23050
rect 17868 22986 17920 22992
rect 17774 22944 17830 22953
rect 17774 22879 17830 22888
rect 17788 22574 17816 22879
rect 17880 22817 17908 22986
rect 17866 22808 17922 22817
rect 17866 22743 17922 22752
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 17682 22264 17738 22273
rect 17682 22199 17738 22208
rect 17696 22001 17724 22199
rect 17776 22024 17828 22030
rect 17682 21992 17738 22001
rect 17776 21966 17828 21972
rect 17682 21927 17738 21936
rect 17788 21593 17816 21966
rect 17774 21584 17830 21593
rect 17684 21548 17736 21554
rect 17774 21519 17830 21528
rect 17684 21490 17736 21496
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17696 21418 17724 21490
rect 17880 21457 17908 22646
rect 17972 22506 18000 23582
rect 18144 23530 18196 23536
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 18064 22166 18092 23462
rect 18156 22710 18184 23530
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 18052 22160 18104 22166
rect 18052 22102 18104 22108
rect 18156 22030 18184 22646
rect 18248 22642 18276 25162
rect 18340 24206 18368 25230
rect 18432 24410 18460 25434
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18418 24304 18474 24313
rect 18418 24239 18474 24248
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18340 23905 18368 24142
rect 18326 23896 18382 23905
rect 18326 23831 18382 23840
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18340 23594 18368 23734
rect 18432 23730 18460 24239
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18328 23588 18380 23594
rect 18328 23530 18380 23536
rect 18326 23352 18382 23361
rect 18326 23287 18382 23296
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18052 22024 18104 22030
rect 17958 21992 18014 22001
rect 18052 21966 18104 21972
rect 18144 22024 18196 22030
rect 18248 22012 18276 22578
rect 18340 22166 18368 23287
rect 18420 23248 18472 23254
rect 18420 23190 18472 23196
rect 18432 22953 18460 23190
rect 18418 22944 18474 22953
rect 18418 22879 18474 22888
rect 18418 22808 18474 22817
rect 18418 22743 18474 22752
rect 18432 22250 18460 22743
rect 18524 22506 18552 25230
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18616 24818 18644 25094
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18602 24576 18658 24585
rect 18602 24511 18658 24520
rect 18616 24206 18644 24511
rect 18708 24342 18736 25622
rect 18800 25294 18828 26726
rect 18892 25906 18920 27639
rect 18984 26926 19012 27911
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 19076 27577 19104 27814
rect 19062 27568 19118 27577
rect 19062 27503 19118 27512
rect 19168 26994 19196 27911
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18892 25673 18920 25842
rect 18878 25664 18934 25673
rect 18878 25599 18934 25608
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 18800 25158 18828 25230
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18786 24984 18842 24993
rect 18786 24919 18842 24928
rect 18800 24886 18828 24919
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 18984 24818 19012 26862
rect 19076 26246 19104 26930
rect 19156 26376 19208 26382
rect 19156 26318 19208 26324
rect 19064 26240 19116 26246
rect 19064 26182 19116 26188
rect 19062 26072 19118 26081
rect 19062 26007 19118 26016
rect 19076 25838 19104 26007
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 19168 25752 19196 26318
rect 19260 25916 19288 28863
rect 19352 28665 19380 29464
rect 19444 28937 19472 29786
rect 19628 29714 19656 31583
rect 19616 29708 19668 29714
rect 19616 29650 19668 29656
rect 19524 29640 19576 29646
rect 19524 29582 19576 29588
rect 19430 28928 19486 28937
rect 19430 28863 19486 28872
rect 19338 28656 19394 28665
rect 19338 28591 19394 28600
rect 19352 28490 19380 28591
rect 19340 28484 19392 28490
rect 19340 28426 19392 28432
rect 19430 28384 19486 28393
rect 19430 28319 19486 28328
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 19352 28082 19380 28154
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 19352 27470 19380 27542
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19444 26790 19472 28319
rect 19432 26784 19484 26790
rect 19352 26744 19432 26772
rect 19255 25910 19307 25916
rect 19255 25852 19307 25858
rect 19248 25764 19300 25770
rect 19168 25724 19248 25752
rect 19248 25706 19300 25712
rect 19352 25650 19380 26744
rect 19432 26726 19484 26732
rect 19430 26616 19486 26625
rect 19430 26551 19486 26560
rect 19444 25702 19472 26551
rect 19536 25786 19564 29582
rect 19720 28626 19748 31980
rect 19892 31962 19944 31968
rect 19984 32020 20036 32026
rect 20534 31991 20590 32000
rect 19984 31962 20036 31968
rect 19892 31680 19944 31686
rect 19892 31622 19944 31628
rect 19800 31136 19852 31142
rect 19800 31078 19852 31084
rect 19812 30326 19840 31078
rect 19904 30376 19932 31622
rect 19996 31113 20024 31962
rect 20076 31952 20128 31958
rect 20076 31894 20128 31900
rect 19982 31104 20038 31113
rect 19982 31039 20038 31048
rect 20088 30705 20116 31894
rect 20548 31346 20576 31991
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20155 31036 20463 31045
rect 20155 31034 20161 31036
rect 20217 31034 20241 31036
rect 20297 31034 20321 31036
rect 20377 31034 20401 31036
rect 20457 31034 20463 31036
rect 20217 30982 20219 31034
rect 20399 30982 20401 31034
rect 20155 30980 20161 30982
rect 20217 30980 20241 30982
rect 20297 30980 20321 30982
rect 20377 30980 20401 30982
rect 20457 30980 20463 30982
rect 20155 30971 20463 30980
rect 20534 30968 20590 30977
rect 20180 30912 20534 30920
rect 20180 30903 20590 30912
rect 20180 30892 20576 30903
rect 20074 30696 20130 30705
rect 20074 30631 20130 30640
rect 19904 30348 20024 30376
rect 19800 30320 19852 30326
rect 19800 30262 19852 30268
rect 19890 30288 19946 30297
rect 19708 28620 19760 28626
rect 19708 28562 19760 28568
rect 19616 28416 19668 28422
rect 19616 28358 19668 28364
rect 19628 28218 19656 28358
rect 19616 28212 19668 28218
rect 19616 28154 19668 28160
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19628 27849 19656 27950
rect 19614 27840 19670 27849
rect 19614 27775 19670 27784
rect 19720 27588 19748 28562
rect 19812 27946 19840 30262
rect 19890 30223 19946 30232
rect 19904 29889 19932 30223
rect 19890 29880 19946 29889
rect 19996 29850 20024 30348
rect 20076 30184 20128 30190
rect 20076 30126 20128 30132
rect 19890 29815 19946 29824
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19904 29481 19932 29650
rect 19996 29646 20024 29786
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19890 29472 19946 29481
rect 19890 29407 19946 29416
rect 19904 29170 19932 29407
rect 20088 29170 20116 30126
rect 20180 30104 20208 30892
rect 20350 30832 20406 30841
rect 20350 30767 20406 30776
rect 20364 30598 20392 30767
rect 20352 30592 20404 30598
rect 20350 30560 20352 30569
rect 20404 30560 20406 30569
rect 20350 30495 20406 30504
rect 20258 30424 20314 30433
rect 20258 30359 20314 30368
rect 20442 30424 20498 30433
rect 20442 30359 20498 30368
rect 20272 30172 20300 30359
rect 20456 30326 20484 30359
rect 20640 30326 20668 32302
rect 21088 32224 21140 32230
rect 21088 32166 21140 32172
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20718 31104 20774 31113
rect 20718 31039 20774 31048
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20628 30320 20680 30326
rect 20732 30297 20760 31039
rect 20628 30262 20680 30268
rect 20718 30288 20774 30297
rect 20718 30223 20774 30232
rect 20272 30144 20760 30172
rect 20180 30076 20576 30104
rect 20155 29948 20463 29957
rect 20155 29946 20161 29948
rect 20217 29946 20241 29948
rect 20297 29946 20321 29948
rect 20377 29946 20401 29948
rect 20457 29946 20463 29948
rect 20217 29894 20219 29946
rect 20399 29894 20401 29946
rect 20155 29892 20161 29894
rect 20217 29892 20241 29894
rect 20297 29892 20321 29894
rect 20377 29892 20401 29894
rect 20457 29892 20463 29894
rect 20155 29883 20463 29892
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20260 29776 20312 29782
rect 20260 29718 20312 29724
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 20180 29050 20208 29514
rect 19904 29022 20208 29050
rect 20272 29034 20300 29718
rect 20364 29578 20392 29786
rect 20352 29572 20404 29578
rect 20352 29514 20404 29520
rect 20444 29572 20496 29578
rect 20444 29514 20496 29520
rect 20456 29306 20484 29514
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20456 29170 20484 29242
rect 20444 29164 20496 29170
rect 20444 29106 20496 29112
rect 20260 29028 20312 29034
rect 19800 27940 19852 27946
rect 19800 27882 19852 27888
rect 19798 27704 19854 27713
rect 19798 27639 19854 27648
rect 19628 27560 19748 27588
rect 19628 27554 19656 27560
rect 19619 27526 19656 27554
rect 19619 27384 19647 27526
rect 19619 27356 19656 27384
rect 19628 26994 19656 27356
rect 19616 26988 19668 26994
rect 19812 26976 19840 27639
rect 19904 27470 19932 29022
rect 20260 28970 20312 28976
rect 20155 28860 20463 28869
rect 20155 28858 20161 28860
rect 20217 28858 20241 28860
rect 20297 28858 20321 28860
rect 20377 28858 20401 28860
rect 20457 28858 20463 28860
rect 20217 28806 20219 28858
rect 20399 28806 20401 28858
rect 20155 28804 20161 28806
rect 20217 28804 20241 28806
rect 20297 28804 20321 28806
rect 20377 28804 20401 28806
rect 20457 28804 20463 28806
rect 19982 28792 20038 28801
rect 20155 28795 20463 28804
rect 20548 28762 20576 30076
rect 20626 30016 20682 30025
rect 20626 29951 20682 29960
rect 20640 29714 20668 29951
rect 20732 29850 20760 30144
rect 20720 29844 20772 29850
rect 20824 29832 20852 31758
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20994 30560 21050 30569
rect 20916 30297 20944 30534
rect 20994 30495 21050 30504
rect 20902 30288 20958 30297
rect 20902 30223 20958 30232
rect 20824 29804 20944 29832
rect 20720 29786 20772 29792
rect 20810 29744 20866 29753
rect 20628 29708 20680 29714
rect 20810 29679 20866 29688
rect 20628 29650 20680 29656
rect 20720 29640 20772 29646
rect 20626 29608 20682 29617
rect 20720 29582 20772 29588
rect 20626 29543 20682 29552
rect 20640 29306 20668 29543
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 20732 29170 20760 29582
rect 20824 29345 20852 29679
rect 20810 29336 20866 29345
rect 20810 29271 20866 29280
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20626 28928 20682 28937
rect 20626 28863 20682 28872
rect 19982 28727 20038 28736
rect 20260 28756 20312 28762
rect 19996 28558 20024 28727
rect 20260 28698 20312 28704
rect 20536 28756 20588 28762
rect 20536 28698 20588 28704
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 20272 28370 20300 28698
rect 20350 28656 20406 28665
rect 20350 28591 20406 28600
rect 20444 28620 20496 28626
rect 20364 28490 20392 28591
rect 20640 28608 20668 28863
rect 20718 28792 20774 28801
rect 20718 28727 20774 28736
rect 20732 28626 20760 28727
rect 20824 28626 20852 29271
rect 20496 28580 20668 28608
rect 20720 28620 20772 28626
rect 20444 28562 20496 28568
rect 20720 28562 20772 28568
rect 20812 28620 20864 28626
rect 20812 28562 20864 28568
rect 20916 28529 20944 29804
rect 21008 29578 21036 30495
rect 20996 29572 21048 29578
rect 20996 29514 21048 29520
rect 20994 29472 21050 29481
rect 20994 29407 21050 29416
rect 20718 28520 20774 28529
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 20444 28484 20496 28490
rect 20444 28426 20496 28432
rect 20548 28478 20718 28506
rect 20456 28370 20484 28426
rect 20272 28342 20484 28370
rect 20548 28200 20576 28478
rect 20718 28455 20774 28464
rect 20902 28520 20958 28529
rect 20902 28455 20958 28464
rect 20720 28416 20772 28422
rect 20720 28358 20772 28364
rect 20812 28416 20864 28422
rect 21008 28404 21036 29407
rect 21100 29220 21128 32166
rect 21192 32026 21220 32302
rect 21180 32020 21232 32026
rect 21180 31962 21232 31968
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 21192 31414 21220 31758
rect 21180 31408 21232 31414
rect 21180 31350 21232 31356
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 21192 29782 21220 30126
rect 21180 29776 21232 29782
rect 21180 29718 21232 29724
rect 21284 29714 21312 32506
rect 21456 32496 21508 32502
rect 21362 32464 21418 32473
rect 21456 32438 21508 32444
rect 21362 32399 21418 32408
rect 21376 30870 21404 32399
rect 21468 31482 21496 32438
rect 21548 32292 21600 32298
rect 21548 32234 21600 32240
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21364 30864 21416 30870
rect 21364 30806 21416 30812
rect 21456 30864 21508 30870
rect 21456 30806 21508 30812
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 21376 29850 21404 30330
rect 21364 29844 21416 29850
rect 21364 29786 21416 29792
rect 21468 29753 21496 30806
rect 21560 30433 21588 32234
rect 21546 30424 21602 30433
rect 21546 30359 21602 30368
rect 21548 30116 21600 30122
rect 21548 30058 21600 30064
rect 21454 29744 21510 29753
rect 21272 29708 21324 29714
rect 21454 29679 21510 29688
rect 21272 29650 21324 29656
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21192 29322 21220 29582
rect 21468 29481 21496 29582
rect 21454 29472 21510 29481
rect 21454 29407 21510 29416
rect 21560 29322 21588 30058
rect 21192 29294 21312 29322
rect 21100 29192 21220 29220
rect 21088 29028 21140 29034
rect 21088 28970 21140 28976
rect 20812 28358 20864 28364
rect 20916 28376 21036 28404
rect 20180 28172 20576 28200
rect 20180 28064 20208 28172
rect 20167 28036 20208 28064
rect 20260 28076 20312 28082
rect 20076 28008 20128 28014
rect 19996 27968 20076 27996
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19892 27124 19944 27130
rect 19892 27066 19944 27072
rect 19616 26930 19668 26936
rect 19720 26948 19840 26976
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 19720 26738 19748 26948
rect 19798 26888 19854 26897
rect 19904 26874 19932 27066
rect 19854 26846 19932 26874
rect 19798 26823 19854 26832
rect 19892 26784 19944 26790
rect 19628 26625 19656 26726
rect 19720 26710 19833 26738
rect 19892 26726 19944 26732
rect 19614 26616 19670 26625
rect 19614 26551 19670 26560
rect 19616 26512 19668 26518
rect 19805 26500 19833 26710
rect 19805 26472 19840 26500
rect 19616 26454 19668 26460
rect 19628 25906 19656 26454
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19720 25922 19748 26318
rect 19812 26024 19840 26472
rect 19904 26314 19932 26726
rect 19996 26382 20024 27968
rect 20076 27950 20128 27956
rect 20167 27928 20195 28036
rect 20260 28018 20312 28024
rect 20536 28076 20588 28082
rect 20588 28036 20668 28064
rect 20536 28018 20588 28024
rect 20167 27900 20208 27928
rect 20180 27860 20208 27900
rect 20088 27832 20208 27860
rect 20272 27860 20300 28018
rect 20272 27832 20576 27860
rect 20088 27606 20116 27832
rect 20155 27772 20463 27781
rect 20155 27770 20161 27772
rect 20217 27770 20241 27772
rect 20297 27770 20321 27772
rect 20377 27770 20401 27772
rect 20457 27770 20463 27772
rect 20217 27718 20219 27770
rect 20399 27718 20401 27770
rect 20155 27716 20161 27718
rect 20217 27716 20241 27718
rect 20297 27716 20321 27718
rect 20377 27716 20401 27718
rect 20457 27716 20463 27718
rect 20155 27707 20463 27716
rect 20260 27668 20312 27674
rect 20312 27628 20392 27656
rect 20260 27610 20312 27616
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 20258 27568 20314 27577
rect 20258 27503 20314 27512
rect 20272 27470 20300 27503
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20168 27396 20220 27402
rect 20168 27338 20220 27344
rect 20180 27062 20208 27338
rect 20168 27056 20220 27062
rect 20168 26998 20220 27004
rect 20076 26784 20128 26790
rect 20364 26772 20392 27628
rect 20548 26858 20576 27832
rect 20640 26976 20668 28036
rect 20732 27538 20760 28358
rect 20824 28082 20852 28358
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20824 27849 20852 28018
rect 20916 28014 20944 28376
rect 20904 28008 20956 28014
rect 20904 27950 20956 27956
rect 20994 27976 21050 27985
rect 20994 27911 21050 27920
rect 20810 27840 20866 27849
rect 20810 27775 20866 27784
rect 20812 27668 20864 27674
rect 20812 27610 20864 27616
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20732 27334 20760 27474
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20640 26948 20760 26976
rect 20536 26852 20588 26858
rect 20536 26794 20588 26800
rect 20444 26784 20496 26790
rect 20364 26744 20444 26772
rect 20076 26726 20128 26732
rect 20444 26726 20496 26732
rect 20534 26752 20590 26761
rect 20088 26568 20116 26726
rect 20155 26684 20463 26693
rect 20534 26687 20590 26696
rect 20155 26682 20161 26684
rect 20217 26682 20241 26684
rect 20297 26682 20321 26684
rect 20377 26682 20401 26684
rect 20457 26682 20463 26684
rect 20217 26630 20219 26682
rect 20399 26630 20401 26682
rect 20155 26628 20161 26630
rect 20217 26628 20241 26630
rect 20297 26628 20321 26630
rect 20377 26628 20401 26630
rect 20457 26628 20463 26630
rect 20155 26619 20463 26628
rect 20548 26586 20576 26687
rect 20732 26625 20760 26948
rect 20718 26616 20774 26625
rect 20536 26580 20588 26586
rect 20088 26540 20484 26568
rect 20352 26444 20404 26450
rect 20272 26404 20352 26432
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 20076 26376 20128 26382
rect 20128 26336 20195 26364
rect 20272 26353 20300 26404
rect 20352 26386 20404 26392
rect 20076 26318 20128 26324
rect 20167 26330 20195 26336
rect 20258 26344 20314 26353
rect 19892 26308 19944 26314
rect 20167 26302 20208 26330
rect 19892 26250 19944 26256
rect 19812 25996 20116 26024
rect 19616 25900 19668 25906
rect 19720 25894 20024 25922
rect 20088 25906 20116 25996
rect 19616 25842 19668 25848
rect 19708 25832 19760 25838
rect 19536 25758 19656 25786
rect 19708 25774 19760 25780
rect 19798 25800 19854 25809
rect 19076 25622 19380 25650
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19076 24993 19104 25622
rect 19536 25480 19564 25638
rect 19168 25452 19564 25480
rect 19168 25362 19196 25452
rect 19338 25392 19394 25401
rect 19156 25356 19208 25362
rect 19338 25327 19340 25336
rect 19156 25298 19208 25304
rect 19392 25327 19394 25336
rect 19522 25392 19578 25401
rect 19522 25327 19578 25336
rect 19340 25298 19392 25304
rect 19536 25294 19564 25327
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19062 24984 19118 24993
rect 19062 24919 19118 24928
rect 19248 24880 19300 24886
rect 19168 24840 19248 24868
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18880 24744 18932 24750
rect 18932 24692 19012 24698
rect 18880 24686 19012 24692
rect 18892 24670 19012 24686
rect 18878 24576 18934 24585
rect 18878 24511 18934 24520
rect 18696 24336 18748 24342
rect 18748 24296 18828 24324
rect 18892 24313 18920 24511
rect 18696 24278 18748 24284
rect 18604 24200 18656 24206
rect 18656 24160 18736 24188
rect 18604 24142 18656 24148
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18616 22409 18644 23666
rect 18708 22642 18736 24160
rect 18800 22642 18828 24296
rect 18878 24304 18934 24313
rect 18878 24239 18934 24248
rect 18984 24206 19012 24670
rect 19168 24614 19196 24840
rect 19248 24822 19300 24828
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18602 22400 18658 22409
rect 18602 22335 18658 22344
rect 18786 22264 18842 22273
rect 18432 22222 18786 22250
rect 18786 22199 18842 22208
rect 18328 22160 18380 22166
rect 18420 22160 18472 22166
rect 18328 22102 18380 22108
rect 18418 22128 18420 22137
rect 18472 22128 18474 22137
rect 18892 22098 18920 24142
rect 18984 22642 19012 24142
rect 19062 24032 19118 24041
rect 19062 23967 19118 23976
rect 19076 23662 19104 23967
rect 19168 23798 19196 24278
rect 19260 24070 19288 24618
rect 19352 24206 19380 25162
rect 19444 25106 19472 25230
rect 19628 25226 19656 25758
rect 19616 25220 19668 25226
rect 19616 25162 19668 25168
rect 19720 25106 19748 25774
rect 19854 25758 19932 25786
rect 19798 25735 19854 25744
rect 19800 25696 19852 25702
rect 19800 25638 19852 25644
rect 19444 25078 19564 25106
rect 19430 24984 19486 24993
rect 19430 24919 19486 24928
rect 19444 24585 19472 24919
rect 19430 24576 19486 24585
rect 19430 24511 19486 24520
rect 19536 24449 19564 25078
rect 19628 25078 19748 25106
rect 19812 25106 19840 25638
rect 19904 25226 19932 25758
rect 19996 25430 20024 25894
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25809 20116 25842
rect 20074 25800 20130 25809
rect 20074 25735 20130 25744
rect 20180 25684 20208 26302
rect 20258 26279 20314 26288
rect 20272 25906 20300 26279
rect 20456 26024 20484 26540
rect 20718 26551 20774 26560
rect 20536 26522 20588 26528
rect 20628 26512 20680 26518
rect 20628 26454 20680 26460
rect 20456 25996 20576 26024
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20456 25770 20484 25842
rect 20444 25764 20496 25770
rect 20444 25706 20496 25712
rect 20088 25656 20208 25684
rect 19984 25424 20036 25430
rect 19984 25366 20036 25372
rect 20088 25265 20116 25656
rect 20155 25596 20463 25605
rect 20155 25594 20161 25596
rect 20217 25594 20241 25596
rect 20297 25594 20321 25596
rect 20377 25594 20401 25596
rect 20457 25594 20463 25596
rect 20217 25542 20219 25594
rect 20399 25542 20401 25594
rect 20155 25540 20161 25542
rect 20217 25540 20241 25542
rect 20297 25540 20321 25542
rect 20377 25540 20401 25542
rect 20457 25540 20463 25542
rect 20155 25531 20463 25540
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 20180 25276 20208 25434
rect 20548 25430 20576 25996
rect 20640 25770 20668 26454
rect 20824 25888 20852 27610
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20732 25860 20852 25888
rect 20628 25764 20680 25770
rect 20628 25706 20680 25712
rect 20444 25424 20496 25430
rect 20444 25366 20496 25372
rect 20536 25424 20588 25430
rect 20536 25366 20588 25372
rect 20352 25288 20404 25294
rect 20074 25256 20130 25265
rect 19892 25220 19944 25226
rect 20180 25248 20300 25276
rect 20074 25191 20130 25200
rect 19892 25162 19944 25168
rect 19812 25078 20208 25106
rect 19628 24585 19656 25078
rect 20180 24954 20208 25078
rect 20168 24948 20220 24954
rect 19720 24908 20024 24936
rect 19720 24750 19748 24908
rect 19996 24868 20024 24908
rect 20168 24890 20220 24896
rect 20076 24880 20128 24886
rect 19996 24840 20076 24868
rect 20076 24822 20128 24828
rect 19800 24812 19852 24818
rect 19800 24754 19852 24760
rect 19708 24744 19760 24750
rect 19708 24686 19760 24692
rect 19812 24614 19840 24754
rect 20168 24744 20220 24750
rect 19996 24704 20168 24732
rect 19708 24608 19760 24614
rect 19614 24576 19670 24585
rect 19708 24550 19760 24556
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19890 24576 19946 24585
rect 19614 24511 19670 24520
rect 19522 24440 19578 24449
rect 19522 24375 19578 24384
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 19524 24200 19576 24206
rect 19576 24160 19656 24188
rect 19524 24142 19576 24148
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19246 23760 19302 23769
rect 19246 23695 19302 23704
rect 19260 23662 19288 23695
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19076 23361 19104 23598
rect 19062 23352 19118 23361
rect 19062 23287 19118 23296
rect 19168 23050 19196 23598
rect 19352 23304 19380 24006
rect 19524 23724 19576 23730
rect 19444 23684 19524 23712
rect 19444 23497 19472 23684
rect 19524 23666 19576 23672
rect 19430 23488 19486 23497
rect 19430 23423 19486 23432
rect 19352 23276 19472 23304
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19064 23044 19116 23050
rect 19064 22986 19116 22992
rect 19156 23044 19208 23050
rect 19156 22986 19208 22992
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18418 22063 18474 22072
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18328 22024 18380 22030
rect 18248 21984 18328 22012
rect 18144 21966 18196 21972
rect 18328 21966 18380 21972
rect 17958 21927 17960 21936
rect 18012 21927 18014 21936
rect 17960 21898 18012 21904
rect 18064 21865 18092 21966
rect 18788 21956 18840 21962
rect 18788 21898 18840 21904
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18050 21856 18106 21865
rect 18050 21791 18106 21800
rect 18156 21814 18736 21842
rect 18156 21690 18184 21814
rect 18708 21729 18736 21814
rect 18234 21720 18290 21729
rect 18144 21684 18196 21690
rect 18234 21655 18236 21664
rect 18144 21626 18196 21632
rect 18288 21655 18290 21664
rect 18510 21720 18566 21729
rect 18694 21720 18750 21729
rect 18566 21678 18644 21706
rect 18510 21655 18566 21664
rect 18236 21626 18288 21632
rect 18340 21542 18552 21570
rect 18236 21480 18288 21486
rect 17866 21448 17922 21457
rect 17684 21412 17736 21418
rect 17684 21354 17736 21360
rect 17776 21412 17828 21418
rect 18340 21468 18368 21542
rect 18524 21486 18552 21542
rect 18288 21440 18368 21468
rect 18420 21480 18472 21486
rect 18236 21422 18288 21428
rect 18420 21422 18472 21428
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 17866 21383 17922 21392
rect 17776 21354 17828 21360
rect 17788 21078 17816 21354
rect 18432 21350 18460 21422
rect 18420 21344 18472 21350
rect 18616 21332 18644 21678
rect 18694 21655 18750 21664
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18708 21486 18736 21558
rect 18800 21486 18828 21898
rect 18892 21729 18920 21898
rect 18878 21720 18934 21729
rect 18878 21655 18934 21664
rect 18984 21554 19012 22578
rect 19076 21729 19104 22986
rect 19168 22234 19196 22986
rect 19352 22817 19380 23122
rect 19338 22808 19394 22817
rect 19338 22743 19394 22752
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 19260 22098 19288 22510
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19248 22092 19300 22098
rect 19168 22052 19248 22080
rect 19062 21720 19118 21729
rect 19062 21655 19118 21664
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18696 21480 18748 21486
rect 18696 21422 18748 21428
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18472 21304 18644 21332
rect 18420 21286 18472 21292
rect 18432 21221 18460 21286
rect 17868 21140 17920 21146
rect 18052 21140 18104 21146
rect 17920 21100 18052 21128
rect 17868 21082 17920 21088
rect 18052 21082 18104 21088
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 17776 21072 17828 21078
rect 17776 21014 17828 21020
rect 17592 21004 17644 21010
rect 17236 20964 17448 20992
rect 17512 20964 17592 20992
rect 17236 20890 17264 20964
rect 17420 20924 17448 20964
rect 17592 20946 17644 20952
rect 17880 20998 18368 21026
rect 16960 20862 17264 20890
rect 17314 20904 17370 20913
rect 16960 20602 16988 20862
rect 17420 20896 17467 20924
rect 17439 20890 17467 20896
rect 17682 20904 17738 20913
rect 17439 20862 17632 20890
rect 17314 20839 17370 20848
rect 17224 20800 17276 20806
rect 17052 20748 17224 20754
rect 17328 20788 17356 20839
rect 17328 20760 17448 20788
rect 17052 20742 17276 20748
rect 17052 20726 17264 20742
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17052 20482 17080 20726
rect 17420 20584 17448 20760
rect 17604 20754 17632 20862
rect 17880 20856 17908 20998
rect 18340 20942 18368 20998
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18328 20936 18380 20942
rect 18604 20936 18656 20942
rect 18328 20878 18380 20884
rect 18524 20896 18604 20924
rect 17682 20839 17684 20848
rect 17736 20839 17738 20848
rect 17684 20810 17736 20816
rect 17788 20828 17908 20856
rect 18144 20868 18196 20874
rect 17788 20754 17816 20828
rect 18144 20810 18196 20816
rect 18156 20777 18184 20810
rect 17604 20726 17816 20754
rect 18142 20768 18198 20777
rect 18142 20703 18198 20712
rect 17960 20596 18012 20602
rect 17420 20556 17960 20584
rect 17960 20538 18012 20544
rect 16868 20454 17080 20482
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 16764 20392 16816 20398
rect 17144 20346 17172 20402
rect 16816 20340 17172 20346
rect 16764 20334 17172 20340
rect 16212 20324 16264 20330
rect 16776 20318 17172 20334
rect 16212 20266 16264 20272
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16040 19718 16068 20198
rect 16224 19922 16252 20266
rect 17236 20244 17264 20470
rect 18248 20466 18276 20878
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18340 20534 18368 20742
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 17408 20460 17460 20466
rect 17960 20460 18012 20466
rect 17460 20420 17960 20448
rect 17408 20402 17460 20408
rect 17960 20402 18012 20408
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 17420 20330 18276 20346
rect 17408 20324 18276 20330
rect 17460 20318 18276 20324
rect 17408 20266 17460 20272
rect 18248 20262 18276 20318
rect 17144 20216 17264 20244
rect 17500 20256 17552 20262
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 15936 19712 15988 19718
rect 15842 19680 15898 19689
rect 15936 19654 15988 19660
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15842 19615 15898 19624
rect 15856 19378 15884 19615
rect 15948 19378 15976 19654
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15750 18864 15806 18873
rect 15660 18828 15712 18834
rect 15750 18799 15806 18808
rect 15660 18770 15712 18776
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15476 18420 15528 18426
rect 15948 18408 15976 18906
rect 16040 18698 16068 19654
rect 16118 19544 16174 19553
rect 16118 19479 16174 19488
rect 16224 19496 16252 19858
rect 17144 19854 17172 20216
rect 17500 20198 17552 20204
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 18052 20256 18104 20262
rect 18236 20256 18288 20262
rect 18052 20198 18104 20204
rect 18142 20224 18198 20233
rect 17512 20040 17540 20198
rect 17420 20012 17540 20040
rect 17420 19961 17448 20012
rect 17696 19972 17724 20198
rect 17406 19952 17462 19961
rect 17224 19916 17276 19922
rect 17696 19944 17816 19972
rect 17406 19887 17462 19896
rect 17224 19858 17276 19864
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 16762 19680 16818 19689
rect 16314 19612 16622 19621
rect 16762 19615 16818 19624
rect 16314 19610 16320 19612
rect 16376 19610 16400 19612
rect 16456 19610 16480 19612
rect 16536 19610 16560 19612
rect 16616 19610 16622 19612
rect 16376 19558 16378 19610
rect 16558 19558 16560 19610
rect 16314 19556 16320 19558
rect 16376 19556 16400 19558
rect 16456 19556 16480 19558
rect 16536 19556 16560 19558
rect 16616 19556 16622 19558
rect 16314 19547 16622 19556
rect 16776 19514 16804 19615
rect 16854 19544 16910 19553
rect 16764 19508 16816 19514
rect 16132 19258 16160 19479
rect 16224 19468 16528 19496
rect 16302 19408 16358 19417
rect 16302 19343 16304 19352
rect 16356 19343 16358 19352
rect 16304 19314 16356 19320
rect 16132 19230 16436 19258
rect 16132 18822 16344 18850
rect 16132 18766 16160 18822
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16212 18760 16264 18766
rect 16316 18748 16344 18822
rect 16408 18816 16436 19230
rect 16500 18884 16528 19468
rect 16854 19479 16910 19488
rect 16948 19508 17000 19514
rect 16764 19450 16816 19456
rect 16868 19394 16896 19479
rect 16948 19450 17000 19456
rect 16592 19366 16896 19394
rect 16592 19009 16620 19366
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16776 19009 16804 19246
rect 16856 19236 16908 19242
rect 16960 19224 16988 19450
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16908 19196 16988 19224
rect 16856 19178 16908 19184
rect 16578 19000 16634 19009
rect 16578 18935 16634 18944
rect 16762 19000 16818 19009
rect 16762 18935 16818 18944
rect 16500 18856 16804 18884
rect 16776 18816 16804 18856
rect 16408 18788 16620 18816
rect 16776 18788 16807 18816
rect 16316 18720 16528 18748
rect 16212 18702 16264 18708
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15476 18362 15528 18368
rect 15764 18380 15976 18408
rect 16026 18456 16082 18465
rect 16026 18391 16028 18400
rect 15200 17274 15252 17280
rect 15304 17292 15424 17320
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14738 16416 14794 16425
rect 14738 16351 14794 16360
rect 14740 16244 14792 16250
rect 14568 16204 14688 16232
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14384 14346 14412 14486
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14384 14006 14412 14282
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14476 13938 14504 14350
rect 14568 13977 14596 16050
rect 14660 14940 14688 16204
rect 14740 16186 14792 16192
rect 14752 15162 14780 16186
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14660 14912 14780 14940
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14660 14414 14688 14758
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14554 13968 14610 13977
rect 14464 13932 14516 13938
rect 14554 13903 14610 13912
rect 14464 13874 14516 13880
rect 14752 13870 14780 14912
rect 14740 13864 14792 13870
rect 14738 13832 14740 13841
rect 14792 13832 14794 13841
rect 14738 13767 14794 13776
rect 14844 13462 14872 16526
rect 14936 15706 14964 17138
rect 15304 17134 15332 17292
rect 15488 17270 15516 18362
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15580 17746 15608 17818
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15120 16658 15148 16934
rect 15212 16726 15240 16934
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15028 16250 15056 16526
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14936 15314 14964 15642
rect 15028 15502 15056 16186
rect 15120 15706 15148 16594
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15212 16289 15240 16526
rect 15198 16280 15254 16289
rect 15198 16215 15254 16224
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15212 15609 15240 16050
rect 15304 16046 15332 16730
rect 15396 16289 15424 17138
rect 15488 16708 15516 17206
rect 15580 16776 15608 17546
rect 15672 17082 15700 18022
rect 15764 17921 15792 18380
rect 16080 18391 16082 18400
rect 16224 18408 16252 18702
rect 16500 18630 16528 18720
rect 16488 18624 16540 18630
rect 16592 18612 16620 18788
rect 16592 18584 16712 18612
rect 16488 18566 16540 18572
rect 16314 18524 16622 18533
rect 16314 18522 16320 18524
rect 16376 18522 16400 18524
rect 16456 18522 16480 18524
rect 16536 18522 16560 18524
rect 16616 18522 16622 18524
rect 16376 18470 16378 18522
rect 16558 18470 16560 18522
rect 16314 18468 16320 18470
rect 16376 18468 16400 18470
rect 16456 18468 16480 18470
rect 16536 18468 16560 18470
rect 16616 18468 16622 18470
rect 16314 18459 16622 18468
rect 16684 18442 16712 18584
rect 16779 18578 16807 18788
rect 16868 18766 16896 19178
rect 16946 19136 17002 19145
rect 16946 19071 17002 19080
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16779 18550 16896 18578
rect 16762 18456 16818 18465
rect 16684 18414 16762 18442
rect 16224 18380 16528 18408
rect 16762 18391 16818 18400
rect 16028 18362 16080 18368
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15750 17912 15806 17921
rect 15948 17882 15976 18022
rect 15750 17847 15806 17856
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16040 17762 16068 18226
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16132 17814 16160 18158
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 15764 17734 16068 17762
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 15764 17678 15792 17734
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 17377 15884 17614
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15842 17368 15898 17377
rect 15842 17303 15898 17312
rect 15750 17096 15806 17105
rect 15672 17054 15750 17082
rect 15750 17031 15806 17040
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15660 16992 15712 16998
rect 15856 16946 15884 17002
rect 15948 16969 15976 17546
rect 16040 17490 16068 17734
rect 16316 17678 16344 18022
rect 16408 17921 16436 18158
rect 16394 17912 16450 17921
rect 16394 17847 16450 17856
rect 16500 17785 16528 18380
rect 16868 18358 16896 18550
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16856 18352 16908 18358
rect 16960 18340 16988 19071
rect 17052 18465 17080 19314
rect 17144 19122 17172 19790
rect 17236 19378 17264 19858
rect 17684 19848 17736 19854
rect 17328 19796 17684 19802
rect 17328 19790 17736 19796
rect 17328 19774 17724 19790
rect 17328 19446 17356 19774
rect 17408 19712 17460 19718
rect 17460 19660 17540 19666
rect 17408 19654 17540 19660
rect 17420 19638 17540 19654
rect 17512 19496 17540 19638
rect 17512 19468 17632 19496
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17420 19122 17448 19382
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17144 19094 17448 19122
rect 17144 18958 17356 18986
rect 17144 18902 17172 18958
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17222 18864 17278 18873
rect 17222 18799 17278 18808
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17038 18456 17094 18465
rect 17038 18391 17094 18400
rect 16960 18312 17080 18340
rect 16856 18294 16908 18300
rect 16592 17814 16620 18294
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16580 17808 16632 17814
rect 16486 17776 16542 17785
rect 16580 17750 16632 17756
rect 16486 17711 16542 17720
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 17536 16264 17542
rect 16040 17462 16160 17490
rect 16212 17478 16264 17484
rect 16026 17368 16082 17377
rect 16026 17303 16082 17312
rect 16040 16998 16068 17303
rect 16028 16992 16080 16998
rect 15712 16940 15884 16946
rect 15660 16934 15884 16940
rect 15672 16918 15884 16934
rect 15934 16960 15990 16969
rect 16028 16934 16080 16940
rect 15934 16895 15990 16904
rect 15844 16788 15896 16794
rect 15580 16748 15700 16776
rect 15488 16680 15608 16708
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15382 16280 15438 16289
rect 15382 16215 15438 16224
rect 15488 16046 15516 16390
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15304 15745 15332 15982
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15290 15736 15346 15745
rect 15290 15671 15346 15680
rect 15198 15600 15254 15609
rect 15198 15535 15254 15544
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14936 15286 15056 15314
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 13648 12406 13768 12434
rect 13924 12406 14320 12434
rect 13740 12374 13768 12406
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12473 9276 12781 9285
rect 12473 9274 12479 9276
rect 12535 9274 12559 9276
rect 12615 9274 12639 9276
rect 12695 9274 12719 9276
rect 12775 9274 12781 9276
rect 12535 9222 12537 9274
rect 12717 9222 12719 9274
rect 12473 9220 12479 9222
rect 12535 9220 12559 9222
rect 12615 9220 12639 9222
rect 12695 9220 12719 9222
rect 12775 9220 12781 9222
rect 12473 9211 12781 9220
rect 14292 8430 14320 12406
rect 14936 12170 14964 14826
rect 15028 14385 15056 15286
rect 15396 15162 15424 15914
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15450 15516 15846
rect 15580 15638 15608 16680
rect 15672 16454 15700 16748
rect 15844 16730 15896 16736
rect 15660 16448 15712 16454
rect 15856 16425 15884 16730
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15660 16390 15712 16396
rect 15842 16416 15898 16425
rect 15842 16351 15898 16360
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15488 15422 15608 15450
rect 15672 15434 15700 15982
rect 15580 15366 15608 15422
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15014 14376 15070 14385
rect 15014 14311 15070 14320
rect 14924 12164 14976 12170
rect 14924 12106 14976 12112
rect 15120 11558 15148 15030
rect 15212 14890 15240 15098
rect 15580 15026 15608 15302
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15212 13530 15240 13942
rect 15304 13530 15332 14962
rect 15396 13734 15424 14962
rect 15474 14648 15530 14657
rect 15474 14583 15476 14592
rect 15528 14583 15530 14592
rect 15476 14554 15528 14560
rect 15568 14340 15620 14346
rect 15672 14328 15700 15030
rect 15620 14300 15700 14328
rect 15568 14282 15620 14288
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15672 12617 15700 13874
rect 15658 12608 15714 12617
rect 15658 12543 15714 12552
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15764 10441 15792 16050
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15856 15910 15884 15982
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15948 15706 15976 16526
rect 16040 16454 16068 16526
rect 16028 16448 16080 16454
rect 16026 16416 16028 16425
rect 16080 16416 16082 16425
rect 16026 16351 16082 16360
rect 16132 16266 16160 17462
rect 16224 16794 16252 17478
rect 16314 17436 16622 17445
rect 16314 17434 16320 17436
rect 16376 17434 16400 17436
rect 16456 17434 16480 17436
rect 16536 17434 16560 17436
rect 16616 17434 16622 17436
rect 16376 17382 16378 17434
rect 16558 17382 16560 17434
rect 16314 17380 16320 17382
rect 16376 17380 16400 17382
rect 16456 17380 16480 17382
rect 16536 17380 16560 17382
rect 16616 17380 16622 17382
rect 16314 17371 16622 17380
rect 16684 17202 16712 17818
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16488 17128 16540 17134
rect 16580 17128 16632 17134
rect 16488 17070 16540 17076
rect 16578 17096 16580 17105
rect 16632 17096 16634 17105
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16040 16238 16160 16266
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15856 14822 15884 15642
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15856 14113 15884 14282
rect 15948 14249 15976 15506
rect 16040 14260 16068 16238
rect 16224 15978 16252 16526
rect 16500 16454 16528 17070
rect 16578 17031 16634 17040
rect 16684 16590 16712 17138
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16488 16448 16540 16454
rect 16592 16436 16620 16526
rect 16592 16408 16712 16436
rect 16776 16425 16804 17546
rect 16488 16390 16540 16396
rect 16314 16348 16622 16357
rect 16314 16346 16320 16348
rect 16376 16346 16400 16348
rect 16456 16346 16480 16348
rect 16536 16346 16560 16348
rect 16616 16346 16622 16348
rect 16376 16294 16378 16346
rect 16558 16294 16560 16346
rect 16314 16292 16320 16294
rect 16376 16292 16400 16294
rect 16456 16292 16480 16294
rect 16536 16292 16560 16294
rect 16616 16292 16622 16294
rect 16314 16283 16622 16292
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16120 15904 16172 15910
rect 16408 15858 16436 16186
rect 16684 16046 16712 16408
rect 16762 16416 16818 16425
rect 16762 16351 16818 16360
rect 16868 16250 16896 17818
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16960 17513 16988 17546
rect 16946 17504 17002 17513
rect 16946 17439 17002 17448
rect 16946 17368 17002 17377
rect 16946 17303 16948 17312
rect 17000 17303 17002 17312
rect 16948 17274 17000 17280
rect 17052 17066 17080 18312
rect 17144 17513 17172 18634
rect 17236 18601 17264 18799
rect 17222 18592 17278 18601
rect 17222 18527 17278 18536
rect 17328 18442 17356 18958
rect 17420 18766 17448 19094
rect 17512 18970 17540 19314
rect 17604 19145 17632 19468
rect 17788 19310 17816 19944
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17880 19156 17908 20198
rect 18064 20097 18092 20198
rect 18236 20198 18288 20204
rect 18142 20159 18198 20168
rect 18050 20088 18106 20097
rect 18050 20023 18106 20032
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17972 19786 18000 19926
rect 18156 19854 18184 20159
rect 18234 20088 18290 20097
rect 18234 20023 18236 20032
rect 18288 20023 18290 20032
rect 18236 19994 18288 20000
rect 18234 19952 18290 19961
rect 18234 19887 18290 19896
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17972 19378 18000 19450
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17590 19136 17646 19145
rect 17590 19071 17646 19080
rect 17788 19128 17908 19156
rect 18144 19168 18196 19174
rect 18050 19136 18106 19145
rect 17682 19000 17738 19009
rect 17500 18964 17552 18970
rect 17788 18970 17816 19128
rect 18248 19145 18276 19887
rect 18340 19378 18368 20470
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18432 20233 18460 20402
rect 18418 20224 18474 20233
rect 18418 20159 18474 20168
rect 18418 20088 18474 20097
rect 18418 20023 18474 20032
rect 18432 19446 18460 20023
rect 18524 19718 18552 20896
rect 18604 20878 18656 20884
rect 18708 20330 18736 21082
rect 18788 21072 18840 21078
rect 19076 21060 19104 21655
rect 19168 21622 19196 22052
rect 19248 22034 19300 22040
rect 19352 21690 19380 22442
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 18788 21014 18840 21020
rect 18984 21032 19104 21060
rect 18800 20942 18828 21014
rect 18984 20992 19012 21032
rect 18892 20964 19012 20992
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18892 20641 18920 20964
rect 18878 20632 18934 20641
rect 18878 20567 18934 20576
rect 19156 20528 19208 20534
rect 19156 20470 19208 20476
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 18696 19984 18748 19990
rect 18616 19944 18696 19972
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18144 19110 18196 19116
rect 18234 19136 18290 19145
rect 18050 19071 18106 19080
rect 17682 18935 17738 18944
rect 17776 18964 17828 18970
rect 17500 18906 17552 18912
rect 17696 18766 17724 18935
rect 17776 18906 17828 18912
rect 17788 18766 17816 18906
rect 17868 18828 17920 18834
rect 17920 18788 18000 18816
rect 17868 18770 17920 18776
rect 17408 18760 17460 18766
rect 17684 18760 17736 18766
rect 17460 18720 17632 18748
rect 17408 18702 17460 18708
rect 17604 18442 17632 18720
rect 17684 18702 17736 18708
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17972 18612 18000 18788
rect 18064 18766 18092 19071
rect 18156 19009 18184 19110
rect 18234 19071 18290 19080
rect 18142 19000 18198 19009
rect 18142 18935 18198 18944
rect 18340 18902 18368 19178
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17972 18584 18092 18612
rect 17224 18420 17276 18426
rect 17328 18414 17448 18442
rect 17604 18414 17908 18442
rect 17224 18362 17276 18368
rect 17130 17504 17186 17513
rect 17130 17439 17186 17448
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 16425 16988 16526
rect 16946 16416 17002 16425
rect 16946 16351 17002 16360
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16120 15846 16172 15852
rect 16132 15638 16160 15846
rect 16316 15830 16436 15858
rect 16316 15706 16344 15830
rect 16394 15736 16450 15745
rect 16304 15700 16356 15706
rect 16488 15700 16540 15706
rect 16450 15680 16488 15688
rect 16394 15671 16488 15680
rect 16408 15660 16488 15671
rect 16304 15642 16356 15648
rect 16488 15642 16540 15648
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 15144 16252 15438
rect 16500 15434 16528 15642
rect 16592 15502 16620 15914
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16488 15428 16540 15434
rect 16488 15370 16540 15376
rect 16314 15260 16622 15269
rect 16314 15258 16320 15260
rect 16376 15258 16400 15260
rect 16456 15258 16480 15260
rect 16536 15258 16560 15260
rect 16616 15258 16622 15260
rect 16376 15206 16378 15258
rect 16558 15206 16560 15258
rect 16314 15204 16320 15206
rect 16376 15204 16400 15206
rect 16456 15204 16480 15206
rect 16536 15204 16560 15206
rect 16616 15204 16622 15206
rect 16314 15195 16622 15204
rect 16224 15116 16620 15144
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16132 14414 16160 14894
rect 16316 14482 16344 14894
rect 16500 14822 16528 14894
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16304 14340 16356 14346
rect 16592 14328 16620 15116
rect 16684 14822 16712 15846
rect 16776 15201 16804 16118
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16762 15192 16818 15201
rect 16762 15127 16818 15136
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 14414 16712 14758
rect 16762 14512 16818 14521
rect 16762 14447 16818 14456
rect 16776 14414 16804 14447
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16356 14300 16620 14328
rect 16304 14282 16356 14288
rect 16764 14272 16816 14278
rect 15934 14240 15990 14249
rect 16040 14232 16160 14260
rect 15934 14175 15990 14184
rect 15842 14104 15898 14113
rect 15842 14039 15898 14048
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15856 12986 15884 13330
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15948 11762 15976 14175
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 12481 16068 13330
rect 16026 12472 16082 12481
rect 16026 12407 16082 12416
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 16132 11354 16160 14232
rect 16764 14214 16816 14220
rect 16314 14172 16622 14181
rect 16314 14170 16320 14172
rect 16376 14170 16400 14172
rect 16456 14170 16480 14172
rect 16536 14170 16560 14172
rect 16616 14170 16622 14172
rect 16376 14118 16378 14170
rect 16558 14118 16560 14170
rect 16314 14116 16320 14118
rect 16376 14116 16400 14118
rect 16456 14116 16480 14118
rect 16536 14116 16560 14118
rect 16616 14116 16622 14118
rect 16314 14107 16622 14116
rect 16776 14074 16804 14214
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 13320 16264 13326
rect 16316 13297 16344 13466
rect 16408 13326 16436 13874
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16396 13320 16448 13326
rect 16212 13262 16264 13268
rect 16302 13288 16358 13297
rect 16224 12918 16252 13262
rect 16396 13262 16448 13268
rect 16302 13223 16358 13232
rect 16314 13084 16622 13093
rect 16314 13082 16320 13084
rect 16376 13082 16400 13084
rect 16456 13082 16480 13084
rect 16536 13082 16560 13084
rect 16616 13082 16622 13084
rect 16376 13030 16378 13082
rect 16558 13030 16560 13082
rect 16314 13028 16320 13030
rect 16376 13028 16400 13030
rect 16456 13028 16480 13030
rect 16536 13028 16560 13030
rect 16616 13028 16622 13030
rect 16314 13019 16622 13028
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16224 12442 16252 12854
rect 16684 12714 16712 13806
rect 16776 13161 16804 13806
rect 16762 13152 16818 13161
rect 16762 13087 16818 13096
rect 16868 13025 16896 15846
rect 17052 15706 17080 17002
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17144 16046 17172 16526
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17236 15910 17264 18362
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 17328 18068 17356 18294
rect 17420 18170 17448 18414
rect 17684 18352 17736 18358
rect 17736 18312 17816 18340
rect 17684 18294 17736 18300
rect 17684 18216 17736 18222
rect 17420 18142 17632 18170
rect 17684 18158 17736 18164
rect 17408 18080 17460 18086
rect 17328 18040 17408 18068
rect 17408 18022 17460 18028
rect 17604 17921 17632 18142
rect 17406 17912 17462 17921
rect 17406 17847 17462 17856
rect 17590 17912 17646 17921
rect 17590 17847 17646 17856
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17328 17377 17356 17614
rect 17314 17368 17370 17377
rect 17314 17303 17370 17312
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16960 14550 16988 15506
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 17052 14414 17080 14554
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16960 14249 16988 14350
rect 17144 14346 17172 15302
rect 17328 15194 17356 17303
rect 17420 17270 17448 17847
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17236 15166 17356 15194
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 16946 14240 17002 14249
rect 17236 14226 17264 15166
rect 17420 15026 17448 17070
rect 17512 16969 17540 17274
rect 17498 16960 17554 16969
rect 17498 16895 17554 16904
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17512 15609 17540 15914
rect 17604 15638 17632 17750
rect 17696 17542 17724 18158
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17788 17270 17816 18312
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16522 17724 16934
rect 17788 16833 17816 17206
rect 17880 17134 17908 18414
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 17972 17882 18000 18294
rect 18064 18154 18092 18584
rect 18156 18358 18184 18838
rect 18432 18834 18460 19110
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17960 17536 18012 17542
rect 18012 17496 18092 17524
rect 17960 17478 18012 17484
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17866 16960 17922 16969
rect 17866 16895 17922 16904
rect 17774 16824 17830 16833
rect 17774 16759 17830 16768
rect 17880 16708 17908 16895
rect 17788 16680 17908 16708
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17788 16232 17816 16680
rect 17972 16658 18000 17070
rect 17960 16652 18012 16658
rect 17880 16612 17960 16640
rect 17880 16250 17908 16612
rect 17960 16594 18012 16600
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17696 16204 17816 16232
rect 17868 16244 17920 16250
rect 17696 15910 17724 16204
rect 17868 16186 17920 16192
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17592 15632 17644 15638
rect 17498 15600 17554 15609
rect 17788 15609 17816 16050
rect 17592 15574 17644 15580
rect 17774 15600 17830 15609
rect 17498 15535 17554 15544
rect 17774 15535 17830 15544
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 17328 14618 17356 14826
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17512 14521 17540 15098
rect 17498 14512 17554 14521
rect 17498 14447 17554 14456
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 16946 14175 17002 14184
rect 17144 14198 17264 14226
rect 16946 14104 17002 14113
rect 16946 14039 17002 14048
rect 16960 13462 16988 14039
rect 17144 13938 17172 14198
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17236 13841 17264 13942
rect 17328 13920 17356 14350
rect 17512 13977 17540 14350
rect 17498 13968 17554 13977
rect 17408 13932 17460 13938
rect 17328 13892 17408 13920
rect 17222 13832 17278 13841
rect 17222 13767 17278 13776
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16854 13016 16910 13025
rect 16854 12951 16910 12960
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16314 11996 16622 12005
rect 16314 11994 16320 11996
rect 16376 11994 16400 11996
rect 16456 11994 16480 11996
rect 16536 11994 16560 11996
rect 16616 11994 16622 11996
rect 16376 11942 16378 11994
rect 16558 11942 16560 11994
rect 16314 11940 16320 11942
rect 16376 11940 16400 11942
rect 16456 11940 16480 11942
rect 16536 11940 16560 11942
rect 16616 11940 16622 11942
rect 16314 11931 16622 11940
rect 16960 11626 16988 13194
rect 17052 12442 17080 13262
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17052 12238 17080 12378
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17052 11830 17080 12174
rect 17328 12102 17356 13892
rect 17498 13903 17554 13912
rect 17408 13874 17460 13880
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 17420 11558 17448 12242
rect 17604 11694 17632 15370
rect 17788 15065 17816 15535
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17774 15056 17830 15065
rect 17880 15026 17908 15302
rect 17774 14991 17830 15000
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17696 12442 17724 14894
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17788 12850 17816 14758
rect 17866 14512 17922 14521
rect 17866 14447 17868 14456
rect 17920 14447 17922 14456
rect 17868 14418 17920 14424
rect 17880 13938 17908 14418
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17972 13161 18000 16458
rect 18064 16114 18092 17496
rect 18156 16998 18184 18294
rect 18340 17649 18368 18362
rect 18524 17649 18552 19654
rect 18616 19310 18644 19944
rect 18696 19926 18748 19932
rect 18694 19816 18750 19825
rect 18694 19751 18696 19760
rect 18748 19751 18750 19760
rect 18696 19722 18748 19728
rect 18800 19689 18828 20266
rect 18892 19825 18920 20266
rect 18972 19848 19024 19854
rect 18878 19816 18934 19825
rect 19168 19825 19196 20470
rect 19260 20466 19288 21354
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19260 19961 19288 20402
rect 19246 19952 19302 19961
rect 19246 19887 19302 19896
rect 18972 19790 19024 19796
rect 19154 19816 19210 19825
rect 18878 19751 18934 19760
rect 18984 19689 19012 19790
rect 19352 19802 19380 21490
rect 19444 21418 19472 23276
rect 19524 23248 19576 23254
rect 19524 23190 19576 23196
rect 19536 23118 19564 23190
rect 19524 23112 19576 23118
rect 19524 23054 19576 23060
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19536 22438 19564 22510
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19536 22166 19564 22374
rect 19524 22160 19576 22166
rect 19524 22102 19576 22108
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 19154 19751 19210 19760
rect 19260 19774 19380 19802
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 18786 19680 18842 19689
rect 18786 19615 18842 19624
rect 18970 19680 19026 19689
rect 19260 19666 19288 19774
rect 18970 19615 19026 19624
rect 19076 19638 19288 19666
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 18786 19544 18842 19553
rect 18786 19479 18842 19488
rect 18880 19508 18932 19514
rect 18694 19408 18750 19417
rect 18800 19378 18828 19479
rect 18880 19450 18932 19456
rect 18694 19343 18750 19352
rect 18788 19372 18840 19378
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18326 17640 18382 17649
rect 18326 17575 18382 17584
rect 18510 17640 18566 17649
rect 18510 17575 18566 17584
rect 18236 17536 18288 17542
rect 18708 17490 18736 19343
rect 18788 19314 18840 19320
rect 18800 18766 18828 19314
rect 18892 18850 18920 19450
rect 19076 19242 19104 19638
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19168 19417 19196 19450
rect 19154 19408 19210 19417
rect 19154 19343 19210 19352
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 19168 19145 19196 19246
rect 19352 19224 19380 19654
rect 19260 19196 19380 19224
rect 19154 19136 19210 19145
rect 19154 19071 19210 19080
rect 18892 18822 19104 18850
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 18630 18920 18702
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18236 17478 18288 17484
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18050 15056 18106 15065
rect 18050 14991 18106 15000
rect 18064 14793 18092 14991
rect 18050 14784 18106 14793
rect 18050 14719 18106 14728
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18064 14482 18092 14554
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17958 13152 18014 13161
rect 17958 13087 18014 13096
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 17328 11218 17356 11494
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 16314 10908 16622 10917
rect 16314 10906 16320 10908
rect 16376 10906 16400 10908
rect 16456 10906 16480 10908
rect 16536 10906 16560 10908
rect 16616 10906 16622 10908
rect 16376 10854 16378 10906
rect 16558 10854 16560 10906
rect 16314 10852 16320 10854
rect 16376 10852 16400 10854
rect 16456 10852 16480 10854
rect 16536 10852 16560 10854
rect 16616 10852 16622 10854
rect 16314 10843 16622 10852
rect 17696 10470 17724 12038
rect 17774 11928 17830 11937
rect 17774 11863 17776 11872
rect 17828 11863 17830 11872
rect 17776 11834 17828 11840
rect 17972 11830 18000 12582
rect 18064 12238 18092 13874
rect 18156 12918 18184 16186
rect 18248 15881 18276 17478
rect 18616 17462 18736 17490
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18340 16998 18368 17206
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18328 16992 18380 16998
rect 18432 16969 18460 17070
rect 18328 16934 18380 16940
rect 18418 16960 18474 16969
rect 18340 16114 18368 16934
rect 18418 16895 18474 16904
rect 18418 16280 18474 16289
rect 18418 16215 18474 16224
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18340 15978 18368 16050
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18234 15872 18290 15881
rect 18234 15807 18290 15816
rect 18234 15736 18290 15745
rect 18234 15671 18290 15680
rect 18248 14618 18276 15671
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18248 14414 18276 14554
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18248 12850 18276 14010
rect 18340 13977 18368 15098
rect 18432 14521 18460 16215
rect 18524 15910 18552 17070
rect 18512 15904 18564 15910
rect 18616 15881 18644 17462
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18892 16250 18920 16662
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18512 15846 18564 15852
rect 18602 15872 18658 15881
rect 18602 15807 18658 15816
rect 18708 15434 18736 15982
rect 18878 15736 18934 15745
rect 18984 15706 19012 17274
rect 19076 16998 19104 18822
rect 19260 18816 19288 19196
rect 19338 19136 19394 19145
rect 19338 19071 19394 19080
rect 19352 18970 19380 19071
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19260 18788 19334 18816
rect 19306 18680 19334 18788
rect 19260 18652 19334 18680
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 19062 16280 19118 16289
rect 19168 16250 19196 18226
rect 19260 17746 19288 18652
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19352 17678 19380 18294
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19352 17218 19380 17614
rect 19444 17338 19472 19790
rect 19536 19009 19564 21898
rect 19628 21729 19656 24160
rect 19720 24070 19748 24550
rect 19890 24511 19946 24520
rect 19798 24440 19854 24449
rect 19798 24375 19854 24384
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19706 23896 19762 23905
rect 19706 23831 19762 23840
rect 19720 23361 19748 23831
rect 19812 23798 19840 24375
rect 19904 24324 19932 24511
rect 19996 24449 20024 24704
rect 20168 24686 20220 24692
rect 20272 24596 20300 25248
rect 20352 25230 20404 25236
rect 20364 24993 20392 25230
rect 20350 24984 20406 24993
rect 20350 24919 20406 24928
rect 20456 24854 20484 25366
rect 20732 25242 20760 25860
rect 20812 25764 20864 25770
rect 20812 25706 20864 25712
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20640 25214 20760 25242
rect 20548 24954 20576 25162
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20456 24826 20576 24854
rect 20088 24568 20300 24596
rect 19982 24440 20038 24449
rect 19982 24375 20038 24384
rect 20088 24392 20116 24568
rect 20155 24508 20463 24517
rect 20155 24506 20161 24508
rect 20217 24506 20241 24508
rect 20297 24506 20321 24508
rect 20377 24506 20401 24508
rect 20457 24506 20463 24508
rect 20217 24454 20219 24506
rect 20399 24454 20401 24506
rect 20155 24452 20161 24454
rect 20217 24452 20241 24454
rect 20297 24452 20321 24454
rect 20377 24452 20401 24454
rect 20457 24452 20463 24454
rect 20155 24443 20463 24452
rect 20352 24404 20404 24410
rect 20088 24364 20208 24392
rect 19904 24296 20116 24324
rect 20088 24206 20116 24296
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19800 23792 19852 23798
rect 19904 23764 19932 24006
rect 19800 23734 19852 23740
rect 19898 23758 19950 23764
rect 19898 23700 19950 23706
rect 19996 23610 20024 24142
rect 20180 23610 20208 24364
rect 20352 24346 20404 24352
rect 20260 24200 20312 24206
rect 20260 24142 20312 24148
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19904 23582 20024 23610
rect 20088 23582 20208 23610
rect 20272 23594 20300 24142
rect 20260 23588 20312 23594
rect 19706 23352 19762 23361
rect 19706 23287 19762 23296
rect 19812 23118 19840 23530
rect 19800 23112 19852 23118
rect 19720 23072 19800 23100
rect 19720 22778 19748 23072
rect 19800 23054 19852 23060
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19706 22536 19762 22545
rect 19706 22471 19762 22480
rect 19720 22030 19748 22471
rect 19812 22409 19840 22714
rect 19798 22400 19854 22409
rect 19798 22335 19854 22344
rect 19904 22250 19932 23582
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 19996 22642 20024 23258
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19996 22506 20024 22578
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 20088 22438 20116 23582
rect 20260 23530 20312 23536
rect 20364 23508 20392 24346
rect 20548 23644 20576 24826
rect 20640 23866 20668 25214
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20548 23616 20668 23644
rect 20364 23497 20576 23508
rect 20364 23488 20590 23497
rect 20364 23480 20534 23488
rect 20155 23420 20463 23429
rect 20534 23423 20590 23432
rect 20155 23418 20161 23420
rect 20217 23418 20241 23420
rect 20297 23418 20321 23420
rect 20377 23418 20401 23420
rect 20457 23418 20463 23420
rect 20217 23366 20219 23418
rect 20399 23366 20401 23418
rect 20155 23364 20161 23366
rect 20217 23364 20241 23366
rect 20297 23364 20321 23366
rect 20377 23364 20401 23366
rect 20457 23364 20463 23366
rect 20155 23355 20463 23364
rect 20640 23304 20668 23616
rect 20364 23276 20668 23304
rect 20364 23186 20392 23276
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20364 22710 20392 23122
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20456 22556 20484 23054
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20456 22528 20576 22556
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20155 22332 20463 22341
rect 20155 22330 20161 22332
rect 20217 22330 20241 22332
rect 20297 22330 20321 22332
rect 20377 22330 20401 22332
rect 20457 22330 20463 22332
rect 20217 22278 20219 22330
rect 20399 22278 20401 22330
rect 20155 22276 20161 22278
rect 20217 22276 20241 22278
rect 20297 22276 20321 22278
rect 20377 22276 20401 22278
rect 20457 22276 20463 22278
rect 19812 22222 19932 22250
rect 19982 22264 20038 22273
rect 20155 22267 20463 22276
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19812 21876 19840 22222
rect 20548 22216 20576 22528
rect 20038 22208 20576 22216
rect 19982 22199 20576 22208
rect 19996 22188 20576 22199
rect 19720 21848 19840 21876
rect 19614 21720 19670 21729
rect 19614 21655 19670 21664
rect 19628 20330 19656 21655
rect 19720 20788 19748 21848
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19812 20942 19840 21422
rect 19904 20942 19932 21626
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19996 21321 20024 21558
rect 19982 21312 20038 21321
rect 19982 21247 20038 21256
rect 20534 21312 20590 21321
rect 20155 21244 20463 21253
rect 20534 21247 20590 21256
rect 20155 21242 20161 21244
rect 20217 21242 20241 21244
rect 20297 21242 20321 21244
rect 20377 21242 20401 21244
rect 20457 21242 20463 21244
rect 20217 21190 20219 21242
rect 20399 21190 20401 21242
rect 20155 21188 20161 21190
rect 20217 21188 20241 21190
rect 20297 21188 20321 21190
rect 20377 21188 20401 21190
rect 20457 21188 20463 21190
rect 20155 21179 20463 21188
rect 19984 21140 20036 21146
rect 20548 21128 20576 21247
rect 20036 21100 20576 21128
rect 19984 21082 20036 21088
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19892 20936 19944 20942
rect 20640 20890 20668 22918
rect 20732 22642 20760 25094
rect 20824 23254 20852 25706
rect 20916 25294 20944 27270
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20732 22234 20760 22578
rect 20916 22545 20944 25230
rect 21008 25226 21036 27911
rect 21100 27577 21128 28970
rect 21192 28490 21220 29192
rect 21180 28484 21232 28490
rect 21180 28426 21232 28432
rect 21180 28212 21232 28218
rect 21180 28154 21232 28160
rect 21192 27656 21220 28154
rect 21284 27946 21312 29294
rect 21376 29294 21588 29322
rect 21376 28422 21404 29294
rect 21456 29232 21508 29238
rect 21456 29174 21508 29180
rect 21546 29200 21602 29209
rect 21468 28490 21496 29174
rect 21546 29135 21602 29144
rect 21560 28762 21588 29135
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21272 27668 21324 27674
rect 21192 27628 21272 27656
rect 21272 27610 21324 27616
rect 21086 27568 21142 27577
rect 21362 27568 21418 27577
rect 21272 27532 21324 27538
rect 21086 27503 21142 27512
rect 21192 27492 21272 27520
rect 21088 27464 21140 27470
rect 21086 27432 21088 27441
rect 21140 27432 21142 27441
rect 21086 27367 21142 27376
rect 21192 27112 21220 27492
rect 21362 27503 21418 27512
rect 21272 27474 21324 27480
rect 21272 27396 21324 27402
rect 21272 27338 21324 27344
rect 21100 27084 21220 27112
rect 20996 25220 21048 25226
rect 21100 25208 21128 27084
rect 21178 27024 21234 27033
rect 21178 26959 21234 26968
rect 21192 26518 21220 26959
rect 21180 26512 21232 26518
rect 21284 26489 21312 27338
rect 21376 27130 21404 27503
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 21468 26994 21496 28426
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 21560 27849 21588 28358
rect 21652 28082 21680 32710
rect 21824 31680 21876 31686
rect 21824 31622 21876 31628
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 21640 28076 21692 28082
rect 21640 28018 21692 28024
rect 21546 27840 21602 27849
rect 21546 27775 21602 27784
rect 21638 27704 21694 27713
rect 21548 27668 21600 27674
rect 21638 27639 21640 27648
rect 21548 27610 21600 27616
rect 21692 27639 21694 27648
rect 21640 27610 21692 27616
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 21180 26454 21232 26460
rect 21270 26480 21326 26489
rect 21270 26415 21326 26424
rect 21376 26432 21404 26930
rect 21560 26926 21588 27610
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21548 26920 21600 26926
rect 21548 26862 21600 26868
rect 21652 26772 21680 27270
rect 21560 26744 21680 26772
rect 21376 26404 21494 26432
rect 21180 26376 21232 26382
rect 21178 26344 21180 26353
rect 21232 26344 21234 26353
rect 21178 26279 21234 26288
rect 21364 26240 21416 26246
rect 21178 26208 21234 26217
rect 21178 26143 21234 26152
rect 21362 26208 21364 26217
rect 21416 26208 21418 26217
rect 21362 26143 21418 26152
rect 21192 25498 21220 26143
rect 21466 26058 21494 26404
rect 21284 26030 21494 26058
rect 21284 25945 21312 26030
rect 21364 25968 21416 25974
rect 21270 25936 21326 25945
rect 21364 25910 21416 25916
rect 21270 25871 21326 25880
rect 21272 25832 21324 25838
rect 21376 25809 21404 25910
rect 21272 25774 21324 25780
rect 21362 25800 21418 25809
rect 21180 25492 21232 25498
rect 21180 25434 21232 25440
rect 21284 25362 21312 25774
rect 21560 25786 21588 26744
rect 21744 26432 21772 30602
rect 21836 28801 21864 31622
rect 22112 31414 22140 32914
rect 22480 32434 22508 34350
rect 23570 32736 23626 32745
rect 23570 32671 23626 32680
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 23584 32314 23612 32671
rect 23676 32434 23704 34350
rect 24584 33380 24636 33386
rect 24584 33322 24636 33328
rect 23996 32668 24304 32677
rect 23996 32666 24002 32668
rect 24058 32666 24082 32668
rect 24138 32666 24162 32668
rect 24218 32666 24242 32668
rect 24298 32666 24304 32668
rect 24058 32614 24060 32666
rect 24240 32614 24242 32666
rect 23996 32612 24002 32614
rect 24058 32612 24082 32614
rect 24138 32612 24162 32614
rect 24218 32612 24242 32614
rect 24298 32612 24304 32614
rect 23996 32603 24304 32612
rect 24596 32570 24624 33322
rect 24584 32564 24636 32570
rect 24584 32506 24636 32512
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23848 32428 23900 32434
rect 23848 32370 23900 32376
rect 23112 32292 23164 32298
rect 23584 32286 23704 32314
rect 23112 32234 23164 32240
rect 22376 32224 22428 32230
rect 22376 32166 22428 32172
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 21916 30116 21968 30122
rect 21916 30058 21968 30064
rect 21928 29782 21956 30058
rect 21916 29776 21968 29782
rect 21916 29718 21968 29724
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21822 28792 21878 28801
rect 21822 28727 21878 28736
rect 21824 28688 21876 28694
rect 21928 28676 21956 29582
rect 22020 29152 22048 31078
rect 22112 29850 22140 31214
rect 22204 30569 22232 31214
rect 22388 31210 22416 32166
rect 23124 32026 23152 32234
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23572 32224 23624 32230
rect 23572 32166 23624 32172
rect 22744 32020 22796 32026
rect 22744 31962 22796 31968
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 22650 31920 22706 31929
rect 22650 31855 22706 31864
rect 22376 31204 22428 31210
rect 22376 31146 22428 31152
rect 22468 31204 22520 31210
rect 22468 31146 22520 31152
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 22190 30560 22246 30569
rect 22190 30495 22246 30504
rect 22388 30258 22416 30670
rect 22376 30252 22428 30258
rect 22376 30194 22428 30200
rect 22192 30048 22244 30054
rect 22192 29990 22244 29996
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 22204 29753 22232 29990
rect 22190 29744 22246 29753
rect 22190 29679 22246 29688
rect 22284 29708 22336 29714
rect 22284 29650 22336 29656
rect 22192 29572 22244 29578
rect 22192 29514 22244 29520
rect 22020 29124 22094 29152
rect 22066 28948 22094 29124
rect 22204 29034 22232 29514
rect 22296 29306 22324 29650
rect 22374 29608 22430 29617
rect 22374 29543 22430 29552
rect 22388 29306 22416 29543
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 22376 29300 22428 29306
rect 22376 29242 22428 29248
rect 22296 29186 22324 29242
rect 22296 29158 22416 29186
rect 22192 29028 22244 29034
rect 22192 28970 22244 28976
rect 22284 29028 22336 29034
rect 22284 28970 22336 28976
rect 22066 28920 22140 28948
rect 22112 28914 22140 28920
rect 22112 28886 22232 28914
rect 22006 28792 22062 28801
rect 22006 28727 22008 28736
rect 22060 28727 22062 28736
rect 22008 28698 22060 28704
rect 21876 28648 21956 28676
rect 22204 28642 22232 28886
rect 21824 28630 21876 28636
rect 21836 28218 21864 28630
rect 22112 28614 22232 28642
rect 21916 28552 21968 28558
rect 22112 28506 22140 28614
rect 21916 28494 21968 28500
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 21824 28008 21876 28014
rect 21824 27950 21876 27956
rect 21836 27849 21864 27950
rect 21822 27840 21878 27849
rect 21822 27775 21878 27784
rect 21822 27568 21878 27577
rect 21822 27503 21878 27512
rect 21362 25735 21418 25744
rect 21468 25758 21588 25786
rect 21652 26404 21772 26432
rect 21364 25424 21416 25430
rect 21364 25366 21416 25372
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 21376 25265 21404 25366
rect 21362 25256 21418 25265
rect 21100 25180 21220 25208
rect 21362 25191 21418 25200
rect 20996 25162 21048 25168
rect 21086 24984 21142 24993
rect 20996 24948 21048 24954
rect 21086 24919 21142 24928
rect 20996 24890 21048 24896
rect 21008 24449 21036 24890
rect 21100 24750 21128 24919
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 20994 24440 21050 24449
rect 20994 24375 21050 24384
rect 21086 24304 21142 24313
rect 21086 24239 21142 24248
rect 20994 24168 21050 24177
rect 21100 24138 21128 24239
rect 20994 24103 21050 24112
rect 21088 24132 21140 24138
rect 21008 24018 21036 24103
rect 21088 24074 21140 24080
rect 21008 23990 21128 24018
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 20902 22536 20958 22545
rect 20902 22471 20958 22480
rect 20810 22400 20866 22409
rect 20810 22335 20866 22344
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20732 21010 20760 21354
rect 20824 21350 20852 22335
rect 21008 22234 21036 23734
rect 21100 23662 21128 23990
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 21086 23488 21142 23497
rect 21086 23423 21142 23432
rect 21100 22982 21128 23423
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 21192 22778 21220 25180
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21284 24138 21312 24618
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21284 23322 21312 23802
rect 21376 23798 21404 25094
rect 21468 24732 21496 25758
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21560 25158 21588 25434
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 21546 24984 21602 24993
rect 21652 24970 21680 26404
rect 21836 26330 21864 27503
rect 21928 26432 21956 28494
rect 22020 28478 22140 28506
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22020 27577 22048 28478
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22112 27985 22140 28358
rect 22204 28257 22232 28494
rect 22296 28422 22324 28970
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22190 28248 22246 28257
rect 22190 28183 22246 28192
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22284 28144 22336 28150
rect 22284 28086 22336 28092
rect 22098 27976 22154 27985
rect 22098 27911 22154 27920
rect 22204 27878 22232 28086
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22006 27568 22062 27577
rect 22296 27554 22324 28086
rect 22006 27503 22062 27512
rect 22112 27526 22324 27554
rect 22112 27452 22140 27526
rect 22020 27424 22140 27452
rect 22020 26586 22048 27424
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 22284 27396 22336 27402
rect 22284 27338 22336 27344
rect 22204 27112 22232 27338
rect 22296 27305 22324 27338
rect 22282 27296 22338 27305
rect 22388 27282 22416 29158
rect 22480 27577 22508 31146
rect 22664 31113 22692 31855
rect 22756 31482 22784 31962
rect 23124 31686 23152 31962
rect 23112 31680 23164 31686
rect 23112 31622 23164 31628
rect 22744 31476 22796 31482
rect 22744 31418 22796 31424
rect 22650 31104 22706 31113
rect 22650 31039 22706 31048
rect 22664 30326 22692 31039
rect 22652 30320 22704 30326
rect 22652 30262 22704 30268
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22572 29306 22600 29582
rect 22560 29300 22612 29306
rect 22560 29242 22612 29248
rect 22664 29084 22692 29990
rect 22756 29170 22784 31418
rect 23308 31113 23336 32166
rect 23478 31648 23534 31657
rect 23478 31583 23534 31592
rect 23294 31104 23350 31113
rect 23294 31039 23350 31048
rect 23020 30932 23072 30938
rect 23020 30874 23072 30880
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 22848 29782 22876 30670
rect 22928 30660 22980 30666
rect 22928 30602 22980 30608
rect 22940 30258 22968 30602
rect 23032 30598 23060 30874
rect 23204 30864 23256 30870
rect 23124 30824 23204 30852
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 23124 30394 23152 30824
rect 23204 30806 23256 30812
rect 23388 30796 23440 30802
rect 23388 30738 23440 30744
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 23112 30388 23164 30394
rect 23112 30330 23164 30336
rect 23204 30320 23256 30326
rect 23202 30288 23204 30297
rect 23256 30288 23258 30297
rect 22928 30252 22980 30258
rect 23202 30223 23258 30232
rect 22928 30194 22980 30200
rect 23020 30184 23072 30190
rect 23020 30126 23072 30132
rect 23112 30184 23164 30190
rect 23112 30126 23164 30132
rect 22928 30116 22980 30122
rect 22928 30058 22980 30064
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22940 29617 22968 30058
rect 22926 29608 22982 29617
rect 22926 29543 22982 29552
rect 22836 29504 22888 29510
rect 23032 29492 23060 30126
rect 23124 30054 23152 30126
rect 23112 30048 23164 30054
rect 23204 30048 23256 30054
rect 23112 29990 23164 29996
rect 23202 30016 23204 30025
rect 23256 30016 23258 30025
rect 23202 29951 23258 29960
rect 23308 29832 23336 30670
rect 22888 29464 23060 29492
rect 23216 29804 23336 29832
rect 22836 29446 22888 29452
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22572 29056 22692 29084
rect 22742 29064 22798 29073
rect 22572 28994 22600 29056
rect 22742 28999 22798 29008
rect 22572 28966 22692 28994
rect 22558 28928 22614 28937
rect 22558 28863 22614 28872
rect 22572 28558 22600 28863
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22558 28248 22614 28257
rect 22558 28183 22614 28192
rect 22572 27946 22600 28183
rect 22560 27940 22612 27946
rect 22560 27882 22612 27888
rect 22558 27840 22614 27849
rect 22558 27775 22614 27784
rect 22466 27568 22522 27577
rect 22466 27503 22522 27512
rect 22466 27296 22522 27305
rect 22388 27254 22466 27282
rect 22282 27231 22338 27240
rect 22466 27231 22522 27240
rect 22204 27084 22508 27112
rect 22374 27024 22430 27033
rect 22192 26988 22244 26994
rect 22374 26959 22430 26968
rect 22192 26930 22244 26936
rect 22100 26852 22152 26858
rect 22100 26794 22152 26800
rect 22112 26625 22140 26794
rect 22098 26616 22154 26625
rect 22008 26580 22060 26586
rect 22098 26551 22154 26560
rect 22008 26522 22060 26528
rect 22204 26450 22232 26930
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22296 26625 22324 26862
rect 22282 26616 22338 26625
rect 22282 26551 22338 26560
rect 22388 26489 22416 26959
rect 22374 26480 22430 26489
rect 22192 26444 22244 26450
rect 21928 26404 22140 26432
rect 21836 26302 22048 26330
rect 21916 26240 21968 26246
rect 21916 26182 21968 26188
rect 21732 25968 21784 25974
rect 21732 25910 21784 25916
rect 21822 25936 21878 25945
rect 21744 25838 21772 25910
rect 21822 25871 21878 25880
rect 21732 25832 21784 25838
rect 21732 25774 21784 25780
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 21744 25129 21772 25638
rect 21730 25120 21786 25129
rect 21730 25055 21786 25064
rect 21652 24942 21772 24970
rect 21546 24919 21602 24928
rect 21560 24868 21588 24919
rect 21560 24840 21680 24868
rect 21548 24744 21600 24750
rect 21468 24704 21548 24732
rect 21468 24410 21496 24704
rect 21548 24686 21600 24692
rect 21546 24440 21602 24449
rect 21456 24404 21508 24410
rect 21546 24375 21602 24384
rect 21456 24346 21508 24352
rect 21454 24032 21510 24041
rect 21454 23967 21510 23976
rect 21364 23792 21416 23798
rect 21468 23769 21496 23967
rect 21560 23866 21588 24375
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21364 23734 21416 23740
rect 21454 23760 21510 23769
rect 21454 23695 21510 23704
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 21362 23488 21418 23497
rect 21362 23423 21418 23432
rect 21272 23316 21324 23322
rect 21272 23258 21324 23264
rect 21376 23118 21404 23423
rect 21468 23186 21496 23598
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21284 22778 21312 23054
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21284 22681 21312 22714
rect 21270 22672 21326 22681
rect 21270 22607 21326 22616
rect 21088 22500 21140 22506
rect 21088 22442 21140 22448
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 21008 21622 21036 22034
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 20996 21412 21048 21418
rect 20916 21372 20996 21400
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 19892 20878 19944 20884
rect 19996 20862 20392 20890
rect 20548 20874 20668 20890
rect 19720 20760 19840 20788
rect 19812 20714 19840 20760
rect 19720 20686 19840 20714
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 20097 19656 20266
rect 19614 20088 19670 20097
rect 19720 20058 19748 20686
rect 19892 20528 19944 20534
rect 19996 20516 20024 20862
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 19944 20488 20024 20516
rect 19892 20470 19944 20476
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19892 20256 19944 20262
rect 19890 20224 19892 20233
rect 19944 20224 19946 20233
rect 19890 20159 19946 20168
rect 19614 20023 19670 20032
rect 19708 20052 19760 20058
rect 19760 20012 19932 20040
rect 19708 19994 19760 20000
rect 19904 19786 19932 20012
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19522 19000 19578 19009
rect 19628 18970 19656 19450
rect 19522 18935 19578 18944
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19720 18884 19748 19722
rect 19800 19712 19852 19718
rect 19852 19660 19932 19666
rect 19800 19654 19932 19660
rect 19812 19638 19932 19654
rect 19798 19544 19854 19553
rect 19798 19479 19854 19488
rect 19904 19496 19932 19638
rect 19719 18856 19748 18884
rect 19719 18850 19747 18856
rect 19628 18822 19747 18850
rect 19628 18766 19656 18822
rect 19616 18760 19668 18766
rect 19522 18728 19578 18737
rect 19616 18702 19668 18708
rect 19522 18663 19578 18672
rect 19536 17542 19564 18663
rect 19628 18290 19656 18702
rect 19812 18442 19840 19479
rect 19904 19468 19938 19496
rect 19910 19428 19938 19468
rect 19996 19446 20024 20266
rect 20088 19972 20116 20742
rect 20364 20244 20392 20862
rect 20536 20868 20668 20874
rect 20588 20862 20668 20868
rect 20536 20810 20588 20816
rect 20628 20800 20680 20806
rect 20824 20788 20852 20946
rect 20916 20913 20944 21372
rect 20996 21354 21048 21360
rect 21100 21321 21128 22442
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21192 22094 21220 22374
rect 21376 22137 21404 23054
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21362 22128 21418 22137
rect 21192 22066 21312 22094
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21086 21312 21142 21321
rect 21086 21247 21142 21256
rect 20902 20904 20958 20913
rect 20902 20839 20958 20848
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20680 20760 20852 20788
rect 20904 20800 20956 20806
rect 20628 20742 20680 20748
rect 20904 20742 20956 20748
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20364 20216 20576 20244
rect 20155 20156 20463 20165
rect 20155 20154 20161 20156
rect 20217 20154 20241 20156
rect 20297 20154 20321 20156
rect 20377 20154 20401 20156
rect 20457 20154 20463 20156
rect 20217 20102 20219 20154
rect 20399 20102 20401 20154
rect 20155 20100 20161 20102
rect 20217 20100 20241 20102
rect 20297 20100 20321 20102
rect 20377 20100 20401 20102
rect 20457 20100 20463 20102
rect 20155 20091 20463 20100
rect 20548 20040 20576 20216
rect 20626 20224 20682 20233
rect 20626 20159 20682 20168
rect 20456 20012 20576 20040
rect 20088 19944 20392 19972
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20074 19680 20130 19689
rect 20074 19615 20130 19624
rect 19904 19400 19938 19428
rect 19984 19440 20036 19446
rect 19904 19310 19932 19400
rect 19984 19382 20036 19388
rect 20088 19334 20116 19615
rect 19898 19304 19950 19310
rect 19898 19246 19950 19252
rect 19996 19306 20116 19334
rect 19890 19136 19946 19145
rect 19890 19071 19946 19080
rect 19910 18850 19938 19071
rect 19996 18970 20024 19306
rect 20272 19156 20300 19722
rect 20364 19310 20392 19944
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20088 19128 20300 19156
rect 20456 19156 20484 20012
rect 20640 19514 20668 20159
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20456 19145 20576 19156
rect 20456 19136 20590 19145
rect 20456 19128 20534 19136
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 20088 18850 20116 19128
rect 20155 19068 20463 19077
rect 20534 19071 20590 19080
rect 20155 19066 20161 19068
rect 20217 19066 20241 19068
rect 20297 19066 20321 19068
rect 20377 19066 20401 19068
rect 20457 19066 20463 19068
rect 20217 19014 20219 19066
rect 20399 19014 20401 19066
rect 20155 19012 20161 19014
rect 20217 19012 20241 19014
rect 20297 19012 20321 19014
rect 20377 19012 20401 19014
rect 20457 19012 20463 19014
rect 20155 19003 20463 19012
rect 20732 18850 20760 20470
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20824 19514 20852 20334
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20916 18970 20944 20742
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 19910 18822 20116 18850
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20456 18822 20760 18850
rect 19812 18414 20116 18442
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19628 17814 19656 18226
rect 19798 18048 19854 18057
rect 19798 17983 19854 17992
rect 19616 17808 19668 17814
rect 19616 17750 19668 17756
rect 19812 17678 19840 17983
rect 19904 17921 19932 18294
rect 19890 17912 19946 17921
rect 19890 17847 19946 17856
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19352 17190 19472 17218
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19062 16215 19118 16224
rect 19156 16244 19208 16250
rect 19076 16182 19104 16215
rect 19156 16186 19208 16192
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 18878 15671 18934 15680
rect 18972 15700 19024 15706
rect 18892 15450 18920 15671
rect 18972 15642 19024 15648
rect 19076 15570 19104 15982
rect 19168 15638 19196 15982
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 18696 15428 18748 15434
rect 18892 15422 19012 15450
rect 18696 15370 18748 15376
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18616 14550 18644 14962
rect 18604 14544 18656 14550
rect 18418 14512 18474 14521
rect 18604 14486 18656 14492
rect 18418 14447 18474 14456
rect 18326 13968 18382 13977
rect 18326 13903 18382 13912
rect 18340 13870 18368 13903
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18340 12238 18368 13806
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18616 13682 18644 14486
rect 18708 13938 18736 15370
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18432 13394 18460 13670
rect 18616 13654 18736 13682
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18432 12918 18460 13330
rect 18708 13326 18736 13654
rect 18800 13462 18828 14826
rect 18892 14550 18920 15302
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18878 13968 18934 13977
rect 18878 13903 18934 13912
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18512 13320 18564 13326
rect 18510 13288 18512 13297
rect 18696 13320 18748 13326
rect 18564 13288 18566 13297
rect 18696 13262 18748 13268
rect 18510 13223 18566 13232
rect 18892 13190 18920 13903
rect 18880 13184 18932 13190
rect 18786 13152 18842 13161
rect 18880 13126 18932 13132
rect 18786 13087 18842 13096
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18524 12434 18552 12786
rect 18800 12782 18828 13087
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18432 12406 18552 12434
rect 18878 12472 18934 12481
rect 18878 12407 18934 12416
rect 18432 12238 18460 12406
rect 18892 12374 18920 12407
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18984 12306 19012 15422
rect 19260 14550 19288 16526
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 13734 19196 14214
rect 19156 13728 19208 13734
rect 19352 13682 19380 16458
rect 19444 15638 19472 17190
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 14657 19472 15302
rect 19536 15194 19564 17478
rect 19614 16280 19670 16289
rect 19614 16215 19670 16224
rect 19628 15881 19656 16215
rect 19614 15872 19670 15881
rect 19614 15807 19670 15816
rect 19720 15434 19748 17478
rect 19798 16960 19854 16969
rect 19996 16946 20024 18294
rect 20088 17592 20116 18414
rect 20364 18086 20392 18770
rect 20352 18080 20404 18086
rect 20456 18068 20484 18822
rect 20536 18692 20588 18698
rect 21008 18680 21036 20810
rect 21192 19334 21220 21898
rect 21284 20534 21312 22066
rect 21468 22098 21496 22986
rect 21560 22710 21588 23462
rect 21652 23118 21680 24840
rect 21744 24410 21772 24942
rect 21836 24854 21864 25871
rect 21928 25702 21956 26182
rect 21916 25696 21968 25702
rect 21916 25638 21968 25644
rect 22020 25430 22048 26302
rect 22008 25424 22060 25430
rect 21914 25392 21970 25401
rect 22008 25366 22060 25372
rect 21914 25327 21970 25336
rect 21928 25276 21956 25327
rect 21928 25248 22048 25276
rect 22020 25158 22048 25248
rect 22008 25152 22060 25158
rect 21914 25120 21970 25129
rect 22008 25094 22060 25100
rect 22112 25106 22140 26404
rect 22244 26404 22324 26432
rect 22374 26415 22430 26424
rect 22192 26386 22244 26392
rect 22190 26208 22246 26217
rect 22190 26143 22246 26152
rect 22204 25906 22232 26143
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 22204 25401 22232 25638
rect 22296 25514 22324 26404
rect 22376 26240 22428 26246
rect 22376 26182 22428 26188
rect 22388 26081 22416 26182
rect 22374 26072 22430 26081
rect 22374 26007 22430 26016
rect 22480 25945 22508 27084
rect 22572 26994 22600 27775
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22572 26450 22600 26726
rect 22560 26444 22612 26450
rect 22560 26386 22612 26392
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22572 26081 22600 26250
rect 22558 26072 22614 26081
rect 22558 26007 22614 26016
rect 22466 25936 22522 25945
rect 22466 25871 22522 25880
rect 22664 25888 22692 28966
rect 22756 28490 22784 28999
rect 22744 28484 22796 28490
rect 22744 28426 22796 28432
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 22756 27538 22784 28018
rect 22848 27577 22876 29446
rect 23216 29345 23244 29804
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23308 29481 23336 29582
rect 23294 29472 23350 29481
rect 23294 29407 23350 29416
rect 23018 29336 23074 29345
rect 23018 29271 23074 29280
rect 23202 29336 23258 29345
rect 23202 29271 23258 29280
rect 23032 29152 23060 29271
rect 23216 29152 23244 29271
rect 23296 29164 23348 29170
rect 23032 29124 23079 29152
rect 23216 29124 23296 29152
rect 23051 29084 23079 29124
rect 23296 29106 23348 29112
rect 23051 29073 23152 29084
rect 22926 29064 22982 29073
rect 23051 29064 23166 29073
rect 23051 29056 23110 29064
rect 22982 29008 23060 29016
rect 22926 28999 23060 29008
rect 23110 28999 23166 29008
rect 23294 29064 23350 29073
rect 23294 28999 23296 29008
rect 22940 28988 23060 28999
rect 22928 28688 22980 28694
rect 22928 28630 22980 28636
rect 23032 28642 23060 28988
rect 23348 28999 23350 29008
rect 23296 28970 23348 28976
rect 23110 28928 23166 28937
rect 23400 28914 23428 30738
rect 23110 28863 23166 28872
rect 23296 28886 23428 28914
rect 23124 28762 23152 28863
rect 23112 28756 23164 28762
rect 23112 28698 23164 28704
rect 23204 28756 23256 28762
rect 23204 28698 23256 28704
rect 23216 28642 23244 28698
rect 23296 28676 23324 28886
rect 23492 28762 23520 31583
rect 23584 31346 23612 32166
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23676 31278 23704 32286
rect 23754 32192 23810 32201
rect 23754 32127 23810 32136
rect 23768 31482 23796 32127
rect 23860 32026 23888 32370
rect 24412 32150 24808 32178
rect 23848 32020 23900 32026
rect 23848 31962 23900 31968
rect 24412 31890 24440 32150
rect 24492 32020 24544 32026
rect 24492 31962 24544 31968
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 23848 31680 23900 31686
rect 23846 31648 23848 31657
rect 23900 31648 23902 31657
rect 23846 31583 23902 31592
rect 23996 31580 24304 31589
rect 23996 31578 24002 31580
rect 24058 31578 24082 31580
rect 24138 31578 24162 31580
rect 24218 31578 24242 31580
rect 24298 31578 24304 31580
rect 24058 31526 24060 31578
rect 24240 31526 24242 31578
rect 23996 31524 24002 31526
rect 24058 31524 24082 31526
rect 24138 31524 24162 31526
rect 24218 31524 24242 31526
rect 24298 31524 24304 31526
rect 23846 31512 23902 31521
rect 23996 31515 24304 31524
rect 23756 31476 23808 31482
rect 23846 31447 23848 31456
rect 23756 31418 23808 31424
rect 23900 31447 23902 31456
rect 23848 31418 23900 31424
rect 23768 31346 23796 31418
rect 23756 31340 23808 31346
rect 23756 31282 23808 31288
rect 23664 31272 23716 31278
rect 23664 31214 23716 31220
rect 23848 31272 23900 31278
rect 23848 31214 23900 31220
rect 23860 31142 23888 31214
rect 23756 31136 23808 31142
rect 23756 31078 23808 31084
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 24308 31136 24360 31142
rect 24308 31078 24360 31084
rect 23662 30832 23718 30841
rect 23662 30767 23718 30776
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23584 30122 23612 30670
rect 23572 30116 23624 30122
rect 23572 30058 23624 30064
rect 23584 29714 23612 30058
rect 23572 29708 23624 29714
rect 23572 29650 23624 29656
rect 23676 29646 23704 30767
rect 23768 30569 23796 31078
rect 23848 30592 23900 30598
rect 23754 30560 23810 30569
rect 24320 30580 24348 31078
rect 24412 30648 24440 31826
rect 24504 31657 24532 31962
rect 24780 31958 24808 32150
rect 24584 31952 24636 31958
rect 24584 31894 24636 31900
rect 24768 31952 24820 31958
rect 24768 31894 24820 31900
rect 24490 31648 24546 31657
rect 24490 31583 24546 31592
rect 24490 31512 24546 31521
rect 24596 31482 24624 31894
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 24490 31447 24492 31456
rect 24544 31447 24546 31456
rect 24584 31476 24636 31482
rect 24492 31418 24544 31424
rect 24584 31418 24636 31424
rect 24504 31346 24532 31418
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24596 30938 24624 31078
rect 24584 30932 24636 30938
rect 24688 30920 24716 31758
rect 24780 31142 24808 31758
rect 24872 31142 24900 32438
rect 24964 31657 24992 34439
rect 25134 33280 25190 33289
rect 25134 33215 25190 33224
rect 25148 32502 25176 33215
rect 25228 32836 25280 32842
rect 25228 32778 25280 32784
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 24950 31648 25006 31657
rect 24950 31583 25006 31592
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24860 31136 24912 31142
rect 24860 31078 24912 31084
rect 24768 30932 24820 30938
rect 24688 30892 24768 30920
rect 24584 30874 24636 30880
rect 24768 30874 24820 30880
rect 24492 30660 24544 30666
rect 24412 30620 24492 30648
rect 24492 30602 24544 30608
rect 24596 30648 24624 30874
rect 24780 30841 24808 30874
rect 24766 30832 24822 30841
rect 24766 30767 24822 30776
rect 24676 30660 24728 30666
rect 24596 30620 24676 30648
rect 24320 30552 24440 30580
rect 23848 30534 23900 30540
rect 23754 30495 23810 30504
rect 23754 30424 23810 30433
rect 23754 30359 23810 30368
rect 23768 30282 23796 30359
rect 23756 30276 23808 30282
rect 23756 30218 23808 30224
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 23768 29714 23796 30126
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23572 29572 23624 29578
rect 23572 29514 23624 29520
rect 23584 29034 23612 29514
rect 23676 29345 23704 29582
rect 23754 29472 23810 29481
rect 23754 29407 23810 29416
rect 23662 29336 23718 29345
rect 23662 29271 23718 29280
rect 23662 29200 23718 29209
rect 23662 29135 23664 29144
rect 23716 29135 23718 29144
rect 23664 29106 23716 29112
rect 23572 29028 23624 29034
rect 23572 28970 23624 28976
rect 23664 29028 23716 29034
rect 23664 28970 23716 28976
rect 23570 28928 23626 28937
rect 23570 28863 23626 28872
rect 23388 28756 23440 28762
rect 23388 28698 23440 28704
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 23296 28648 23336 28676
rect 22940 28540 22968 28630
rect 23032 28614 23244 28642
rect 22940 28512 23152 28540
rect 23039 28416 23091 28422
rect 23124 28404 23152 28512
rect 23124 28376 23244 28404
rect 23039 28358 23091 28364
rect 23051 28234 23079 28358
rect 23051 28206 23152 28234
rect 22926 28112 22982 28121
rect 22926 28047 22982 28056
rect 23020 28076 23072 28082
rect 22834 27568 22890 27577
rect 22744 27532 22796 27538
rect 22834 27503 22890 27512
rect 22744 27474 22796 27480
rect 22940 27441 22968 28047
rect 23020 28018 23072 28024
rect 23032 27577 23060 28018
rect 23018 27568 23074 27577
rect 23018 27503 23074 27512
rect 22926 27432 22982 27441
rect 22836 27396 22888 27402
rect 22926 27367 22982 27376
rect 22836 27338 22888 27344
rect 22742 27296 22798 27305
rect 22742 27231 22798 27240
rect 22756 26246 22784 27231
rect 22744 26240 22796 26246
rect 22744 26182 22796 26188
rect 22756 26042 22784 26182
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22848 25956 22876 27338
rect 22928 27328 22980 27334
rect 23032 27305 23060 27503
rect 22928 27270 22980 27276
rect 23018 27296 23074 27305
rect 22940 27130 22968 27270
rect 23018 27231 23074 27240
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22926 27024 22982 27033
rect 22926 26959 22928 26968
rect 22980 26959 22982 26968
rect 22928 26930 22980 26936
rect 23020 26852 23072 26858
rect 23020 26794 23072 26800
rect 23032 26364 23060 26794
rect 23124 26518 23152 28206
rect 23216 28082 23244 28376
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23308 27606 23336 28648
rect 23400 28098 23428 28698
rect 23584 28694 23612 28863
rect 23572 28688 23624 28694
rect 23572 28630 23624 28636
rect 23676 28506 23704 28970
rect 23768 28762 23796 29407
rect 23756 28756 23808 28762
rect 23756 28698 23808 28704
rect 23492 28478 23704 28506
rect 23492 28218 23520 28478
rect 23572 28416 23624 28422
rect 23570 28384 23572 28393
rect 23756 28416 23808 28422
rect 23624 28384 23626 28393
rect 23756 28358 23808 28364
rect 23570 28319 23626 28328
rect 23480 28212 23532 28218
rect 23480 28154 23532 28160
rect 23584 28150 23612 28319
rect 23662 28248 23718 28257
rect 23662 28183 23664 28192
rect 23716 28183 23718 28192
rect 23664 28154 23716 28160
rect 23572 28144 23624 28150
rect 23400 28070 23520 28098
rect 23572 28086 23624 28092
rect 23296 27600 23348 27606
rect 23202 27568 23258 27577
rect 23296 27542 23348 27548
rect 23386 27568 23442 27577
rect 23202 27503 23258 27512
rect 23386 27503 23442 27512
rect 23216 27470 23244 27503
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23294 27432 23350 27441
rect 23216 26994 23244 27406
rect 23294 27367 23350 27376
rect 23308 27010 23336 27367
rect 23400 27130 23428 27503
rect 23492 27130 23520 28070
rect 23570 27976 23626 27985
rect 23570 27911 23626 27920
rect 23584 27674 23612 27911
rect 23572 27668 23624 27674
rect 23572 27610 23624 27616
rect 23768 27441 23796 28358
rect 23754 27432 23810 27441
rect 23754 27367 23810 27376
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23662 27296 23718 27305
rect 23376 27124 23428 27130
rect 23376 27066 23428 27072
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23204 26988 23256 26994
rect 23308 26982 23428 27010
rect 23204 26930 23256 26936
rect 23400 26926 23428 26982
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23204 26852 23256 26858
rect 23204 26794 23256 26800
rect 23112 26512 23164 26518
rect 23112 26454 23164 26460
rect 23032 26336 23152 26364
rect 22848 25928 23060 25956
rect 22664 25860 22876 25888
rect 22560 25832 22612 25838
rect 22612 25792 22784 25820
rect 22560 25774 22612 25780
rect 22376 25764 22428 25770
rect 22428 25724 22508 25752
rect 22376 25706 22428 25712
rect 22480 25684 22508 25724
rect 22480 25656 22600 25684
rect 22296 25486 22416 25514
rect 22388 25480 22416 25486
rect 22388 25452 22508 25480
rect 22284 25424 22336 25430
rect 22190 25392 22246 25401
rect 22336 25384 22416 25412
rect 22284 25366 22336 25372
rect 22190 25327 22246 25336
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22112 25078 22232 25106
rect 21914 25055 21970 25064
rect 21928 24954 21956 25055
rect 22006 24984 22062 24993
rect 21916 24948 21968 24954
rect 22062 24942 22140 24970
rect 22006 24919 22062 24928
rect 21916 24890 21968 24896
rect 21836 24826 21956 24854
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21836 24614 21864 24686
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21732 23792 21784 23798
rect 21732 23734 21784 23740
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21548 22704 21600 22710
rect 21548 22646 21600 22652
rect 21638 22672 21694 22681
rect 21638 22607 21694 22616
rect 21652 22574 21680 22607
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21362 22063 21418 22072
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21376 21690 21404 21966
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 21376 20380 21404 21626
rect 21468 21146 21496 22034
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21560 21010 21588 22510
rect 21638 21856 21694 21865
rect 21638 21791 21694 21800
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21652 20913 21680 21791
rect 21638 20904 21694 20913
rect 21638 20839 21694 20848
rect 21638 20632 21694 20641
rect 21638 20567 21694 20576
rect 21652 20466 21680 20567
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21456 20392 21508 20398
rect 21376 20352 21456 20380
rect 21456 20334 21508 20340
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 20588 18652 21036 18680
rect 21100 19306 21220 19334
rect 20536 18634 20588 18640
rect 21100 18601 21128 19306
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21086 18592 21142 18601
rect 21086 18527 21142 18536
rect 21088 18148 21140 18154
rect 21088 18090 21140 18096
rect 20456 18040 20576 18068
rect 20352 18022 20404 18028
rect 20155 17980 20463 17989
rect 20155 17978 20161 17980
rect 20217 17978 20241 17980
rect 20297 17978 20321 17980
rect 20377 17978 20401 17980
rect 20457 17978 20463 17980
rect 20217 17926 20219 17978
rect 20399 17926 20401 17978
rect 20155 17924 20161 17926
rect 20217 17924 20241 17926
rect 20297 17924 20321 17926
rect 20377 17924 20401 17926
rect 20457 17924 20463 17926
rect 20155 17915 20463 17924
rect 20168 17604 20220 17610
rect 20088 17564 20168 17592
rect 20168 17546 20220 17552
rect 20548 16980 20576 18040
rect 21100 17814 21128 18090
rect 21088 17808 21140 17814
rect 20732 17734 20944 17762
rect 21088 17750 21140 17756
rect 20732 17678 20760 17734
rect 20720 17672 20772 17678
rect 20626 17640 20682 17649
rect 20720 17614 20772 17620
rect 20626 17575 20682 17584
rect 20640 17542 20668 17575
rect 20732 17542 20760 17614
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20824 17270 20852 17546
rect 20628 17264 20680 17270
rect 20628 17206 20680 17212
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 19798 16895 19854 16904
rect 19904 16918 20024 16946
rect 20088 16952 20576 16980
rect 19812 16794 19840 16895
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19904 16708 19932 16918
rect 19982 16824 20038 16833
rect 20088 16810 20116 16952
rect 20155 16892 20463 16901
rect 20155 16890 20161 16892
rect 20217 16890 20241 16892
rect 20297 16890 20321 16892
rect 20377 16890 20401 16892
rect 20457 16890 20463 16892
rect 20217 16838 20219 16890
rect 20399 16838 20401 16890
rect 20155 16836 20161 16838
rect 20217 16836 20241 16838
rect 20297 16836 20321 16838
rect 20377 16836 20401 16838
rect 20457 16836 20463 16838
rect 20155 16827 20463 16836
rect 20038 16782 20116 16810
rect 19982 16759 20038 16768
rect 19904 16680 20024 16708
rect 19800 16516 19852 16522
rect 19852 16476 19932 16504
rect 19800 16458 19852 16464
rect 19904 15745 19932 16476
rect 19890 15736 19946 15745
rect 19890 15671 19946 15680
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19628 15314 19656 15370
rect 19628 15286 19840 15314
rect 19536 15166 19656 15194
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19430 14648 19486 14657
rect 19430 14583 19486 14592
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19156 13670 19208 13676
rect 19260 13654 19380 13682
rect 19154 13560 19210 13569
rect 19260 13530 19288 13654
rect 19154 13495 19210 13504
rect 19248 13524 19300 13530
rect 19062 13288 19118 13297
rect 19062 13223 19118 13232
rect 19076 12646 19104 13223
rect 19168 13002 19196 13495
rect 19248 13466 19300 13472
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19352 13433 19380 13466
rect 19338 13424 19394 13433
rect 19338 13359 19394 13368
rect 19168 12974 19288 13002
rect 19260 12918 19288 12974
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18248 11762 18276 12038
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18340 11762 18368 11834
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 19168 11014 19196 12854
rect 19260 11218 19288 12854
rect 19444 12730 19472 13942
rect 19352 12702 19472 12730
rect 19536 12714 19564 14894
rect 19628 14482 19656 15166
rect 19812 15094 19840 15286
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19720 14657 19748 14758
rect 19706 14648 19762 14657
rect 19706 14583 19762 14592
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19720 14414 19748 14583
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19614 14104 19670 14113
rect 19614 14039 19670 14048
rect 19628 14006 19656 14039
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19616 13456 19668 13462
rect 19616 13398 19668 13404
rect 19628 13190 19656 13398
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19524 12708 19576 12714
rect 19352 12646 19380 12702
rect 19524 12650 19576 12656
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19522 12064 19578 12073
rect 19522 11999 19578 12008
rect 19536 11898 19564 11999
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 17684 10464 17736 10470
rect 15750 10432 15806 10441
rect 19720 10441 19748 14214
rect 19890 14104 19946 14113
rect 19890 14039 19946 14048
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19812 13161 19840 13262
rect 19798 13152 19854 13161
rect 19798 13087 19854 13096
rect 19904 12617 19932 14039
rect 19996 13705 20024 16680
rect 20534 16688 20590 16697
rect 20534 16623 20590 16632
rect 20548 16250 20576 16623
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20640 16182 20668 17206
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20272 15910 20300 15982
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20155 15804 20463 15813
rect 20155 15802 20161 15804
rect 20217 15802 20241 15804
rect 20297 15802 20321 15804
rect 20377 15802 20401 15804
rect 20457 15802 20463 15804
rect 20217 15750 20219 15802
rect 20399 15750 20401 15802
rect 20155 15748 20161 15750
rect 20217 15748 20241 15750
rect 20297 15748 20321 15750
rect 20377 15748 20401 15750
rect 20457 15748 20463 15750
rect 20155 15739 20463 15748
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20088 14822 20116 15506
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 15201 20760 15370
rect 20718 15192 20774 15201
rect 20718 15127 20774 15136
rect 20824 15065 20852 17002
rect 20916 15706 20944 17734
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20810 15056 20866 15065
rect 20810 14991 20866 15000
rect 21008 14929 21036 17614
rect 21100 17202 21128 17750
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21192 17066 21220 19178
rect 21284 19174 21312 19450
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21272 18692 21324 18698
rect 21272 18634 21324 18640
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 21178 16552 21234 16561
rect 21178 16487 21234 16496
rect 21192 16114 21220 16487
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21086 15736 21142 15745
rect 21086 15671 21142 15680
rect 20994 14920 21050 14929
rect 20812 14884 20864 14890
rect 20994 14855 21050 14864
rect 20812 14826 20864 14832
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20155 14716 20463 14725
rect 20155 14714 20161 14716
rect 20217 14714 20241 14716
rect 20297 14714 20321 14716
rect 20377 14714 20401 14716
rect 20457 14714 20463 14716
rect 20217 14662 20219 14714
rect 20399 14662 20401 14714
rect 20155 14660 20161 14662
rect 20217 14660 20241 14662
rect 20297 14660 20321 14662
rect 20377 14660 20401 14662
rect 20457 14660 20463 14662
rect 20155 14651 20463 14660
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20350 14512 20406 14521
rect 20350 14447 20406 14456
rect 20364 14278 20392 14447
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20456 13870 20484 14554
rect 20534 14376 20590 14385
rect 20534 14311 20590 14320
rect 20548 14006 20576 14311
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20444 13864 20496 13870
rect 20088 13824 20444 13852
rect 19982 13696 20038 13705
rect 19982 13631 20038 13640
rect 19984 12640 20036 12646
rect 19890 12608 19946 12617
rect 19984 12582 20036 12588
rect 19890 12543 19946 12552
rect 19904 12442 19932 12543
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19996 12238 20024 12582
rect 20088 12238 20116 13824
rect 20444 13806 20496 13812
rect 20824 13802 20852 14826
rect 21100 14278 21128 15671
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21192 14278 21220 14554
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 20812 13796 20864 13802
rect 20640 13756 20812 13784
rect 20155 13628 20463 13637
rect 20155 13626 20161 13628
rect 20217 13626 20241 13628
rect 20297 13626 20321 13628
rect 20377 13626 20401 13628
rect 20457 13626 20463 13628
rect 20217 13574 20219 13626
rect 20399 13574 20401 13626
rect 20155 13572 20161 13574
rect 20217 13572 20241 13574
rect 20297 13572 20321 13574
rect 20377 13572 20401 13574
rect 20457 13572 20463 13574
rect 20155 13563 20463 13572
rect 20534 13152 20590 13161
rect 20534 13087 20590 13096
rect 20155 12540 20463 12549
rect 20155 12538 20161 12540
rect 20217 12538 20241 12540
rect 20297 12538 20321 12540
rect 20377 12538 20401 12540
rect 20457 12538 20463 12540
rect 20217 12486 20219 12538
rect 20399 12486 20401 12538
rect 20155 12484 20161 12486
rect 20217 12484 20241 12486
rect 20297 12484 20321 12486
rect 20377 12484 20401 12486
rect 20457 12484 20463 12486
rect 20155 12475 20463 12484
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19982 12064 20038 12073
rect 19904 11694 19932 12038
rect 19982 11999 20038 12008
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19904 11150 19932 11630
rect 19996 11529 20024 11999
rect 19982 11520 20038 11529
rect 19982 11455 20038 11464
rect 20155 11452 20463 11461
rect 20155 11450 20161 11452
rect 20217 11450 20241 11452
rect 20297 11450 20321 11452
rect 20377 11450 20401 11452
rect 20457 11450 20463 11452
rect 20217 11398 20219 11450
rect 20399 11398 20401 11450
rect 20155 11396 20161 11398
rect 20217 11396 20241 11398
rect 20297 11396 20321 11398
rect 20377 11396 20401 11398
rect 20457 11396 20463 11398
rect 20155 11387 20463 11396
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 10810 19932 11086
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 20088 10674 20116 10950
rect 20548 10810 20576 13087
rect 20640 12782 20668 13756
rect 20812 13738 20864 13744
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20810 13288 20866 13297
rect 21008 13258 21036 13738
rect 20810 13223 20866 13232
rect 20996 13252 21048 13258
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 12434 20760 12718
rect 20640 12406 20760 12434
rect 20640 12238 20668 12406
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20732 11558 20760 11630
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20824 11150 20852 13223
rect 20996 13194 21048 13200
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20916 11218 20944 11698
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20916 11082 20944 11154
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20902 10840 20958 10849
rect 20536 10804 20588 10810
rect 20902 10775 20904 10784
rect 20536 10746 20588 10752
rect 20956 10775 20958 10784
rect 20904 10746 20956 10752
rect 20902 10704 20958 10713
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20720 10668 20772 10674
rect 20772 10628 20852 10656
rect 20902 10639 20904 10648
rect 20720 10610 20772 10616
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 17684 10406 17736 10412
rect 19706 10432 19762 10441
rect 15750 10367 15806 10376
rect 19706 10367 19762 10376
rect 20155 10364 20463 10373
rect 20155 10362 20161 10364
rect 20217 10362 20241 10364
rect 20297 10362 20321 10364
rect 20377 10362 20401 10364
rect 20457 10362 20463 10364
rect 20217 10310 20219 10362
rect 20399 10310 20401 10362
rect 20155 10308 20161 10310
rect 20217 10308 20241 10310
rect 20297 10308 20321 10310
rect 20377 10308 20401 10310
rect 20457 10308 20463 10310
rect 20155 10299 20463 10308
rect 20732 10266 20760 10474
rect 20824 10470 20852 10628
rect 20956 10639 20958 10648
rect 20904 10610 20956 10616
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20916 10305 20944 10610
rect 20902 10296 20958 10305
rect 20720 10260 20772 10266
rect 21008 10266 21036 12854
rect 21100 11676 21128 14214
rect 21284 11762 21312 18634
rect 21376 16590 21404 19654
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21468 19156 21496 19246
rect 21560 19224 21588 20198
rect 21652 20058 21680 20266
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21560 19196 21680 19224
rect 21468 19128 21588 19156
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21468 17785 21496 18362
rect 21454 17776 21510 17785
rect 21454 17711 21510 17720
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16794 21496 16934
rect 21560 16794 21588 19128
rect 21652 18850 21680 19196
rect 21744 19174 21772 23734
rect 21836 23225 21864 24278
rect 21928 23594 21956 24826
rect 22006 24848 22062 24857
rect 22112 24818 22140 24942
rect 22204 24857 22232 25078
rect 22296 24954 22324 25230
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22190 24848 22246 24857
rect 22006 24783 22062 24792
rect 22100 24812 22152 24818
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 22020 23304 22048 24783
rect 22190 24783 22246 24792
rect 22100 24754 22152 24760
rect 22296 24562 22324 24890
rect 22112 24534 22324 24562
rect 22112 24206 22140 24534
rect 22388 24449 22416 25384
rect 22480 24854 22508 25452
rect 22572 25265 22600 25656
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22558 25256 22614 25265
rect 22664 25226 22692 25298
rect 22558 25191 22614 25200
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22480 24826 22600 24854
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22190 24440 22246 24449
rect 22190 24375 22246 24384
rect 22374 24440 22430 24449
rect 22374 24375 22430 24384
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22098 23760 22154 23769
rect 22204 23730 22232 24375
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22098 23695 22154 23704
rect 22192 23724 22244 23730
rect 21928 23276 22048 23304
rect 21822 23216 21878 23225
rect 21822 23151 21878 23160
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21836 22506 21864 23054
rect 21928 22642 21956 23276
rect 22006 23216 22062 23225
rect 22112 23186 22140 23695
rect 22192 23666 22244 23672
rect 22006 23151 22062 23160
rect 22100 23180 22152 23186
rect 22020 22953 22048 23151
rect 22100 23122 22152 23128
rect 22192 23112 22244 23118
rect 22296 23100 22324 24210
rect 22480 24177 22508 24550
rect 22466 24168 22522 24177
rect 22466 24103 22522 24112
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22388 23526 22416 23802
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22244 23072 22324 23100
rect 22192 23054 22244 23060
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 22006 22944 22062 22953
rect 22006 22879 22062 22888
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21824 22500 21876 22506
rect 21824 22442 21876 22448
rect 21836 21418 21864 22442
rect 21928 22166 21956 22578
rect 21916 22160 21968 22166
rect 22020 22137 22048 22714
rect 21916 22102 21968 22108
rect 22006 22128 22062 22137
rect 22006 22063 22062 22072
rect 22112 21894 22140 22986
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22204 21729 22232 22374
rect 22190 21720 22246 21729
rect 22296 21690 22324 23072
rect 22374 22944 22430 22953
rect 22374 22879 22430 22888
rect 22388 22574 22416 22879
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22480 22438 22508 23666
rect 22572 23254 22600 24826
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22664 24041 22692 24550
rect 22650 24032 22706 24041
rect 22650 23967 22706 23976
rect 22664 23594 22692 23967
rect 22756 23905 22784 25792
rect 22848 24256 22876 25860
rect 23032 24834 23060 25928
rect 23124 25906 23152 26336
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23216 25480 23244 26794
rect 23308 25786 23336 26862
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23400 26450 23428 26726
rect 23492 26518 23520 26930
rect 23584 26858 23612 27270
rect 23662 27231 23718 27240
rect 23669 27062 23697 27231
rect 23664 27056 23716 27062
rect 23664 26998 23716 27004
rect 23754 27024 23810 27033
rect 23754 26959 23810 26968
rect 23572 26852 23624 26858
rect 23572 26794 23624 26800
rect 23768 26738 23796 26959
rect 23860 26926 23888 30534
rect 23996 30492 24304 30501
rect 23996 30490 24002 30492
rect 24058 30490 24082 30492
rect 24138 30490 24162 30492
rect 24218 30490 24242 30492
rect 24298 30490 24304 30492
rect 24058 30438 24060 30490
rect 24240 30438 24242 30490
rect 23996 30436 24002 30438
rect 24058 30436 24082 30438
rect 24138 30436 24162 30438
rect 24218 30436 24242 30438
rect 24298 30436 24304 30438
rect 23996 30427 24304 30436
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24124 30116 24176 30122
rect 24124 30058 24176 30064
rect 23938 30016 23994 30025
rect 23938 29951 23994 29960
rect 23952 29782 23980 29951
rect 24136 29850 24164 30058
rect 24228 29850 24256 30262
rect 24124 29844 24176 29850
rect 24124 29786 24176 29792
rect 24216 29844 24268 29850
rect 24216 29786 24268 29792
rect 23940 29776 23992 29782
rect 23940 29718 23992 29724
rect 24228 29510 24256 29786
rect 24216 29504 24268 29510
rect 24216 29446 24268 29452
rect 23996 29404 24304 29413
rect 23996 29402 24002 29404
rect 24058 29402 24082 29404
rect 24138 29402 24162 29404
rect 24218 29402 24242 29404
rect 24298 29402 24304 29404
rect 24058 29350 24060 29402
rect 24240 29350 24242 29402
rect 23996 29348 24002 29350
rect 24058 29348 24082 29350
rect 24138 29348 24162 29350
rect 24218 29348 24242 29350
rect 24298 29348 24304 29350
rect 23996 29339 24304 29348
rect 24214 29200 24270 29209
rect 24032 29164 24084 29170
rect 24214 29135 24270 29144
rect 24308 29164 24360 29170
rect 24032 29106 24084 29112
rect 24044 29034 24072 29106
rect 24032 29028 24084 29034
rect 24032 28970 24084 28976
rect 23938 28928 23994 28937
rect 23938 28863 23994 28872
rect 23952 28490 23980 28863
rect 24228 28626 24256 29135
rect 24308 29106 24360 29112
rect 24320 29073 24348 29106
rect 24412 29102 24440 30552
rect 24490 30424 24546 30433
rect 24490 30359 24546 30368
rect 24400 29096 24452 29102
rect 24306 29064 24362 29073
rect 24400 29038 24452 29044
rect 24306 28999 24308 29008
rect 24360 28999 24362 29008
rect 24308 28970 24360 28976
rect 24320 28939 24348 28970
rect 24400 28960 24452 28966
rect 24400 28902 24452 28908
rect 24124 28620 24176 28626
rect 24124 28562 24176 28568
rect 24216 28620 24268 28626
rect 24216 28562 24268 28568
rect 24136 28490 24164 28562
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 24124 28484 24176 28490
rect 24124 28426 24176 28432
rect 23996 28316 24304 28325
rect 23996 28314 24002 28316
rect 24058 28314 24082 28316
rect 24138 28314 24162 28316
rect 24218 28314 24242 28316
rect 24298 28314 24304 28316
rect 24058 28262 24060 28314
rect 24240 28262 24242 28314
rect 23996 28260 24002 28262
rect 24058 28260 24082 28262
rect 24138 28260 24162 28262
rect 24218 28260 24242 28262
rect 24298 28260 24304 28262
rect 23996 28251 24304 28260
rect 24216 28212 24268 28218
rect 24268 28172 24348 28200
rect 24216 28154 24268 28160
rect 23940 28144 23992 28150
rect 23940 28086 23992 28092
rect 23952 27402 23980 28086
rect 24124 28076 24176 28082
rect 24124 28018 24176 28024
rect 24136 27849 24164 28018
rect 24320 27985 24348 28172
rect 24412 28150 24440 28902
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24400 28008 24452 28014
rect 24306 27976 24362 27985
rect 24216 27940 24268 27946
rect 24400 27950 24452 27956
rect 24306 27911 24362 27920
rect 24216 27882 24268 27888
rect 24122 27840 24178 27849
rect 24122 27775 24178 27784
rect 24030 27568 24086 27577
rect 24030 27503 24086 27512
rect 23940 27396 23992 27402
rect 23940 27338 23992 27344
rect 24044 27334 24072 27503
rect 24136 27441 24164 27775
rect 24228 27470 24256 27882
rect 24216 27464 24268 27470
rect 24122 27432 24178 27441
rect 24216 27406 24268 27412
rect 24122 27367 24178 27376
rect 24032 27328 24084 27334
rect 24032 27270 24084 27276
rect 23996 27228 24304 27237
rect 23996 27226 24002 27228
rect 24058 27226 24082 27228
rect 24138 27226 24162 27228
rect 24218 27226 24242 27228
rect 24298 27226 24304 27228
rect 24058 27174 24060 27226
rect 24240 27174 24242 27226
rect 23996 27172 24002 27174
rect 24058 27172 24082 27174
rect 24138 27172 24162 27174
rect 24218 27172 24242 27174
rect 24298 27172 24304 27174
rect 23996 27163 24304 27172
rect 24032 27124 24084 27130
rect 24032 27066 24084 27072
rect 23940 27056 23992 27062
rect 24044 27033 24072 27066
rect 23940 26998 23992 27004
rect 24030 27024 24086 27033
rect 23848 26920 23900 26926
rect 23848 26862 23900 26868
rect 23584 26710 23796 26738
rect 23480 26512 23532 26518
rect 23480 26454 23532 26460
rect 23584 26466 23612 26710
rect 23662 26616 23718 26625
rect 23846 26616 23902 26625
rect 23718 26574 23796 26602
rect 23662 26551 23718 26560
rect 23388 26444 23440 26450
rect 23584 26438 23704 26466
rect 23388 26386 23440 26392
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 23308 25758 23440 25786
rect 23412 25514 23440 25758
rect 23124 25452 23244 25480
rect 23308 25486 23440 25514
rect 23124 25362 23152 25452
rect 23112 25356 23164 25362
rect 23112 25298 23164 25304
rect 23204 25356 23256 25362
rect 23204 25298 23256 25304
rect 23216 25158 23244 25298
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23032 24806 23244 24834
rect 23020 24744 23072 24750
rect 23020 24686 23072 24692
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 22940 24410 22968 24618
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 22928 24268 22980 24274
rect 22848 24228 22928 24256
rect 22928 24210 22980 24216
rect 22926 24168 22982 24177
rect 22836 24132 22888 24138
rect 22926 24103 22982 24112
rect 22836 24074 22888 24080
rect 22848 24041 22876 24074
rect 22834 24032 22890 24041
rect 22834 23967 22890 23976
rect 22742 23896 22798 23905
rect 22742 23831 22798 23840
rect 22940 23798 22968 24103
rect 22928 23792 22980 23798
rect 22742 23760 22798 23769
rect 22928 23734 22980 23740
rect 22742 23695 22798 23704
rect 22756 23662 22784 23695
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 22744 23520 22796 23526
rect 23032 23474 23060 24686
rect 23124 23526 23152 24686
rect 23216 23905 23244 24806
rect 23202 23896 23258 23905
rect 23202 23831 23258 23840
rect 23204 23588 23256 23594
rect 23204 23530 23256 23536
rect 22744 23462 22796 23468
rect 22560 23248 22612 23254
rect 22560 23190 22612 23196
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22572 22250 22600 23190
rect 22756 22778 22784 23462
rect 22848 23446 23060 23474
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22742 22672 22798 22681
rect 22652 22636 22704 22642
rect 22848 22658 22876 23446
rect 23124 23186 23152 23462
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 22798 22630 22876 22658
rect 22742 22607 22798 22616
rect 22652 22578 22704 22584
rect 22480 22222 22600 22250
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22190 21655 22246 21664
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21822 21312 21878 21321
rect 21822 21247 21878 21256
rect 21732 19168 21784 19174
rect 21836 19156 21864 21247
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21928 20210 21956 20402
rect 22006 20360 22062 20369
rect 22112 20346 22140 21490
rect 22190 21176 22246 21185
rect 22388 21162 22416 21898
rect 22480 21418 22508 22222
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22246 21134 22416 21162
rect 22190 21111 22246 21120
rect 22466 20768 22522 20777
rect 22466 20703 22522 20712
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22282 20496 22338 20505
rect 22282 20431 22338 20440
rect 22296 20398 22324 20431
rect 22388 20398 22416 20538
rect 22062 20318 22140 20346
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22006 20295 22062 20304
rect 22374 20224 22430 20233
rect 21928 20182 22374 20210
rect 22374 20159 22430 20168
rect 22480 19990 22508 20703
rect 21916 19984 21968 19990
rect 22468 19984 22520 19990
rect 21916 19926 21968 19932
rect 22006 19952 22062 19961
rect 21928 19224 21956 19926
rect 22062 19910 22324 19938
rect 22468 19926 22520 19932
rect 22006 19887 22062 19896
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22112 19689 22140 19722
rect 22098 19680 22154 19689
rect 22098 19615 22154 19624
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 21928 19196 22048 19224
rect 21836 19128 21956 19156
rect 21732 19110 21784 19116
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21652 18822 21772 18850
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21652 18222 21680 18702
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21744 18057 21772 18822
rect 21836 18630 21864 18906
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 21836 18086 21864 18294
rect 21824 18080 21876 18086
rect 21730 18048 21786 18057
rect 21824 18022 21876 18028
rect 21730 17983 21786 17992
rect 21744 17270 21772 17983
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21376 14482 21404 16390
rect 21468 15706 21496 16458
rect 21560 16046 21588 16730
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21560 15201 21588 15982
rect 21546 15192 21602 15201
rect 21546 15127 21602 15136
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21468 14618 21496 14894
rect 21560 14793 21588 14894
rect 21546 14784 21602 14793
rect 21546 14719 21602 14728
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13394 21404 13670
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21376 13161 21404 13194
rect 21362 13152 21418 13161
rect 21362 13087 21418 13096
rect 21468 12481 21496 14282
rect 21546 13696 21602 13705
rect 21546 13631 21602 13640
rect 21560 12889 21588 13631
rect 21546 12880 21602 12889
rect 21546 12815 21602 12824
rect 21546 12608 21602 12617
rect 21546 12543 21602 12552
rect 21454 12472 21510 12481
rect 21454 12407 21510 12416
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21180 11688 21232 11694
rect 21100 11648 21180 11676
rect 21180 11630 21232 11636
rect 21454 11656 21510 11665
rect 21454 11591 21510 11600
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21100 11014 21128 11494
rect 21468 11150 21496 11591
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21100 10470 21128 10950
rect 21560 10470 21588 12543
rect 21652 11354 21680 17002
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21744 14822 21772 15098
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21744 14006 21772 14758
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 21744 13297 21772 13806
rect 21730 13288 21786 13297
rect 21730 13223 21786 13232
rect 21730 12608 21786 12617
rect 21730 12543 21786 12552
rect 21744 12102 21772 12543
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21836 11286 21864 16458
rect 21928 11762 21956 19128
rect 22020 18698 22048 19196
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 22020 16998 22048 17818
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22008 16720 22060 16726
rect 22112 16708 22140 19314
rect 22204 18358 22232 19382
rect 22296 18630 22324 19910
rect 22480 18902 22508 19926
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22296 16833 22324 18566
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22388 17746 22416 18158
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22480 17524 22508 17682
rect 22388 17496 22508 17524
rect 22282 16824 22338 16833
rect 22282 16759 22338 16768
rect 22060 16680 22140 16708
rect 22388 16697 22416 17496
rect 22468 16992 22520 16998
rect 22466 16960 22468 16969
rect 22520 16960 22522 16969
rect 22466 16895 22522 16904
rect 22572 16810 22600 21626
rect 22664 19514 22692 22578
rect 22744 22568 22796 22574
rect 22928 22568 22980 22574
rect 22796 22528 22876 22556
rect 22744 22510 22796 22516
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22756 20262 22784 21626
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22756 19961 22784 20198
rect 22742 19952 22798 19961
rect 22742 19887 22798 19896
rect 22848 19854 22876 22528
rect 22928 22510 22980 22516
rect 22940 22409 22968 22510
rect 23112 22432 23164 22438
rect 22926 22400 22982 22409
rect 22926 22335 22982 22344
rect 23110 22400 23112 22409
rect 23164 22400 23166 22409
rect 23110 22335 23166 22344
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22756 18902 22784 19790
rect 22940 19786 22968 22335
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23032 21350 23060 21830
rect 23216 21350 23244 23530
rect 23308 21962 23336 25486
rect 23386 25392 23442 25401
rect 23386 25327 23442 25336
rect 23400 24041 23428 25327
rect 23492 24449 23520 26250
rect 23584 25265 23612 26318
rect 23676 25498 23704 26438
rect 23768 25514 23796 26574
rect 23846 26551 23902 26560
rect 23860 26382 23888 26551
rect 23952 26382 23980 26998
rect 24412 26994 24440 27950
rect 24030 26959 24086 26968
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24124 26920 24176 26926
rect 24124 26862 24176 26868
rect 24136 26625 24164 26862
rect 24122 26616 24178 26625
rect 24122 26551 24178 26560
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 23940 26376 23992 26382
rect 24228 26353 24256 26930
rect 24308 26920 24360 26926
rect 24306 26888 24308 26897
rect 24360 26888 24362 26897
rect 24306 26823 24362 26832
rect 24400 26852 24452 26858
rect 24400 26794 24452 26800
rect 23940 26318 23992 26324
rect 24214 26344 24270 26353
rect 23952 26228 23980 26318
rect 24214 26279 24270 26288
rect 23860 26200 23980 26228
rect 23860 25650 23888 26200
rect 23996 26140 24304 26149
rect 23996 26138 24002 26140
rect 24058 26138 24082 26140
rect 24138 26138 24162 26140
rect 24218 26138 24242 26140
rect 24298 26138 24304 26140
rect 24058 26086 24060 26138
rect 24240 26086 24242 26138
rect 23996 26084 24002 26086
rect 24058 26084 24082 26086
rect 24138 26084 24162 26086
rect 24218 26084 24242 26086
rect 24298 26084 24304 26086
rect 23996 26075 24304 26084
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 24214 25800 24270 25809
rect 23860 25622 23980 25650
rect 23664 25492 23716 25498
rect 23768 25486 23888 25514
rect 23952 25498 23980 25622
rect 23664 25434 23716 25440
rect 23756 25424 23808 25430
rect 23662 25392 23718 25401
rect 23756 25366 23808 25372
rect 23662 25327 23718 25336
rect 23570 25256 23626 25265
rect 23570 25191 23626 25200
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23584 24993 23612 25094
rect 23570 24984 23626 24993
rect 23570 24919 23626 24928
rect 23572 24880 23624 24886
rect 23572 24822 23624 24828
rect 23478 24440 23534 24449
rect 23478 24375 23534 24384
rect 23584 24342 23612 24822
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 23676 24206 23704 25327
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23572 24064 23624 24070
rect 23386 24032 23442 24041
rect 23768 24052 23796 25366
rect 23860 24886 23888 25486
rect 23940 25492 23992 25498
rect 23940 25434 23992 25440
rect 24044 25265 24072 25774
rect 24214 25735 24270 25744
rect 24122 25528 24178 25537
rect 24122 25463 24124 25472
rect 24176 25463 24178 25472
rect 24124 25434 24176 25440
rect 24030 25256 24086 25265
rect 24030 25191 24086 25200
rect 24228 25158 24256 25735
rect 24306 25392 24362 25401
rect 24306 25327 24362 25336
rect 24320 25294 24348 25327
rect 24308 25288 24360 25294
rect 24308 25230 24360 25236
rect 24216 25152 24268 25158
rect 24412 25129 24440 26794
rect 24504 25974 24532 30359
rect 24596 28694 24624 30620
rect 24676 30602 24728 30608
rect 24872 30308 24900 31078
rect 24964 30938 24992 31583
rect 25056 31210 25084 32166
rect 25044 31204 25096 31210
rect 25044 31146 25096 31152
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 24950 30560 25006 30569
rect 24950 30495 25006 30504
rect 24964 30394 24992 30495
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 24780 30280 24900 30308
rect 24676 30252 24728 30258
rect 24780 30240 24808 30280
rect 24952 30252 25004 30258
rect 24728 30212 24808 30240
rect 24872 30212 24952 30240
rect 24676 30194 24728 30200
rect 24768 30116 24820 30122
rect 24872 30104 24900 30212
rect 24952 30194 25004 30200
rect 24820 30076 24900 30104
rect 24950 30152 25006 30161
rect 24950 30087 25006 30096
rect 24768 30058 24820 30064
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24688 29753 24716 29990
rect 24766 29880 24822 29889
rect 24766 29815 24822 29824
rect 24860 29844 24912 29850
rect 24674 29744 24730 29753
rect 24674 29679 24730 29688
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24688 29345 24716 29582
rect 24674 29336 24730 29345
rect 24674 29271 24730 29280
rect 24780 29209 24808 29815
rect 24860 29786 24912 29792
rect 24872 29753 24900 29786
rect 24858 29744 24914 29753
rect 24858 29679 24914 29688
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24766 29200 24822 29209
rect 24676 29164 24728 29170
rect 24766 29135 24822 29144
rect 24676 29106 24728 29112
rect 24584 28688 24636 28694
rect 24584 28630 24636 28636
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24596 28257 24624 28494
rect 24582 28248 24638 28257
rect 24582 28183 24638 28192
rect 24584 28008 24636 28014
rect 24584 27950 24636 27956
rect 24596 27713 24624 27950
rect 24688 27849 24716 29106
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24674 27840 24730 27849
rect 24674 27775 24730 27784
rect 24582 27704 24638 27713
rect 24582 27639 24638 27648
rect 24584 27532 24636 27538
rect 24584 27474 24636 27480
rect 24596 26314 24624 27474
rect 24674 27432 24730 27441
rect 24674 27367 24730 27376
rect 24584 26308 24636 26314
rect 24584 26250 24636 26256
rect 24688 26246 24716 27367
rect 24676 26240 24728 26246
rect 24596 26188 24676 26194
rect 24596 26182 24728 26188
rect 24596 26166 24716 26182
rect 24492 25968 24544 25974
rect 24492 25910 24544 25916
rect 24490 25528 24546 25537
rect 24490 25463 24546 25472
rect 24504 25265 24532 25463
rect 24596 25430 24624 26166
rect 24780 26081 24808 28494
rect 24872 28200 24900 29582
rect 24964 29481 24992 30087
rect 24950 29472 25006 29481
rect 24950 29407 25006 29416
rect 24950 29200 25006 29209
rect 24950 29135 24952 29144
rect 25004 29135 25006 29144
rect 24952 29106 25004 29112
rect 25056 28694 25084 30330
rect 25148 29170 25176 32438
rect 25240 32230 25268 32778
rect 25332 32434 25360 34575
rect 26054 34350 26110 35150
rect 27250 34350 27306 35150
rect 28446 34350 28502 35150
rect 29090 34368 29146 34377
rect 25412 33244 25464 33250
rect 25412 33186 25464 33192
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25240 32026 25268 32166
rect 25228 32020 25280 32026
rect 25424 32008 25452 33186
rect 25688 33176 25740 33182
rect 25688 33118 25740 33124
rect 25228 31962 25280 31968
rect 25332 31980 25452 32008
rect 25226 31376 25282 31385
rect 25226 31311 25282 31320
rect 25240 30938 25268 31311
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 25228 30592 25280 30598
rect 25228 30534 25280 30540
rect 25240 30433 25268 30534
rect 25226 30424 25282 30433
rect 25332 30394 25360 31980
rect 25410 31920 25466 31929
rect 25410 31855 25466 31864
rect 25226 30359 25282 30368
rect 25320 30388 25372 30394
rect 25320 30330 25372 30336
rect 25424 30274 25452 31855
rect 25504 31136 25556 31142
rect 25502 31104 25504 31113
rect 25556 31104 25558 31113
rect 25502 31039 25558 31048
rect 25504 30592 25556 30598
rect 25556 30552 25636 30580
rect 25504 30534 25556 30540
rect 25504 30388 25556 30394
rect 25504 30330 25556 30336
rect 25332 30246 25452 30274
rect 25516 30258 25544 30330
rect 25504 30252 25556 30258
rect 25228 30184 25280 30190
rect 25226 30152 25228 30161
rect 25280 30152 25282 30161
rect 25226 30087 25282 30096
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 25240 29753 25268 29786
rect 25226 29744 25282 29753
rect 25226 29679 25282 29688
rect 25226 29472 25282 29481
rect 25226 29407 25282 29416
rect 25240 29238 25268 29407
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 25136 29164 25188 29170
rect 25136 29106 25188 29112
rect 25228 29096 25280 29102
rect 25228 29038 25280 29044
rect 24952 28688 25004 28694
rect 24952 28630 25004 28636
rect 25044 28688 25096 28694
rect 25044 28630 25096 28636
rect 24964 28540 24992 28630
rect 24964 28512 25084 28540
rect 25056 28506 25084 28512
rect 25056 28478 25176 28506
rect 24872 28172 25084 28200
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24872 27674 24900 27814
rect 24860 27668 24912 27674
rect 24860 27610 24912 27616
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24766 26072 24822 26081
rect 24766 26007 24822 26016
rect 24872 25956 24900 27270
rect 24964 26625 24992 28018
rect 24950 26616 25006 26625
rect 25056 26586 25084 28172
rect 25148 27169 25176 28478
rect 25240 28082 25268 29038
rect 25332 28966 25360 30246
rect 25504 30194 25556 30200
rect 25412 30184 25464 30190
rect 25608 30138 25636 30552
rect 25412 30126 25464 30132
rect 25320 28960 25372 28966
rect 25320 28902 25372 28908
rect 25320 28620 25372 28626
rect 25320 28562 25372 28568
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25228 27872 25280 27878
rect 25226 27840 25228 27849
rect 25280 27840 25282 27849
rect 25226 27775 25282 27784
rect 25332 27713 25360 28562
rect 25424 28558 25452 30126
rect 25516 30110 25636 30138
rect 25412 28552 25464 28558
rect 25412 28494 25464 28500
rect 25516 28506 25544 30110
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25608 29481 25636 29582
rect 25594 29472 25650 29481
rect 25594 29407 25650 29416
rect 25608 28994 25636 29407
rect 25700 29170 25728 33118
rect 26068 32434 26096 34350
rect 26790 34096 26846 34105
rect 26790 34031 26846 34040
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26516 32360 26568 32366
rect 26516 32302 26568 32308
rect 26528 32026 26556 32302
rect 26332 32020 26384 32026
rect 26332 31962 26384 31968
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 25792 29617 25820 31758
rect 26160 31346 26188 31758
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 25884 30394 25912 31282
rect 26160 30841 26188 31282
rect 26240 30864 26292 30870
rect 26146 30832 26202 30841
rect 26240 30806 26292 30812
rect 26146 30767 26202 30776
rect 25964 30592 26016 30598
rect 25964 30534 26016 30540
rect 25872 30388 25924 30394
rect 25872 30330 25924 30336
rect 25884 29850 25912 30330
rect 25872 29844 25924 29850
rect 25872 29786 25924 29792
rect 25778 29608 25834 29617
rect 25778 29543 25834 29552
rect 25688 29164 25740 29170
rect 25688 29106 25740 29112
rect 25608 28966 25728 28994
rect 25596 28756 25648 28762
rect 25596 28698 25648 28704
rect 25608 28626 25636 28698
rect 25596 28620 25648 28626
rect 25596 28562 25648 28568
rect 25424 28404 25452 28494
rect 25516 28478 25636 28506
rect 25424 28376 25544 28404
rect 25412 28144 25464 28150
rect 25412 28086 25464 28092
rect 25424 28014 25452 28086
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25410 27840 25466 27849
rect 25410 27775 25466 27784
rect 25318 27704 25374 27713
rect 25318 27639 25374 27648
rect 25228 27464 25280 27470
rect 25228 27406 25280 27412
rect 25134 27160 25190 27169
rect 25134 27095 25190 27104
rect 25134 26888 25190 26897
rect 25134 26823 25190 26832
rect 24950 26551 25006 26560
rect 25044 26580 25096 26586
rect 24688 25928 24900 25956
rect 24688 25702 24716 25928
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24676 25696 24728 25702
rect 24676 25638 24728 25644
rect 24780 25514 24808 25774
rect 24964 25752 24992 26551
rect 25044 26522 25096 26528
rect 25148 26382 25176 26823
rect 25136 26376 25188 26382
rect 25042 26344 25098 26353
rect 25136 26318 25188 26324
rect 25042 26279 25098 26288
rect 25056 26042 25084 26279
rect 25044 26036 25096 26042
rect 25044 25978 25096 25984
rect 24688 25486 24808 25514
rect 24872 25724 24992 25752
rect 24872 25498 24900 25724
rect 24950 25664 25006 25673
rect 24950 25599 25006 25608
rect 24964 25498 24992 25599
rect 24860 25492 24912 25498
rect 24584 25424 24636 25430
rect 24584 25366 24636 25372
rect 24584 25288 24636 25294
rect 24490 25256 24546 25265
rect 24688 25276 24716 25486
rect 24860 25434 24912 25440
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24636 25248 24716 25276
rect 24584 25230 24636 25236
rect 24490 25191 24546 25200
rect 24216 25094 24268 25100
rect 24398 25120 24454 25129
rect 23996 25052 24304 25061
rect 24398 25055 24454 25064
rect 23996 25050 24002 25052
rect 24058 25050 24082 25052
rect 24138 25050 24162 25052
rect 24218 25050 24242 25052
rect 24298 25050 24304 25052
rect 24058 24998 24060 25050
rect 24240 24998 24242 25050
rect 23996 24996 24002 24998
rect 24058 24996 24082 24998
rect 24138 24996 24162 24998
rect 24218 24996 24242 24998
rect 24298 24996 24304 24998
rect 23996 24987 24304 24996
rect 24398 24984 24454 24993
rect 24596 24954 24624 25230
rect 24398 24919 24454 24928
rect 24584 24948 24636 24954
rect 23848 24880 23900 24886
rect 23848 24822 23900 24828
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24320 24290 24348 24550
rect 24412 24410 24440 24919
rect 24584 24890 24636 24896
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24492 24336 24544 24342
rect 24320 24262 24440 24290
rect 24492 24278 24544 24284
rect 23624 24024 23796 24052
rect 23846 24032 23902 24041
rect 23572 24006 23624 24012
rect 23386 23967 23442 23976
rect 23846 23967 23902 23976
rect 23570 23896 23626 23905
rect 23570 23831 23626 23840
rect 23754 23896 23810 23905
rect 23754 23831 23810 23840
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23296 21956 23348 21962
rect 23296 21898 23348 21904
rect 23400 21690 23428 23734
rect 23584 23662 23612 23831
rect 23768 23798 23796 23831
rect 23756 23792 23808 23798
rect 23756 23734 23808 23740
rect 23480 23656 23532 23662
rect 23478 23624 23480 23633
rect 23572 23656 23624 23662
rect 23532 23624 23534 23633
rect 23572 23598 23624 23604
rect 23478 23559 23534 23568
rect 23478 23488 23534 23497
rect 23478 23423 23534 23432
rect 23492 22545 23520 23423
rect 23664 23180 23716 23186
rect 23584 23140 23664 23168
rect 23478 22536 23534 22545
rect 23478 22471 23534 22480
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 23204 21344 23256 21350
rect 23584 21321 23612 23140
rect 23664 23122 23716 23128
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23676 22234 23704 22442
rect 23664 22228 23716 22234
rect 23664 22170 23716 22176
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23676 21690 23704 21966
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23204 21286 23256 21292
rect 23570 21312 23626 21321
rect 23570 21247 23626 21256
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22744 18896 22796 18902
rect 22744 18838 22796 18844
rect 23032 18601 23060 19994
rect 23492 19990 23520 20334
rect 23768 20330 23796 22578
rect 23860 21690 23888 23967
rect 23996 23964 24304 23973
rect 23996 23962 24002 23964
rect 24058 23962 24082 23964
rect 24138 23962 24162 23964
rect 24218 23962 24242 23964
rect 24298 23962 24304 23964
rect 24058 23910 24060 23962
rect 24240 23910 24242 23962
rect 23996 23908 24002 23910
rect 24058 23908 24082 23910
rect 24138 23908 24162 23910
rect 24218 23908 24242 23910
rect 24298 23908 24304 23910
rect 23996 23899 24304 23908
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 24032 23248 24084 23254
rect 24032 23190 24084 23196
rect 24044 22982 24072 23190
rect 24136 23118 24164 23462
rect 24412 23361 24440 24262
rect 24504 23905 24532 24278
rect 24596 24206 24624 24890
rect 24780 24721 24808 25327
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24766 24712 24822 24721
rect 24676 24676 24728 24682
rect 24766 24647 24822 24656
rect 24676 24618 24728 24624
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24490 23896 24546 23905
rect 24490 23831 24546 23840
rect 24398 23352 24454 23361
rect 24398 23287 24454 23296
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 24688 23050 24716 24618
rect 24872 23798 24900 25094
rect 24952 24948 25004 24954
rect 24952 24890 25004 24896
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 24964 23644 24992 24890
rect 25056 24886 25084 25978
rect 25148 25158 25176 26318
rect 25240 25362 25268 27406
rect 25332 27334 25360 27639
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25228 25356 25280 25362
rect 25228 25298 25280 25304
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 25056 24614 25084 24686
rect 25044 24608 25096 24614
rect 25042 24576 25044 24585
rect 25096 24576 25098 24585
rect 25042 24511 25098 24520
rect 25226 24576 25282 24585
rect 25226 24511 25282 24520
rect 25044 24404 25096 24410
rect 25096 24364 25176 24392
rect 25044 24346 25096 24352
rect 25044 24064 25096 24070
rect 25044 24006 25096 24012
rect 24780 23616 24992 23644
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 24582 22944 24638 22953
rect 23996 22876 24304 22885
rect 24582 22879 24638 22888
rect 23996 22874 24002 22876
rect 24058 22874 24082 22876
rect 24138 22874 24162 22876
rect 24218 22874 24242 22876
rect 24298 22874 24304 22876
rect 24058 22822 24060 22874
rect 24240 22822 24242 22874
rect 23996 22820 24002 22822
rect 24058 22820 24082 22822
rect 24138 22820 24162 22822
rect 24218 22820 24242 22822
rect 24298 22820 24304 22822
rect 23996 22811 24304 22820
rect 24596 22642 24624 22879
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24780 22488 24808 23616
rect 25056 23526 25084 24006
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24872 23168 24900 23258
rect 25044 23180 25096 23186
rect 24872 23140 25044 23168
rect 25044 23122 25096 23128
rect 25148 23066 25176 24364
rect 25240 23769 25268 24511
rect 25226 23760 25282 23769
rect 25226 23695 25282 23704
rect 25332 23526 25360 26930
rect 25424 25702 25452 27775
rect 25516 27470 25544 28376
rect 25608 28234 25636 28478
rect 25700 28422 25728 28966
rect 25792 28762 25820 29543
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29238 25912 29446
rect 25872 29232 25924 29238
rect 25872 29174 25924 29180
rect 25884 28762 25912 29174
rect 25780 28756 25832 28762
rect 25780 28698 25832 28704
rect 25872 28756 25924 28762
rect 25872 28698 25924 28704
rect 25778 28656 25834 28665
rect 25778 28591 25780 28600
rect 25832 28591 25834 28600
rect 25780 28562 25832 28568
rect 25780 28484 25832 28490
rect 25780 28426 25832 28432
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25608 28206 25728 28234
rect 25596 27872 25648 27878
rect 25594 27840 25596 27849
rect 25648 27840 25650 27849
rect 25594 27775 25650 27784
rect 25596 27668 25648 27674
rect 25596 27610 25648 27616
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25504 26988 25556 26994
rect 25608 26976 25636 27610
rect 25700 27334 25728 28206
rect 25792 27946 25820 28426
rect 25872 28416 25924 28422
rect 25872 28358 25924 28364
rect 25780 27940 25832 27946
rect 25780 27882 25832 27888
rect 25778 27840 25834 27849
rect 25778 27775 25834 27784
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25556 26948 25636 26976
rect 25504 26930 25556 26936
rect 25516 26217 25544 26930
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25608 26586 25636 26726
rect 25596 26580 25648 26586
rect 25596 26522 25648 26528
rect 25502 26208 25558 26217
rect 25502 26143 25558 26152
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25056 23038 25176 23066
rect 24860 22500 24912 22506
rect 24780 22460 24860 22488
rect 24860 22442 24912 22448
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23952 22273 23980 22374
rect 23938 22264 23994 22273
rect 23938 22199 23994 22208
rect 24676 22228 24728 22234
rect 24676 22170 24728 22176
rect 24492 21956 24544 21962
rect 24492 21898 24544 21904
rect 23996 21788 24304 21797
rect 23996 21786 24002 21788
rect 24058 21786 24082 21788
rect 24138 21786 24162 21788
rect 24218 21786 24242 21788
rect 24298 21786 24304 21788
rect 24058 21734 24060 21786
rect 24240 21734 24242 21786
rect 23996 21732 24002 21734
rect 24058 21732 24082 21734
rect 24138 21732 24162 21734
rect 24218 21732 24242 21734
rect 24298 21732 24304 21734
rect 23996 21723 24304 21732
rect 23848 21684 23900 21690
rect 23848 21626 23900 21632
rect 24504 21321 24532 21898
rect 24584 21888 24636 21894
rect 24688 21865 24716 22170
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24584 21830 24636 21836
rect 24674 21856 24730 21865
rect 24596 21729 24624 21830
rect 24674 21791 24730 21800
rect 24582 21720 24638 21729
rect 24582 21655 24638 21664
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24490 21312 24546 21321
rect 24490 21247 24546 21256
rect 23996 20700 24304 20709
rect 23996 20698 24002 20700
rect 24058 20698 24082 20700
rect 24138 20698 24162 20700
rect 24218 20698 24242 20700
rect 24298 20698 24304 20700
rect 24058 20646 24060 20698
rect 24240 20646 24242 20698
rect 23996 20644 24002 20646
rect 24058 20644 24082 20646
rect 24138 20644 24162 20646
rect 24218 20644 24242 20646
rect 24298 20644 24304 20646
rect 23996 20635 24304 20644
rect 23756 20324 23808 20330
rect 23756 20266 23808 20272
rect 23480 19984 23532 19990
rect 23480 19926 23532 19932
rect 23756 19916 23808 19922
rect 23756 19858 23808 19864
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23110 19000 23166 19009
rect 23110 18935 23166 18944
rect 23124 18737 23152 18935
rect 23216 18834 23244 19450
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23110 18728 23166 18737
rect 23110 18663 23166 18672
rect 23018 18592 23074 18601
rect 23018 18527 23074 18536
rect 22744 18352 22796 18358
rect 22742 18320 22744 18329
rect 22796 18320 22798 18329
rect 22742 18255 22798 18264
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 22928 18080 22980 18086
rect 22928 18022 22980 18028
rect 22940 17746 22968 18022
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22664 17626 22692 17682
rect 22664 17598 22876 17626
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22480 16782 22600 16810
rect 22374 16688 22430 16697
rect 22008 16662 22060 16668
rect 22020 16114 22048 16662
rect 22374 16623 22430 16632
rect 22284 16176 22336 16182
rect 22282 16144 22284 16153
rect 22336 16144 22338 16153
rect 22008 16108 22060 16114
rect 22282 16079 22338 16088
rect 22008 16050 22060 16056
rect 22020 15434 22048 16050
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22020 14822 22048 15370
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22020 14074 22048 14214
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 22020 13938 22048 14010
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22020 13394 22048 13874
rect 22098 13424 22154 13433
rect 22008 13388 22060 13394
rect 22098 13359 22154 13368
rect 22008 13330 22060 13336
rect 22020 12850 22048 13330
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 22020 11286 22048 11834
rect 22112 11626 22140 13359
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 22204 11354 22232 15370
rect 22388 14890 22416 15982
rect 22480 15065 22508 16782
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22466 15056 22522 15065
rect 22466 14991 22522 15000
rect 22376 14884 22428 14890
rect 22376 14826 22428 14832
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 13190 22324 14758
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22388 13297 22416 14486
rect 22480 13841 22508 14991
rect 22466 13832 22522 13841
rect 22466 13767 22522 13776
rect 22374 13288 22430 13297
rect 22374 13223 22430 13232
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22284 12368 22336 12374
rect 22284 12310 22336 12316
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10674 22048 11086
rect 22296 10849 22324 12310
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22388 11830 22416 12038
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22282 10840 22338 10849
rect 22282 10775 22338 10784
rect 22480 10742 22508 12106
rect 22572 10810 22600 16118
rect 22664 14260 22692 17478
rect 22848 17134 22876 17598
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22742 16688 22798 16697
rect 22742 16623 22798 16632
rect 22756 14958 22784 16623
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22848 15162 22876 16458
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22744 14952 22796 14958
rect 22744 14894 22796 14900
rect 22756 14414 22784 14894
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22836 14340 22888 14346
rect 22836 14282 22888 14288
rect 22664 14232 22784 14260
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22664 10810 22692 13194
rect 22756 12374 22784 14232
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11898 22784 12174
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22848 11082 22876 14282
rect 22940 11898 22968 17206
rect 23032 17134 23060 18158
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23032 16697 23060 17070
rect 23018 16688 23074 16697
rect 23018 16623 23074 16632
rect 23018 16552 23074 16561
rect 23018 16487 23074 16496
rect 23032 14482 23060 16487
rect 23124 15722 23152 17818
rect 23202 17776 23258 17785
rect 23202 17711 23258 17720
rect 23216 17105 23244 17711
rect 23202 17096 23258 17105
rect 23202 17031 23258 17040
rect 23308 16402 23336 19654
rect 23400 19514 23428 19790
rect 23570 19544 23626 19553
rect 23388 19508 23440 19514
rect 23570 19479 23626 19488
rect 23388 19450 23440 19456
rect 23386 18728 23442 18737
rect 23386 18663 23442 18672
rect 23400 17241 23428 18663
rect 23584 18358 23612 19479
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23386 17232 23442 17241
rect 23386 17167 23442 17176
rect 23492 16794 23520 18090
rect 23676 18057 23704 18566
rect 23768 18290 23796 19858
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 23996 19612 24304 19621
rect 23996 19610 24002 19612
rect 24058 19610 24082 19612
rect 24138 19610 24162 19612
rect 24218 19610 24242 19612
rect 24298 19610 24304 19612
rect 24058 19558 24060 19610
rect 24240 19558 24242 19610
rect 23996 19556 24002 19558
rect 24058 19556 24082 19558
rect 24138 19556 24162 19558
rect 24218 19556 24242 19558
rect 24298 19556 24304 19558
rect 23996 19547 24304 19556
rect 24596 19553 24624 19790
rect 24582 19544 24638 19553
rect 24582 19479 24638 19488
rect 23848 19440 23900 19446
rect 24688 19394 24716 21490
rect 23848 19382 23900 19388
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23756 18080 23808 18086
rect 23662 18048 23718 18057
rect 23756 18022 23808 18028
rect 23662 17983 23718 17992
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23584 17377 23612 17750
rect 23570 17368 23626 17377
rect 23570 17303 23626 17312
rect 23768 16833 23796 18022
rect 23754 16824 23810 16833
rect 23480 16788 23532 16794
rect 23754 16759 23810 16768
rect 23480 16730 23532 16736
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23308 16374 23428 16402
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23308 16017 23336 16186
rect 23294 16008 23350 16017
rect 23400 15978 23428 16374
rect 23294 15943 23350 15952
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23124 15694 23336 15722
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23032 12238 23060 12718
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22468 10736 22520 10742
rect 22468 10678 22520 10684
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 20902 10231 20958 10240
rect 20996 10260 21048 10266
rect 20720 10202 20772 10208
rect 20916 10130 20944 10231
rect 20996 10202 21048 10208
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 16314 9820 16622 9829
rect 16314 9818 16320 9820
rect 16376 9818 16400 9820
rect 16456 9818 16480 9820
rect 16536 9818 16560 9820
rect 16616 9818 16622 9820
rect 16376 9766 16378 9818
rect 16558 9766 16560 9818
rect 16314 9764 16320 9766
rect 16376 9764 16400 9766
rect 16456 9764 16480 9766
rect 16536 9764 16560 9766
rect 16616 9764 16622 9766
rect 16314 9755 16622 9764
rect 21100 9722 21128 10406
rect 22020 10266 22048 10610
rect 22192 10532 22244 10538
rect 22192 10474 22244 10480
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 22204 10441 22232 10474
rect 22190 10432 22246 10441
rect 22190 10367 22246 10376
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22192 10192 22244 10198
rect 22296 10180 22324 10474
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22244 10152 22324 10180
rect 22192 10134 22244 10140
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22112 9722 22140 9998
rect 22664 9722 22692 10202
rect 23124 10130 23152 15574
rect 23308 11354 23336 15694
rect 23492 15484 23520 16594
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23676 16436 23704 16526
rect 23676 16408 23796 16436
rect 23662 16144 23718 16153
rect 23662 16079 23718 16088
rect 23676 15978 23704 16079
rect 23768 16046 23796 16408
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23572 15972 23624 15978
rect 23572 15914 23624 15920
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23584 15638 23612 15914
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 23756 15496 23808 15502
rect 23492 15456 23612 15484
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23400 13920 23428 15030
rect 23478 14376 23534 14385
rect 23478 14311 23534 14320
rect 23492 14278 23520 14311
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23400 13892 23520 13920
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23400 12238 23428 13738
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23400 11558 23428 12174
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23492 11354 23520 13892
rect 23584 13705 23612 15456
rect 23756 15438 23808 15444
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23676 14074 23704 14758
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23570 13696 23626 13705
rect 23570 13631 23626 13640
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23584 12050 23612 12378
rect 23676 12238 23704 13806
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23584 12022 23704 12050
rect 23570 11928 23626 11937
rect 23570 11863 23572 11872
rect 23624 11863 23626 11872
rect 23572 11834 23624 11840
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23584 11150 23612 11698
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 23216 10538 23244 10746
rect 23676 10674 23704 12022
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 23202 10432 23258 10441
rect 23202 10367 23258 10376
rect 23216 10130 23244 10367
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 23676 10062 23704 10610
rect 23768 10266 23796 15438
rect 23860 14657 23888 19382
rect 24596 19366 24716 19394
rect 24032 19168 24084 19174
rect 24030 19136 24032 19145
rect 24216 19168 24268 19174
rect 24084 19136 24086 19145
rect 24216 19110 24268 19116
rect 24030 19071 24086 19080
rect 24228 18766 24256 19110
rect 24490 19000 24546 19009
rect 24490 18935 24546 18944
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24504 18601 24532 18935
rect 24490 18592 24546 18601
rect 23996 18524 24304 18533
rect 24490 18527 24546 18536
rect 23996 18522 24002 18524
rect 24058 18522 24082 18524
rect 24138 18522 24162 18524
rect 24218 18522 24242 18524
rect 24298 18522 24304 18524
rect 24058 18470 24060 18522
rect 24240 18470 24242 18522
rect 23996 18468 24002 18470
rect 24058 18468 24082 18470
rect 24138 18468 24162 18470
rect 24218 18468 24242 18470
rect 24298 18468 24304 18470
rect 23996 18459 24304 18468
rect 24398 18456 24454 18465
rect 24398 18391 24454 18400
rect 24412 18290 24440 18391
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 23996 17436 24304 17445
rect 23996 17434 24002 17436
rect 24058 17434 24082 17436
rect 24138 17434 24162 17436
rect 24218 17434 24242 17436
rect 24298 17434 24304 17436
rect 24058 17382 24060 17434
rect 24240 17382 24242 17434
rect 23996 17380 24002 17382
rect 24058 17380 24082 17382
rect 24138 17380 24162 17382
rect 24218 17380 24242 17382
rect 24298 17380 24304 17382
rect 23996 17371 24304 17380
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 23952 16794 23980 17274
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 24044 16794 24072 17138
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 24030 16552 24086 16561
rect 24030 16487 24086 16496
rect 24044 16454 24072 16487
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 23996 16348 24304 16357
rect 23996 16346 24002 16348
rect 24058 16346 24082 16348
rect 24138 16346 24162 16348
rect 24218 16346 24242 16348
rect 24298 16346 24304 16348
rect 24058 16294 24060 16346
rect 24240 16294 24242 16346
rect 23996 16292 24002 16294
rect 24058 16292 24082 16294
rect 24138 16292 24162 16294
rect 24218 16292 24242 16294
rect 24298 16292 24304 16294
rect 23996 16283 24304 16292
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23940 16176 23992 16182
rect 23940 16118 23992 16124
rect 23952 15609 23980 16118
rect 23938 15600 23994 15609
rect 23938 15535 23994 15544
rect 24044 15473 24072 16186
rect 24030 15464 24086 15473
rect 24030 15399 24086 15408
rect 23996 15260 24304 15269
rect 23996 15258 24002 15260
rect 24058 15258 24082 15260
rect 24138 15258 24162 15260
rect 24218 15258 24242 15260
rect 24298 15258 24304 15260
rect 24058 15206 24060 15258
rect 24240 15206 24242 15258
rect 23996 15204 24002 15206
rect 24058 15204 24082 15206
rect 24138 15204 24162 15206
rect 24218 15204 24242 15206
rect 24298 15204 24304 15206
rect 23996 15195 24304 15204
rect 23846 14648 23902 14657
rect 23846 14583 23902 14592
rect 23860 14346 24164 14362
rect 23860 14340 24176 14346
rect 23860 14334 24124 14340
rect 23860 14074 23888 14334
rect 24124 14282 24176 14288
rect 23996 14172 24304 14181
rect 23996 14170 24002 14172
rect 24058 14170 24082 14172
rect 24138 14170 24162 14172
rect 24218 14170 24242 14172
rect 24298 14170 24304 14172
rect 24058 14118 24060 14170
rect 24240 14118 24242 14170
rect 23996 14116 24002 14118
rect 24058 14116 24082 14118
rect 24138 14116 24162 14118
rect 24218 14116 24242 14118
rect 24298 14116 24304 14118
rect 23996 14107 24304 14116
rect 23848 14068 23900 14074
rect 24412 14056 24440 18226
rect 24490 18184 24546 18193
rect 24490 18119 24546 18128
rect 24504 17338 24532 18119
rect 24596 17626 24624 19366
rect 24676 18080 24728 18086
rect 24780 18057 24808 21898
rect 24872 19922 24900 22442
rect 24952 21412 25004 21418
rect 24952 21354 25004 21360
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24872 19417 24900 19722
rect 24858 19408 24914 19417
rect 24858 19343 24914 19352
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 24676 18022 24728 18028
rect 24766 18048 24822 18057
rect 24688 17728 24716 18022
rect 24766 17983 24822 17992
rect 24688 17700 24808 17728
rect 24780 17649 24808 17700
rect 24766 17640 24822 17649
rect 24596 17598 24716 17626
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 24504 15745 24532 16458
rect 24490 15736 24546 15745
rect 24490 15671 24546 15680
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24504 14822 24532 15438
rect 24596 15094 24624 17478
rect 24688 17377 24716 17598
rect 24766 17575 24822 17584
rect 24872 17513 24900 19178
rect 24964 18902 24992 21354
rect 25056 20058 25084 23038
rect 25240 22964 25268 23462
rect 25424 23225 25452 24210
rect 25516 24041 25544 26143
rect 25608 26042 25636 26522
rect 25700 26518 25728 27270
rect 25688 26512 25740 26518
rect 25688 26454 25740 26460
rect 25688 26376 25740 26382
rect 25688 26318 25740 26324
rect 25700 26217 25728 26318
rect 25792 26246 25820 27775
rect 25884 27010 25912 28358
rect 25976 27588 26004 30534
rect 26252 30394 26280 30806
rect 26344 30569 26372 31962
rect 26700 31272 26752 31278
rect 26700 31214 26752 31220
rect 26608 31204 26660 31210
rect 26608 31146 26660 31152
rect 26514 30968 26570 30977
rect 26514 30903 26570 30912
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26330 30560 26386 30569
rect 26330 30495 26386 30504
rect 26240 30388 26292 30394
rect 26240 30330 26292 30336
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 26068 30025 26096 30126
rect 26240 30116 26292 30122
rect 26240 30058 26292 30064
rect 26054 30016 26110 30025
rect 26054 29951 26110 29960
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 26056 29776 26108 29782
rect 26056 29718 26108 29724
rect 26068 28082 26096 29718
rect 26160 29617 26188 29786
rect 26146 29608 26202 29617
rect 26252 29578 26280 30058
rect 26330 30016 26386 30025
rect 26330 29951 26386 29960
rect 26344 29850 26372 29951
rect 26332 29844 26384 29850
rect 26332 29786 26384 29792
rect 26332 29708 26384 29714
rect 26332 29650 26384 29656
rect 26146 29543 26202 29552
rect 26240 29572 26292 29578
rect 26240 29514 26292 29520
rect 26146 29472 26202 29481
rect 26146 29407 26202 29416
rect 26160 29220 26188 29407
rect 26252 29345 26280 29514
rect 26238 29336 26294 29345
rect 26344 29306 26372 29650
rect 26238 29271 26294 29280
rect 26332 29300 26384 29306
rect 26332 29242 26384 29248
rect 26160 29192 26280 29220
rect 26148 29028 26200 29034
rect 26148 28970 26200 28976
rect 26160 28082 26188 28970
rect 26252 28558 26280 29192
rect 26332 29096 26384 29102
rect 26332 29038 26384 29044
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 26238 28384 26294 28393
rect 26238 28319 26294 28328
rect 26052 28076 26104 28082
rect 26052 28018 26104 28024
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 26160 27849 26188 28018
rect 26146 27840 26202 27849
rect 26146 27775 26202 27784
rect 26252 27690 26280 28319
rect 26160 27674 26280 27690
rect 26148 27668 26280 27674
rect 26200 27662 26280 27668
rect 26148 27610 26200 27616
rect 26240 27600 26292 27606
rect 25976 27560 26092 27588
rect 26064 27520 26092 27560
rect 26238 27568 26240 27577
rect 26292 27568 26294 27577
rect 26064 27492 26096 27520
rect 26238 27503 26294 27512
rect 25964 27464 26016 27470
rect 25964 27406 26016 27412
rect 25976 27169 26004 27406
rect 25962 27160 26018 27169
rect 25962 27095 26018 27104
rect 25884 26982 26004 27010
rect 25870 26888 25926 26897
rect 25870 26823 25872 26832
rect 25924 26823 25926 26832
rect 25872 26794 25924 26800
rect 25872 26444 25924 26450
rect 25872 26386 25924 26392
rect 25780 26240 25832 26246
rect 25686 26208 25742 26217
rect 25780 26182 25832 26188
rect 25686 26143 25742 26152
rect 25884 26081 25912 26386
rect 25870 26072 25926 26081
rect 25596 26036 25648 26042
rect 25870 26007 25926 26016
rect 25596 25978 25648 25984
rect 25688 25968 25740 25974
rect 25594 25936 25650 25945
rect 25688 25910 25740 25916
rect 25870 25936 25926 25945
rect 25594 25871 25650 25880
rect 25608 24818 25636 25871
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25594 24440 25650 24449
rect 25594 24375 25650 24384
rect 25502 24032 25558 24041
rect 25502 23967 25558 23976
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 25410 23216 25466 23225
rect 25410 23151 25466 23160
rect 25148 22936 25268 22964
rect 25412 22976 25464 22982
rect 25148 22234 25176 22936
rect 25412 22918 25464 22924
rect 25320 22704 25372 22710
rect 25320 22646 25372 22652
rect 25226 22400 25282 22409
rect 25226 22335 25282 22344
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25240 21049 25268 22335
rect 25332 22137 25360 22646
rect 25318 22128 25374 22137
rect 25318 22063 25374 22072
rect 25226 21040 25282 21049
rect 25226 20975 25282 20984
rect 25228 20868 25280 20874
rect 25228 20810 25280 20816
rect 25240 20714 25268 20810
rect 25148 20686 25268 20714
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25042 19816 25098 19825
rect 25042 19751 25098 19760
rect 25056 19417 25084 19751
rect 25042 19408 25098 19417
rect 25042 19343 25098 19352
rect 24952 18896 25004 18902
rect 24952 18838 25004 18844
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24858 17504 24914 17513
rect 24858 17439 24914 17448
rect 24674 17368 24730 17377
rect 24674 17303 24730 17312
rect 24676 17264 24728 17270
rect 24728 17224 24808 17252
rect 24676 17206 24728 17212
rect 24674 16824 24730 16833
rect 24674 16759 24730 16768
rect 24688 15706 24716 16759
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24780 15162 24808 17224
rect 24858 17232 24914 17241
rect 24858 17167 24914 17176
rect 24872 16590 24900 17167
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24858 16416 24914 16425
rect 24858 16351 24914 16360
rect 24872 16250 24900 16351
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24858 16008 24914 16017
rect 24858 15943 24914 15952
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24584 15088 24636 15094
rect 24584 15030 24636 15036
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24490 14648 24546 14657
rect 24490 14583 24546 14592
rect 23848 14010 23900 14016
rect 24320 14028 24440 14056
rect 23860 13938 23888 14010
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 24030 13832 24086 13841
rect 24030 13767 24086 13776
rect 24044 13326 24072 13767
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24228 13394 24256 13670
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24320 13172 24348 14028
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24412 13240 24440 13874
rect 24504 13308 24532 14583
rect 24596 13433 24624 14894
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24780 13938 24808 14418
rect 24872 14278 24900 15943
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24872 14113 24900 14214
rect 24858 14104 24914 14113
rect 24858 14039 24914 14048
rect 24858 13968 24914 13977
rect 24768 13932 24820 13938
rect 24858 13903 24914 13912
rect 24768 13874 24820 13880
rect 24766 13832 24822 13841
rect 24766 13767 24768 13776
rect 24820 13767 24822 13776
rect 24768 13738 24820 13744
rect 24872 13512 24900 13903
rect 24780 13484 24900 13512
rect 24582 13424 24638 13433
rect 24582 13359 24638 13368
rect 24504 13280 24716 13308
rect 24412 13212 24624 13240
rect 23846 13152 23902 13161
rect 24320 13144 24532 13172
rect 23846 13087 23902 13096
rect 23860 12986 23888 13087
rect 23996 13084 24304 13093
rect 23996 13082 24002 13084
rect 24058 13082 24082 13084
rect 24138 13082 24162 13084
rect 24218 13082 24242 13084
rect 24298 13082 24304 13084
rect 24058 13030 24060 13082
rect 24240 13030 24242 13082
rect 23996 13028 24002 13030
rect 24058 13028 24082 13030
rect 24138 13028 24162 13030
rect 24218 13028 24242 13030
rect 24298 13028 24304 13030
rect 23996 13019 24304 13028
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 24214 12880 24270 12889
rect 24214 12815 24216 12824
rect 24268 12815 24270 12824
rect 24216 12786 24268 12792
rect 23846 12472 23902 12481
rect 23846 12407 23902 12416
rect 23860 11898 23888 12407
rect 24228 12186 24256 12786
rect 24400 12708 24452 12714
rect 24400 12650 24452 12656
rect 24412 12442 24440 12650
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24228 12158 24440 12186
rect 23996 11996 24304 12005
rect 23996 11994 24002 11996
rect 24058 11994 24082 11996
rect 24138 11994 24162 11996
rect 24218 11994 24242 11996
rect 24298 11994 24304 11996
rect 24058 11942 24060 11994
rect 24240 11942 24242 11994
rect 23996 11940 24002 11942
rect 24058 11940 24082 11942
rect 24138 11940 24162 11942
rect 24218 11940 24242 11942
rect 24298 11940 24304 11942
rect 23996 11931 24304 11940
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23860 10441 23888 11698
rect 23996 10908 24304 10917
rect 23996 10906 24002 10908
rect 24058 10906 24082 10908
rect 24138 10906 24162 10908
rect 24218 10906 24242 10908
rect 24298 10906 24304 10908
rect 24058 10854 24060 10906
rect 24240 10854 24242 10906
rect 23996 10852 24002 10854
rect 24058 10852 24082 10854
rect 24138 10852 24162 10854
rect 24218 10852 24242 10854
rect 24298 10852 24304 10854
rect 23996 10843 24304 10852
rect 24306 10704 24362 10713
rect 24306 10639 24362 10648
rect 24320 10470 24348 10639
rect 24308 10464 24360 10470
rect 23846 10432 23902 10441
rect 24308 10406 24360 10412
rect 23846 10367 23902 10376
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 23112 9716 23164 9722
rect 23112 9658 23164 9664
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20155 9276 20463 9285
rect 20155 9274 20161 9276
rect 20217 9274 20241 9276
rect 20297 9274 20321 9276
rect 20377 9274 20401 9276
rect 20457 9274 20463 9276
rect 20217 9222 20219 9274
rect 20399 9222 20401 9274
rect 20155 9220 20161 9222
rect 20217 9220 20241 9222
rect 20297 9220 20321 9222
rect 20377 9220 20401 9222
rect 20457 9220 20463 9222
rect 20155 9211 20463 9220
rect 20640 8974 20668 9590
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 21928 8838 21956 9658
rect 23124 9178 23152 9658
rect 23768 9450 23796 10202
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 16314 8732 16622 8741
rect 16314 8730 16320 8732
rect 16376 8730 16400 8732
rect 16456 8730 16480 8732
rect 16536 8730 16560 8732
rect 16616 8730 16622 8732
rect 16376 8678 16378 8730
rect 16558 8678 16560 8730
rect 16314 8676 16320 8678
rect 16376 8676 16400 8678
rect 16456 8676 16480 8678
rect 16536 8676 16560 8678
rect 16616 8676 16622 8678
rect 16314 8667 16622 8676
rect 19522 8664 19578 8673
rect 19522 8599 19578 8608
rect 14280 8424 14332 8430
rect 19536 8401 19564 8599
rect 22572 8430 22600 8774
rect 22940 8498 22968 9114
rect 23124 8634 23152 9114
rect 23860 9042 23888 10367
rect 24320 10146 24348 10406
rect 24412 10266 24440 12158
rect 24504 11914 24532 13144
rect 24596 12102 24624 13212
rect 24688 12442 24716 13280
rect 24780 12782 24808 13484
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24872 12850 24900 13330
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24780 12238 24808 12582
rect 24872 12442 24900 12786
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24964 12374 24992 18702
rect 25056 18290 25084 19343
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 25044 17876 25096 17882
rect 25044 17818 25096 17824
rect 25056 17270 25084 17818
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25056 16425 25084 16526
rect 25042 16416 25098 16425
rect 25042 16351 25098 16360
rect 25044 16176 25096 16182
rect 25044 16118 25096 16124
rect 25056 15337 25084 16118
rect 25042 15328 25098 15337
rect 25042 15263 25098 15272
rect 25044 14340 25096 14346
rect 25044 14282 25096 14288
rect 25056 13802 25084 14282
rect 25044 13796 25096 13802
rect 25044 13738 25096 13744
rect 25042 13016 25098 13025
rect 25042 12951 25098 12960
rect 25056 12850 25084 12951
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24504 11886 24716 11914
rect 24584 11620 24636 11626
rect 24584 11562 24636 11568
rect 24596 11218 24624 11562
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24596 10674 24624 11154
rect 24688 11082 24716 11886
rect 24780 11762 24808 12174
rect 24872 11762 24900 12174
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24688 10810 24716 11018
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24872 10554 24900 11698
rect 24964 11642 24992 12038
rect 25056 11762 25084 12786
rect 25148 12442 25176 20686
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25240 18057 25268 18566
rect 25332 18222 25360 19994
rect 25424 19666 25452 22918
rect 25516 21146 25544 23666
rect 25608 23225 25636 24375
rect 25700 24177 25728 25910
rect 25870 25871 25926 25880
rect 25884 25770 25912 25871
rect 25976 25838 26004 26982
rect 26068 26024 26096 27492
rect 26148 27464 26200 27470
rect 26146 27432 26148 27441
rect 26200 27432 26202 27441
rect 26344 27402 26372 29038
rect 26436 29034 26464 30602
rect 26528 29646 26556 30903
rect 26620 30734 26648 31146
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26608 29844 26660 29850
rect 26608 29786 26660 29792
rect 26516 29640 26568 29646
rect 26516 29582 26568 29588
rect 26514 29472 26570 29481
rect 26514 29407 26570 29416
rect 26528 29170 26556 29407
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26514 29064 26570 29073
rect 26424 29028 26476 29034
rect 26514 28999 26570 29008
rect 26424 28970 26476 28976
rect 26436 28257 26464 28970
rect 26528 28966 26556 28999
rect 26516 28960 26568 28966
rect 26620 28937 26648 29786
rect 26712 29174 26740 31214
rect 26804 30841 26832 34031
rect 27066 32464 27122 32473
rect 27264 32434 27292 34350
rect 29642 34350 29698 35150
rect 30838 34490 30894 35150
rect 30838 34462 30972 34490
rect 30838 34350 30894 34462
rect 29090 34303 29146 34312
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27066 32399 27122 32408
rect 27252 32428 27304 32434
rect 26884 32292 26936 32298
rect 26884 32234 26936 32240
rect 26896 31210 26924 32234
rect 26976 31748 27028 31754
rect 26976 31690 27028 31696
rect 26884 31204 26936 31210
rect 26884 31146 26936 31152
rect 26790 30832 26846 30841
rect 26790 30767 26846 30776
rect 26896 30546 26924 31146
rect 26804 30518 26924 30546
rect 26804 30326 26832 30518
rect 26884 30388 26936 30394
rect 26884 30330 26936 30336
rect 26792 30320 26844 30326
rect 26792 30262 26844 30268
rect 26792 30116 26844 30122
rect 26792 30058 26844 30064
rect 26804 29889 26832 30058
rect 26790 29880 26846 29889
rect 26790 29815 26846 29824
rect 26712 29146 26832 29174
rect 26804 29102 26832 29146
rect 26792 29096 26844 29102
rect 26792 29038 26844 29044
rect 26700 29028 26752 29034
rect 26700 28970 26752 28976
rect 26516 28902 26568 28908
rect 26606 28928 26662 28937
rect 26606 28863 26662 28872
rect 26606 28792 26662 28801
rect 26516 28756 26568 28762
rect 26712 28778 26740 28970
rect 26792 28960 26844 28966
rect 26790 28928 26792 28937
rect 26844 28928 26846 28937
rect 26790 28863 26846 28872
rect 26790 28792 26846 28801
rect 26712 28750 26790 28778
rect 26606 28727 26662 28736
rect 26896 28762 26924 30330
rect 26988 29850 27016 31690
rect 27080 31249 27108 32399
rect 27252 32370 27304 32376
rect 27540 32366 27568 33458
rect 27620 33312 27672 33318
rect 27620 33254 27672 33260
rect 27528 32360 27580 32366
rect 27528 32302 27580 32308
rect 27434 32192 27490 32201
rect 27434 32127 27490 32136
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27066 31240 27122 31249
rect 27066 31175 27122 31184
rect 27080 30258 27108 31175
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 27068 30048 27120 30054
rect 27066 30016 27068 30025
rect 27120 30016 27122 30025
rect 27066 29951 27122 29960
rect 26976 29844 27028 29850
rect 26976 29786 27028 29792
rect 26988 29170 27016 29786
rect 27080 29481 27108 29951
rect 27066 29472 27122 29481
rect 27066 29407 27122 29416
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 26976 28960 27028 28966
rect 26976 28902 27028 28908
rect 26988 28762 27016 28902
rect 26790 28727 26846 28736
rect 26884 28756 26936 28762
rect 26516 28698 26568 28704
rect 26422 28248 26478 28257
rect 26422 28183 26478 28192
rect 26422 27976 26478 27985
rect 26422 27911 26478 27920
rect 26436 27588 26464 27911
rect 26528 27849 26556 28698
rect 26620 28393 26648 28727
rect 26884 28698 26936 28704
rect 26976 28756 27028 28762
rect 26976 28698 27028 28704
rect 26792 28688 26844 28694
rect 26844 28636 26924 28642
rect 26792 28630 26924 28636
rect 26804 28614 26924 28630
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 26606 28384 26662 28393
rect 26606 28319 26662 28328
rect 26804 28257 26832 28494
rect 26896 28422 26924 28614
rect 27080 28608 27108 28970
rect 26988 28580 27108 28608
rect 26884 28416 26936 28422
rect 26884 28358 26936 28364
rect 26790 28248 26846 28257
rect 26790 28183 26846 28192
rect 26608 28144 26660 28150
rect 26608 28086 26660 28092
rect 26700 28144 26752 28150
rect 26700 28086 26752 28092
rect 26620 28014 26648 28086
rect 26608 28008 26660 28014
rect 26608 27950 26660 27956
rect 26712 27878 26740 28086
rect 26988 28082 27016 28580
rect 27068 28416 27120 28422
rect 27068 28358 27120 28364
rect 26792 28076 26844 28082
rect 26792 28018 26844 28024
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 26804 27985 26832 28018
rect 26790 27976 26846 27985
rect 26790 27911 26846 27920
rect 26884 27940 26936 27946
rect 26884 27882 26936 27888
rect 26700 27872 26752 27878
rect 26514 27840 26570 27849
rect 26792 27872 26844 27878
rect 26700 27814 26752 27820
rect 26790 27840 26792 27849
rect 26844 27840 26846 27849
rect 26514 27775 26570 27784
rect 26790 27775 26846 27784
rect 26896 27606 26924 27882
rect 26974 27704 27030 27713
rect 26974 27639 27030 27648
rect 26988 27606 27016 27639
rect 26884 27600 26936 27606
rect 26436 27560 26740 27588
rect 26146 27367 26202 27376
rect 26332 27396 26384 27402
rect 26160 27130 26188 27367
rect 26608 27396 26660 27402
rect 26332 27338 26384 27344
rect 26528 27356 26608 27384
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26344 26994 26372 27338
rect 26422 27296 26478 27305
rect 26422 27231 26478 27240
rect 26436 26994 26464 27231
rect 26332 26988 26384 26994
rect 26332 26930 26384 26936
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26238 26888 26294 26897
rect 26238 26823 26294 26832
rect 26252 26790 26280 26823
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26148 26376 26200 26382
rect 26200 26336 26280 26364
rect 26148 26318 26200 26324
rect 26068 25996 26188 26024
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 25964 25832 26016 25838
rect 25964 25774 26016 25780
rect 25872 25764 25924 25770
rect 25872 25706 25924 25712
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25976 25430 26004 25638
rect 25964 25424 26016 25430
rect 25964 25366 26016 25372
rect 25778 25120 25834 25129
rect 25778 25055 25834 25064
rect 25792 24614 25820 25055
rect 25962 24848 26018 24857
rect 25872 24812 25924 24818
rect 25962 24783 26018 24792
rect 25872 24754 25924 24760
rect 25884 24721 25912 24754
rect 25870 24712 25926 24721
rect 25870 24647 25926 24656
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 25870 24440 25926 24449
rect 25870 24375 25926 24384
rect 25884 24342 25912 24375
rect 25872 24336 25924 24342
rect 25872 24278 25924 24284
rect 25976 24206 26004 24783
rect 25964 24200 26016 24206
rect 25686 24168 25742 24177
rect 25964 24142 26016 24148
rect 25686 24103 25742 24112
rect 25688 23792 25740 23798
rect 25686 23760 25688 23769
rect 25872 23792 25924 23798
rect 25740 23760 25742 23769
rect 25872 23734 25924 23740
rect 25686 23695 25742 23704
rect 25884 23633 25912 23734
rect 26068 23730 26096 25842
rect 26160 25838 26188 25996
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 26148 25696 26200 25702
rect 26148 25638 26200 25644
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 25870 23624 25926 23633
rect 25870 23559 25926 23568
rect 26160 23338 26188 25638
rect 26252 24154 26280 26336
rect 26344 24868 26372 26930
rect 26436 26518 26464 26930
rect 26424 26512 26476 26518
rect 26424 26454 26476 26460
rect 26424 26376 26476 26382
rect 26424 26318 26476 26324
rect 26436 25498 26464 26318
rect 26528 25974 26556 27356
rect 26608 27338 26660 27344
rect 26712 27282 26740 27560
rect 26620 27254 26740 27282
rect 26804 27560 26884 27588
rect 26620 26382 26648 27254
rect 26804 26926 26832 27560
rect 26884 27542 26936 27548
rect 26976 27600 27028 27606
rect 27080 27577 27108 28358
rect 26976 27542 27028 27548
rect 27066 27568 27122 27577
rect 27066 27503 27122 27512
rect 27080 27418 27108 27503
rect 26988 27390 27108 27418
rect 26988 27334 27016 27390
rect 26976 27328 27028 27334
rect 26896 27288 26976 27316
rect 26896 26994 26924 27288
rect 26976 27270 27028 27276
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 26974 27160 27030 27169
rect 26974 27095 27030 27104
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 26792 26920 26844 26926
rect 26698 26888 26754 26897
rect 26792 26862 26844 26868
rect 26698 26823 26754 26832
rect 26712 26518 26740 26823
rect 26792 26784 26844 26790
rect 26792 26726 26844 26732
rect 26884 26784 26936 26790
rect 26884 26726 26936 26732
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 26608 26376 26660 26382
rect 26608 26318 26660 26324
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 26516 25832 26568 25838
rect 26514 25800 26516 25809
rect 26568 25800 26570 25809
rect 26514 25735 26570 25744
rect 26514 25664 26570 25673
rect 26514 25599 26570 25608
rect 26424 25492 26476 25498
rect 26424 25434 26476 25440
rect 26424 25152 26476 25158
rect 26424 25094 26476 25100
rect 26436 24993 26464 25094
rect 26422 24984 26478 24993
rect 26528 24954 26556 25599
rect 26422 24919 26478 24928
rect 26516 24948 26568 24954
rect 26516 24890 26568 24896
rect 26344 24840 26464 24868
rect 26252 24126 26372 24154
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26252 23798 26280 24006
rect 26240 23792 26292 23798
rect 26240 23734 26292 23740
rect 26344 23633 26372 24126
rect 26330 23624 26386 23633
rect 26330 23559 26386 23568
rect 26160 23310 26280 23338
rect 25594 23216 25650 23225
rect 25594 23151 25650 23160
rect 26056 23044 26108 23050
rect 26056 22986 26108 22992
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25596 22092 25648 22098
rect 25596 22034 25648 22040
rect 25608 21146 25636 22034
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25596 21140 25648 21146
rect 25596 21082 25648 21088
rect 25516 20641 25544 21082
rect 25502 20632 25558 20641
rect 25700 20618 25728 22918
rect 25964 22704 26016 22710
rect 25964 22646 26016 22652
rect 25976 22574 26004 22646
rect 25964 22568 26016 22574
rect 25964 22510 26016 22516
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25792 21049 25820 22170
rect 25872 21956 25924 21962
rect 25872 21898 25924 21904
rect 25778 21040 25834 21049
rect 25778 20975 25834 20984
rect 25608 20602 25728 20618
rect 25502 20567 25558 20576
rect 25596 20596 25728 20602
rect 25648 20590 25728 20596
rect 25596 20538 25648 20544
rect 25688 20528 25740 20534
rect 25688 20470 25740 20476
rect 25700 19825 25728 20470
rect 25884 20398 25912 21898
rect 26068 20806 26096 22986
rect 26148 22228 26200 22234
rect 26252 22216 26280 23310
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 26344 22642 26372 23054
rect 26436 22982 26464 24840
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 26528 23746 26556 24754
rect 26620 23905 26648 26318
rect 26712 25226 26740 26454
rect 26804 26217 26832 26726
rect 26790 26208 26846 26217
rect 26790 26143 26846 26152
rect 26700 25220 26752 25226
rect 26700 25162 26752 25168
rect 26698 25120 26754 25129
rect 26698 25055 26754 25064
rect 26712 24954 26740 25055
rect 26700 24948 26752 24954
rect 26700 24890 26752 24896
rect 26804 24886 26832 26143
rect 26792 24880 26844 24886
rect 26792 24822 26844 24828
rect 26698 24576 26754 24585
rect 26698 24511 26754 24520
rect 26712 24410 26740 24511
rect 26700 24404 26752 24410
rect 26700 24346 26752 24352
rect 26790 24168 26846 24177
rect 26790 24103 26846 24112
rect 26606 23896 26662 23905
rect 26606 23831 26662 23840
rect 26804 23798 26832 24103
rect 26896 24018 26924 26726
rect 26988 25514 27016 27095
rect 27080 26790 27108 27270
rect 27068 26784 27120 26790
rect 27068 26726 27120 26732
rect 27066 26616 27122 26625
rect 27066 26551 27122 26560
rect 27080 26382 27108 26551
rect 27172 26382 27200 31282
rect 27252 31136 27304 31142
rect 27344 31136 27396 31142
rect 27252 31078 27304 31084
rect 27342 31104 27344 31113
rect 27396 31104 27398 31113
rect 27264 28966 27292 31078
rect 27342 31039 27398 31048
rect 27448 30734 27476 32127
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27436 30728 27488 30734
rect 27342 30696 27398 30705
rect 27436 30670 27488 30676
rect 27342 30631 27398 30640
rect 27356 30054 27384 30631
rect 27448 30190 27476 30670
rect 27436 30184 27488 30190
rect 27436 30126 27488 30132
rect 27344 30048 27396 30054
rect 27344 29990 27396 29996
rect 27356 29889 27384 29990
rect 27342 29880 27398 29889
rect 27342 29815 27398 29824
rect 27448 29714 27476 30126
rect 27540 29714 27568 31962
rect 27436 29708 27488 29714
rect 27436 29650 27488 29656
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27344 29504 27396 29510
rect 27344 29446 27396 29452
rect 27434 29472 27490 29481
rect 27252 28960 27304 28966
rect 27252 28902 27304 28908
rect 27264 26994 27292 28902
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 27068 25900 27120 25906
rect 27264 25888 27292 26930
rect 27120 25860 27292 25888
rect 27068 25842 27120 25848
rect 27356 25820 27384 29446
rect 27434 29407 27490 29416
rect 27448 29034 27476 29407
rect 27526 29336 27582 29345
rect 27526 29271 27582 29280
rect 27540 29238 27568 29271
rect 27528 29232 27580 29238
rect 27528 29174 27580 29180
rect 27632 29102 27660 33254
rect 28172 32496 28224 32502
rect 28172 32438 28224 32444
rect 27837 32124 28145 32133
rect 27837 32122 27843 32124
rect 27899 32122 27923 32124
rect 27979 32122 28003 32124
rect 28059 32122 28083 32124
rect 28139 32122 28145 32124
rect 27899 32070 27901 32122
rect 28081 32070 28083 32122
rect 27837 32068 27843 32070
rect 27899 32068 27923 32070
rect 27979 32068 28003 32070
rect 28059 32068 28083 32070
rect 28139 32068 28145 32070
rect 27710 32056 27766 32065
rect 27837 32059 28145 32068
rect 27710 31991 27766 32000
rect 27724 31890 27752 31991
rect 27712 31884 27764 31890
rect 27712 31826 27764 31832
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 27724 29832 27752 31690
rect 27837 31036 28145 31045
rect 27837 31034 27843 31036
rect 27899 31034 27923 31036
rect 27979 31034 28003 31036
rect 28059 31034 28083 31036
rect 28139 31034 28145 31036
rect 27899 30982 27901 31034
rect 28081 30982 28083 31034
rect 27837 30980 27843 30982
rect 27899 30980 27923 30982
rect 27979 30980 28003 30982
rect 28059 30980 28083 30982
rect 28139 30980 28145 30982
rect 27837 30971 28145 30980
rect 28184 30818 28212 32438
rect 28354 32328 28410 32337
rect 28354 32263 28356 32272
rect 28408 32263 28410 32272
rect 28356 32234 28408 32240
rect 28724 31748 28776 31754
rect 28724 31690 28776 31696
rect 28264 31476 28316 31482
rect 28264 31418 28316 31424
rect 28092 30790 28212 30818
rect 27894 30424 27950 30433
rect 27894 30359 27950 30368
rect 27988 30388 28040 30394
rect 27908 30190 27936 30359
rect 27988 30330 28040 30336
rect 28000 30258 28028 30330
rect 27988 30252 28040 30258
rect 27988 30194 28040 30200
rect 27896 30184 27948 30190
rect 27896 30126 27948 30132
rect 28092 30054 28120 30790
rect 28172 30728 28224 30734
rect 28172 30670 28224 30676
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 27837 29948 28145 29957
rect 27837 29946 27843 29948
rect 27899 29946 27923 29948
rect 27979 29946 28003 29948
rect 28059 29946 28083 29948
rect 28139 29946 28145 29948
rect 27899 29894 27901 29946
rect 28081 29894 28083 29946
rect 27837 29892 27843 29894
rect 27899 29892 27923 29894
rect 27979 29892 28003 29894
rect 28059 29892 28083 29894
rect 28139 29892 28145 29894
rect 27837 29883 28145 29892
rect 27724 29804 27844 29832
rect 27712 29708 27764 29714
rect 27712 29650 27764 29656
rect 27724 29102 27752 29650
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27712 29096 27764 29102
rect 27712 29038 27764 29044
rect 27436 29028 27488 29034
rect 27436 28970 27488 28976
rect 27620 28960 27672 28966
rect 27816 28948 27844 29804
rect 28078 29744 28134 29753
rect 28078 29679 28134 29688
rect 28092 29646 28120 29679
rect 27896 29640 27948 29646
rect 28080 29640 28132 29646
rect 27896 29582 27948 29588
rect 27986 29608 28042 29617
rect 27908 29186 27936 29582
rect 28080 29582 28132 29588
rect 27986 29543 28042 29552
rect 28000 29492 28028 29543
rect 28000 29464 28120 29492
rect 27988 29300 28040 29306
rect 28092 29288 28120 29464
rect 28040 29260 28120 29288
rect 27988 29242 28040 29248
rect 27908 29158 28120 29186
rect 27620 28902 27672 28908
rect 27724 28920 27844 28948
rect 28092 28948 28120 29158
rect 28184 29016 28212 30670
rect 28276 29753 28304 31418
rect 28736 31113 28764 31690
rect 28816 31680 28868 31686
rect 28816 31622 28868 31628
rect 28722 31104 28778 31113
rect 28722 31039 28778 31048
rect 28446 30968 28502 30977
rect 28828 30938 28856 31622
rect 28446 30903 28502 30912
rect 28724 30932 28776 30938
rect 28354 30832 28410 30841
rect 28460 30802 28488 30903
rect 28724 30874 28776 30880
rect 28816 30932 28868 30938
rect 28816 30874 28868 30880
rect 28354 30767 28410 30776
rect 28448 30796 28500 30802
rect 28368 30734 28396 30767
rect 28448 30738 28500 30744
rect 28356 30728 28408 30734
rect 28356 30670 28408 30676
rect 28354 30424 28410 30433
rect 28354 30359 28410 30368
rect 28368 29782 28396 30359
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 28446 29880 28502 29889
rect 28446 29815 28502 29824
rect 28356 29776 28408 29782
rect 28262 29744 28318 29753
rect 28356 29718 28408 29724
rect 28262 29679 28318 29688
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 28262 29472 28318 29481
rect 28262 29407 28318 29416
rect 28276 29306 28304 29407
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 28368 29186 28396 29514
rect 28460 29306 28488 29815
rect 28448 29300 28500 29306
rect 28448 29242 28500 29248
rect 28368 29170 28404 29186
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 28184 28988 28396 29016
rect 28092 28937 28304 28948
rect 28092 28928 28318 28937
rect 28092 28920 28262 28928
rect 27526 28792 27582 28801
rect 27526 28727 27582 28736
rect 27436 27872 27488 27878
rect 27436 27814 27488 27820
rect 27448 26234 27476 27814
rect 27540 27470 27568 28727
rect 27632 28422 27660 28902
rect 27724 28490 27752 28920
rect 27837 28860 28145 28869
rect 28262 28863 28318 28872
rect 27837 28858 27843 28860
rect 27899 28858 27923 28860
rect 27979 28858 28003 28860
rect 28059 28858 28083 28860
rect 28139 28858 28145 28860
rect 27899 28806 27901 28858
rect 28081 28806 28083 28858
rect 27837 28804 27843 28806
rect 27899 28804 27923 28806
rect 27979 28804 28003 28806
rect 28059 28804 28083 28806
rect 28139 28804 28145 28806
rect 27837 28795 28145 28804
rect 28368 28744 28396 28988
rect 28460 28801 28488 29106
rect 28092 28716 28396 28744
rect 28446 28792 28502 28801
rect 28446 28727 28502 28736
rect 27804 28552 27856 28558
rect 27804 28494 27856 28500
rect 27712 28484 27764 28490
rect 27712 28426 27764 28432
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27632 27713 27660 28018
rect 27816 28014 27844 28494
rect 27896 28484 27948 28490
rect 27896 28426 27948 28432
rect 27804 28008 27856 28014
rect 27804 27950 27856 27956
rect 27908 27860 27936 28426
rect 27988 28212 28040 28218
rect 27988 28154 28040 28160
rect 28000 27928 28028 28154
rect 28092 28082 28120 28716
rect 28184 28614 28396 28642
rect 28184 28218 28212 28614
rect 28368 28608 28396 28614
rect 28552 28608 28580 30194
rect 28632 30048 28684 30054
rect 28632 29990 28684 29996
rect 28644 29714 28672 29990
rect 28632 29708 28684 29714
rect 28632 29650 28684 29656
rect 28632 29572 28684 29578
rect 28632 29514 28684 29520
rect 28644 29306 28672 29514
rect 28632 29300 28684 29306
rect 28632 29242 28684 29248
rect 28632 29096 28684 29102
rect 28632 29038 28684 29044
rect 28368 28580 28580 28608
rect 28264 28552 28316 28558
rect 28264 28494 28316 28500
rect 28276 28422 28304 28494
rect 28368 28478 28580 28506
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28368 28082 28396 28478
rect 28552 28422 28580 28478
rect 28540 28416 28592 28422
rect 28446 28384 28502 28393
rect 28540 28358 28592 28364
rect 28446 28319 28502 28328
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 28000 27900 28396 27928
rect 27710 27840 27766 27849
rect 27908 27832 28205 27860
rect 28177 27826 28205 27832
rect 28258 27840 28314 27849
rect 28177 27798 28258 27826
rect 27710 27775 27766 27784
rect 27618 27704 27674 27713
rect 27618 27639 27674 27648
rect 27724 27656 27752 27775
rect 27837 27772 28145 27781
rect 28258 27775 28314 27784
rect 27837 27770 27843 27772
rect 27899 27770 27923 27772
rect 27979 27770 28003 27772
rect 28059 27770 28083 27772
rect 28139 27770 28145 27772
rect 27899 27718 27901 27770
rect 28081 27718 28083 27770
rect 27837 27716 27843 27718
rect 27899 27716 27923 27718
rect 27979 27716 28003 27718
rect 28059 27716 28083 27718
rect 28139 27716 28145 27718
rect 27837 27707 28145 27716
rect 27724 27628 28304 27656
rect 27894 27568 27950 27577
rect 27620 27532 27672 27538
rect 27672 27492 27844 27520
rect 27894 27503 27950 27512
rect 27620 27474 27672 27480
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27816 27402 27844 27492
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 27804 27396 27856 27402
rect 27804 27338 27856 27344
rect 27526 27160 27582 27169
rect 27526 27095 27582 27104
rect 27540 26994 27568 27095
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27540 26790 27568 26930
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 27528 26444 27580 26450
rect 27528 26386 27580 26392
rect 27540 26353 27568 26386
rect 27526 26344 27582 26353
rect 27526 26279 27582 26288
rect 27632 26296 27660 27338
rect 27908 27130 27936 27503
rect 28172 27464 28224 27470
rect 28092 27424 28172 27452
rect 27986 27160 28042 27169
rect 27896 27124 27948 27130
rect 28092 27146 28120 27424
rect 28172 27406 28224 27412
rect 28042 27118 28120 27146
rect 28170 27160 28226 27169
rect 27986 27095 27988 27104
rect 27896 27066 27948 27072
rect 28040 27095 28042 27104
rect 28170 27095 28226 27104
rect 27988 27066 28040 27072
rect 28177 27010 28205 27095
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 28092 26982 28205 27010
rect 28276 27010 28304 27628
rect 28368 27130 28396 27900
rect 28460 27878 28488 28319
rect 28644 28064 28672 29038
rect 28637 28036 28672 28064
rect 28637 27962 28665 28036
rect 28552 27934 28665 27962
rect 28448 27872 28500 27878
rect 28448 27814 28500 27820
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 28276 26982 28396 27010
rect 27724 26450 27752 26930
rect 27908 26790 27936 26930
rect 28092 26790 28120 26982
rect 28368 26976 28396 26982
rect 28368 26948 28404 26976
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 28173 26784 28225 26790
rect 28376 26772 28404 26948
rect 28368 26744 28404 26772
rect 28368 26738 28396 26744
rect 28173 26726 28225 26732
rect 28177 26710 28213 26726
rect 27837 26684 28145 26693
rect 27837 26682 27843 26684
rect 27899 26682 27923 26684
rect 27979 26682 28003 26684
rect 28059 26682 28083 26684
rect 28139 26682 28145 26684
rect 27899 26630 27901 26682
rect 28081 26630 28083 26682
rect 27837 26628 27843 26630
rect 27899 26628 27923 26630
rect 27979 26628 28003 26630
rect 28059 26628 28083 26630
rect 28139 26628 28145 26630
rect 27837 26619 28145 26628
rect 28185 26568 28213 26710
rect 27816 26540 28213 26568
rect 28276 26710 28396 26738
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 27632 26268 27752 26296
rect 27448 26206 27685 26234
rect 27657 26024 27685 26206
rect 27631 25996 27685 26024
rect 27631 25956 27659 25996
rect 27724 25974 27752 26268
rect 27712 25968 27764 25974
rect 27631 25928 27660 25956
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27264 25792 27384 25820
rect 27540 25809 27568 25842
rect 27632 25838 27660 25928
rect 27712 25910 27764 25916
rect 27620 25832 27672 25838
rect 27526 25800 27582 25809
rect 27160 25764 27212 25770
rect 27264 25752 27292 25792
rect 27436 25764 27488 25770
rect 27212 25724 27292 25752
rect 27356 25724 27436 25752
rect 27160 25706 27212 25712
rect 26988 25486 27200 25514
rect 27068 25424 27120 25430
rect 27068 25366 27120 25372
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 26988 25129 27016 25230
rect 26974 25120 27030 25129
rect 26974 25055 27030 25064
rect 27080 24936 27108 25366
rect 27172 25294 27200 25486
rect 27252 25424 27304 25430
rect 27252 25366 27304 25372
rect 27264 25294 27292 25366
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 27252 25288 27304 25294
rect 27252 25230 27304 25236
rect 27080 24908 27200 24936
rect 26976 24880 27028 24886
rect 26976 24822 27028 24828
rect 26988 24585 27016 24822
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 26974 24576 27030 24585
rect 26974 24511 27030 24520
rect 26896 23990 27016 24018
rect 26884 23860 26936 23866
rect 26884 23802 26936 23808
rect 26792 23792 26844 23798
rect 26698 23760 26754 23769
rect 26528 23718 26648 23746
rect 26516 23656 26568 23662
rect 26516 23598 26568 23604
rect 26528 23497 26556 23598
rect 26514 23488 26570 23497
rect 26514 23423 26570 23432
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 26200 22188 26280 22216
rect 26148 22170 26200 22176
rect 26344 22148 26372 22578
rect 26424 22568 26476 22574
rect 26424 22510 26476 22516
rect 26436 22438 26464 22510
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26424 22160 26476 22166
rect 26146 22128 26202 22137
rect 26344 22120 26424 22148
rect 26424 22102 26476 22108
rect 26146 22063 26148 22072
rect 26200 22063 26202 22072
rect 26148 22034 26200 22040
rect 26332 21616 26384 21622
rect 26332 21558 26384 21564
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 26056 20800 26108 20806
rect 26252 20777 26280 20810
rect 26056 20742 26108 20748
rect 26238 20768 26294 20777
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 25686 19816 25742 19825
rect 25686 19751 25742 19760
rect 25424 19638 25544 19666
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25226 18048 25282 18057
rect 25226 17983 25282 17992
rect 25228 17672 25280 17678
rect 25228 17614 25280 17620
rect 25240 16590 25268 17614
rect 25332 17134 25360 18158
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25318 16824 25374 16833
rect 25318 16759 25374 16768
rect 25332 16658 25360 16759
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25228 16584 25280 16590
rect 25424 16561 25452 19450
rect 25516 17882 25544 19638
rect 25792 19553 25820 20198
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25594 19544 25650 19553
rect 25594 19479 25596 19488
rect 25648 19479 25650 19488
rect 25778 19544 25834 19553
rect 25778 19479 25834 19488
rect 25596 19450 25648 19456
rect 25688 19440 25740 19446
rect 25688 19382 25740 19388
rect 25504 17876 25556 17882
rect 25504 17818 25556 17824
rect 25596 17808 25648 17814
rect 25596 17750 25648 17756
rect 25504 17740 25556 17746
rect 25504 17682 25556 17688
rect 25516 16969 25544 17682
rect 25608 17066 25636 17750
rect 25596 17060 25648 17066
rect 25596 17002 25648 17008
rect 25502 16960 25558 16969
rect 25502 16895 25558 16904
rect 25608 16726 25636 17002
rect 25596 16720 25648 16726
rect 25596 16662 25648 16668
rect 25700 16561 25728 19382
rect 25778 18456 25834 18465
rect 25778 18391 25780 18400
rect 25832 18391 25834 18400
rect 25780 18362 25832 18368
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25792 17746 25820 18158
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25780 17604 25832 17610
rect 25780 17546 25832 17552
rect 25792 16658 25820 17546
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25228 16526 25280 16532
rect 25410 16552 25466 16561
rect 25320 16516 25372 16522
rect 25410 16487 25466 16496
rect 25686 16552 25742 16561
rect 25686 16487 25742 16496
rect 25320 16458 25372 16464
rect 25228 15088 25280 15094
rect 25228 15030 25280 15036
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25134 12200 25190 12209
rect 25134 12135 25190 12144
rect 25148 11898 25176 12135
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 24964 11614 25084 11642
rect 24872 10526 24992 10554
rect 24400 10260 24452 10266
rect 24400 10202 24452 10208
rect 24320 10118 24440 10146
rect 23996 9820 24304 9829
rect 23996 9818 24002 9820
rect 24058 9818 24082 9820
rect 24138 9818 24162 9820
rect 24218 9818 24242 9820
rect 24298 9818 24304 9820
rect 24058 9766 24060 9818
rect 24240 9766 24242 9818
rect 23996 9764 24002 9766
rect 24058 9764 24082 9766
rect 24138 9764 24162 9766
rect 24218 9764 24242 9766
rect 24298 9764 24304 9766
rect 23996 9755 24304 9764
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23996 8732 24304 8741
rect 23996 8730 24002 8732
rect 24058 8730 24082 8732
rect 24138 8730 24162 8732
rect 24218 8730 24242 8732
rect 24298 8730 24304 8732
rect 24058 8678 24060 8730
rect 24240 8678 24242 8730
rect 23996 8676 24002 8678
rect 24058 8676 24082 8678
rect 24138 8676 24162 8678
rect 24218 8676 24242 8678
rect 24298 8676 24304 8678
rect 23996 8667 24304 8676
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22560 8424 22612 8430
rect 14280 8366 14332 8372
rect 19522 8392 19578 8401
rect 22560 8366 22612 8372
rect 19522 8327 19578 8336
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 12473 8188 12781 8197
rect 12473 8186 12479 8188
rect 12535 8186 12559 8188
rect 12615 8186 12639 8188
rect 12695 8186 12719 8188
rect 12775 8186 12781 8188
rect 12535 8134 12537 8186
rect 12717 8134 12719 8186
rect 12473 8132 12479 8134
rect 12535 8132 12559 8134
rect 12615 8132 12639 8134
rect 12695 8132 12719 8134
rect 12775 8132 12781 8134
rect 12473 8123 12781 8132
rect 20155 8188 20463 8197
rect 20155 8186 20161 8188
rect 20217 8186 20241 8188
rect 20297 8186 20321 8188
rect 20377 8186 20401 8188
rect 20457 8186 20463 8188
rect 20217 8134 20219 8186
rect 20399 8134 20401 8186
rect 20155 8132 20161 8134
rect 20217 8132 20241 8134
rect 20297 8132 20321 8134
rect 20377 8132 20401 8134
rect 20457 8132 20463 8134
rect 20155 8123 20463 8132
rect 21376 7954 21404 8230
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 16314 7644 16622 7653
rect 16314 7642 16320 7644
rect 16376 7642 16400 7644
rect 16456 7642 16480 7644
rect 16536 7642 16560 7644
rect 16616 7642 16622 7644
rect 16376 7590 16378 7642
rect 16558 7590 16560 7642
rect 16314 7588 16320 7590
rect 16376 7588 16400 7590
rect 16456 7588 16480 7590
rect 16536 7588 16560 7590
rect 16616 7588 16622 7590
rect 16314 7579 16622 7588
rect 23996 7644 24304 7653
rect 23996 7642 24002 7644
rect 24058 7642 24082 7644
rect 24138 7642 24162 7644
rect 24218 7642 24242 7644
rect 24298 7642 24304 7644
rect 24058 7590 24060 7642
rect 24240 7590 24242 7642
rect 23996 7588 24002 7590
rect 24058 7588 24082 7590
rect 24138 7588 24162 7590
rect 24218 7588 24242 7590
rect 24298 7588 24304 7590
rect 23996 7579 24304 7588
rect 12473 7100 12781 7109
rect 12473 7098 12479 7100
rect 12535 7098 12559 7100
rect 12615 7098 12639 7100
rect 12695 7098 12719 7100
rect 12775 7098 12781 7100
rect 12535 7046 12537 7098
rect 12717 7046 12719 7098
rect 12473 7044 12479 7046
rect 12535 7044 12559 7046
rect 12615 7044 12639 7046
rect 12695 7044 12719 7046
rect 12775 7044 12781 7046
rect 12473 7035 12781 7044
rect 20155 7100 20463 7109
rect 20155 7098 20161 7100
rect 20217 7098 20241 7100
rect 20297 7098 20321 7100
rect 20377 7098 20401 7100
rect 20457 7098 20463 7100
rect 20217 7046 20219 7098
rect 20399 7046 20401 7098
rect 20155 7044 20161 7046
rect 20217 7044 20241 7046
rect 20297 7044 20321 7046
rect 20377 7044 20401 7046
rect 20457 7044 20463 7046
rect 20155 7035 20463 7044
rect 12084 6886 12204 6914
rect 8632 6556 8940 6565
rect 8632 6554 8638 6556
rect 8694 6554 8718 6556
rect 8774 6554 8798 6556
rect 8854 6554 8878 6556
rect 8934 6554 8940 6556
rect 8694 6502 8696 6554
rect 8876 6502 8878 6554
rect 8632 6500 8638 6502
rect 8694 6500 8718 6502
rect 8774 6500 8798 6502
rect 8854 6500 8878 6502
rect 8934 6500 8940 6502
rect 8632 6491 8940 6500
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8632 5468 8940 5477
rect 8632 5466 8638 5468
rect 8694 5466 8718 5468
rect 8774 5466 8798 5468
rect 8854 5466 8878 5468
rect 8934 5466 8940 5468
rect 8694 5414 8696 5466
rect 8876 5414 8878 5466
rect 8632 5412 8638 5414
rect 8694 5412 8718 5414
rect 8774 5412 8798 5414
rect 8854 5412 8878 5414
rect 8934 5412 8940 5414
rect 8632 5403 8940 5412
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 12176 5302 12204 6886
rect 16314 6556 16622 6565
rect 16314 6554 16320 6556
rect 16376 6554 16400 6556
rect 16456 6554 16480 6556
rect 16536 6554 16560 6556
rect 16616 6554 16622 6556
rect 16376 6502 16378 6554
rect 16558 6502 16560 6554
rect 16314 6500 16320 6502
rect 16376 6500 16400 6502
rect 16456 6500 16480 6502
rect 16536 6500 16560 6502
rect 16616 6500 16622 6502
rect 16314 6491 16622 6500
rect 23996 6556 24304 6565
rect 23996 6554 24002 6556
rect 24058 6554 24082 6556
rect 24138 6554 24162 6556
rect 24218 6554 24242 6556
rect 24298 6554 24304 6556
rect 24058 6502 24060 6554
rect 24240 6502 24242 6554
rect 23996 6500 24002 6502
rect 24058 6500 24082 6502
rect 24138 6500 24162 6502
rect 24218 6500 24242 6502
rect 24298 6500 24304 6502
rect 23996 6491 24304 6500
rect 12473 6012 12781 6021
rect 12473 6010 12479 6012
rect 12535 6010 12559 6012
rect 12615 6010 12639 6012
rect 12695 6010 12719 6012
rect 12775 6010 12781 6012
rect 12535 5958 12537 6010
rect 12717 5958 12719 6010
rect 12473 5956 12479 5958
rect 12535 5956 12559 5958
rect 12615 5956 12639 5958
rect 12695 5956 12719 5958
rect 12775 5956 12781 5958
rect 12473 5947 12781 5956
rect 20155 6012 20463 6021
rect 20155 6010 20161 6012
rect 20217 6010 20241 6012
rect 20297 6010 20321 6012
rect 20377 6010 20401 6012
rect 20457 6010 20463 6012
rect 20217 5958 20219 6010
rect 20399 5958 20401 6010
rect 20155 5956 20161 5958
rect 20217 5956 20241 5958
rect 20297 5956 20321 5958
rect 20377 5956 20401 5958
rect 20457 5956 20463 5958
rect 20155 5947 20463 5956
rect 16314 5468 16622 5477
rect 16314 5466 16320 5468
rect 16376 5466 16400 5468
rect 16456 5466 16480 5468
rect 16536 5466 16560 5468
rect 16616 5466 16622 5468
rect 16376 5414 16378 5466
rect 16558 5414 16560 5466
rect 16314 5412 16320 5414
rect 16376 5412 16400 5414
rect 16456 5412 16480 5414
rect 16536 5412 16560 5414
rect 16616 5412 16622 5414
rect 16314 5403 16622 5412
rect 23996 5468 24304 5477
rect 23996 5466 24002 5468
rect 24058 5466 24082 5468
rect 24138 5466 24162 5468
rect 24218 5466 24242 5468
rect 24298 5466 24304 5468
rect 24058 5414 24060 5466
rect 24240 5414 24242 5466
rect 23996 5412 24002 5414
rect 24058 5412 24082 5414
rect 24138 5412 24162 5414
rect 24218 5412 24242 5414
rect 24298 5412 24304 5414
rect 23996 5403 24304 5412
rect 12164 5296 12216 5302
rect 5170 5264 5226 5273
rect 12164 5238 12216 5244
rect 24412 5234 24440 10118
rect 24964 9518 24992 10526
rect 24952 9512 25004 9518
rect 25056 9489 25084 11614
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 25148 10470 25176 10610
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25148 10305 25176 10406
rect 25134 10296 25190 10305
rect 25134 10231 25190 10240
rect 25240 10198 25268 15030
rect 25332 12646 25360 16458
rect 25410 16416 25466 16425
rect 25410 16351 25466 16360
rect 25424 14940 25452 16351
rect 25594 16008 25650 16017
rect 25594 15943 25650 15952
rect 25608 15910 25636 15943
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 25504 14952 25556 14958
rect 25424 14912 25504 14940
rect 25504 14894 25556 14900
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25502 14648 25558 14657
rect 25412 14612 25464 14618
rect 25700 14634 25728 14894
rect 25502 14583 25558 14592
rect 25608 14606 25728 14634
rect 25412 14554 25464 14560
rect 25424 13938 25452 14554
rect 25516 14550 25544 14583
rect 25504 14544 25556 14550
rect 25504 14486 25556 14492
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25424 13569 25452 13670
rect 25410 13560 25466 13569
rect 25410 13495 25466 13504
rect 25516 13258 25544 13874
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 25502 13152 25558 13161
rect 25424 12850 25452 13126
rect 25502 13087 25558 13096
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25424 12753 25452 12786
rect 25410 12744 25466 12753
rect 25410 12679 25466 12688
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25320 12368 25372 12374
rect 25320 12310 25372 12316
rect 25228 10192 25280 10198
rect 25228 10134 25280 10140
rect 25228 9512 25280 9518
rect 24952 9454 25004 9460
rect 25042 9480 25098 9489
rect 24964 8242 24992 9454
rect 25228 9454 25280 9460
rect 25042 9415 25098 9424
rect 25240 8945 25268 9454
rect 25332 9110 25360 12310
rect 25424 9738 25452 12679
rect 25516 12170 25544 13087
rect 25504 12164 25556 12170
rect 25504 12106 25556 12112
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25516 10266 25544 10950
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25424 9722 25544 9738
rect 25424 9716 25556 9722
rect 25424 9710 25504 9716
rect 25504 9658 25556 9664
rect 25412 9648 25464 9654
rect 25410 9616 25412 9625
rect 25464 9616 25466 9625
rect 25410 9551 25466 9560
rect 25320 9104 25372 9110
rect 25424 9081 25452 9551
rect 25320 9046 25372 9052
rect 25410 9072 25466 9081
rect 25410 9007 25466 9016
rect 25226 8936 25282 8945
rect 25226 8871 25282 8880
rect 25240 8838 25268 8871
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 24872 8214 24992 8242
rect 24872 7750 24900 8214
rect 25240 8090 25268 8774
rect 25516 8634 25544 9658
rect 25608 9450 25636 14606
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25700 13977 25728 14214
rect 25686 13968 25742 13977
rect 25686 13903 25742 13912
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25700 13297 25728 13670
rect 25686 13288 25742 13297
rect 25686 13223 25742 13232
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25596 9444 25648 9450
rect 25596 9386 25648 9392
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24872 7410 24900 7686
rect 25700 7546 25728 12922
rect 25792 11014 25820 16594
rect 25884 12986 25912 19722
rect 25976 18630 26004 20742
rect 26238 20703 26294 20712
rect 26148 20528 26200 20534
rect 26068 20488 26148 20516
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 26068 18442 26096 20488
rect 26148 20470 26200 20476
rect 26344 20244 26372 21558
rect 26422 21312 26478 21321
rect 26422 21247 26478 21256
rect 26436 20777 26464 21247
rect 26422 20768 26478 20777
rect 26422 20703 26478 20712
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26436 20369 26464 20538
rect 26422 20360 26478 20369
rect 26422 20295 26478 20304
rect 26160 20216 26372 20244
rect 26160 20097 26188 20216
rect 26146 20088 26202 20097
rect 26528 20058 26556 22578
rect 26620 22545 26648 23718
rect 26896 23769 26924 23802
rect 26792 23734 26844 23740
rect 26882 23760 26938 23769
rect 26698 23695 26754 23704
rect 26988 23730 27016 23990
rect 26882 23695 26938 23704
rect 26976 23724 27028 23730
rect 26712 23662 26740 23695
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26712 23118 26740 23598
rect 26792 23316 26844 23322
rect 26792 23258 26844 23264
rect 26700 23112 26752 23118
rect 26700 23054 26752 23060
rect 26606 22536 26662 22545
rect 26606 22471 26662 22480
rect 26700 22432 26752 22438
rect 26700 22374 26752 22380
rect 26712 22234 26740 22374
rect 26700 22228 26752 22234
rect 26700 22170 26752 22176
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 26620 21554 26648 22102
rect 26700 22092 26752 22098
rect 26700 22034 26752 22040
rect 26712 21622 26740 22034
rect 26804 21622 26832 23258
rect 26700 21616 26752 21622
rect 26700 21558 26752 21564
rect 26792 21616 26844 21622
rect 26792 21558 26844 21564
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26620 20874 26648 21490
rect 26698 21040 26754 21049
rect 26698 20975 26754 20984
rect 26712 20942 26740 20975
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 26608 20868 26660 20874
rect 26608 20810 26660 20816
rect 26620 20398 26648 20810
rect 26712 20466 26740 20878
rect 26896 20714 26924 23695
rect 26976 23666 27028 23672
rect 26976 23248 27028 23254
rect 27080 23236 27108 24754
rect 27172 23712 27200 24908
rect 27228 24880 27280 24886
rect 27280 24828 27292 24868
rect 27228 24822 27292 24828
rect 27264 24614 27292 24822
rect 27252 24608 27304 24614
rect 27252 24550 27304 24556
rect 27250 24032 27306 24041
rect 27250 23967 27306 23976
rect 27264 23866 27292 23967
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27356 23780 27384 25724
rect 27620 25774 27672 25780
rect 27712 25832 27764 25838
rect 27712 25774 27764 25780
rect 27526 25735 27582 25744
rect 27436 25706 27488 25712
rect 27434 25664 27490 25673
rect 27724 25650 27752 25774
rect 27816 25770 27844 26540
rect 28276 26518 28304 26710
rect 28354 26616 28410 26625
rect 28354 26551 28410 26560
rect 28264 26512 28316 26518
rect 28264 26454 28316 26460
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 27896 26376 27948 26382
rect 27894 26344 27896 26353
rect 27948 26344 27950 26353
rect 27894 26279 27950 26288
rect 27988 26308 28040 26314
rect 27988 26250 28040 26256
rect 28000 26024 28028 26250
rect 28092 26194 28120 26386
rect 28172 26376 28224 26382
rect 28368 26364 28396 26551
rect 28224 26336 28396 26364
rect 28172 26318 28224 26324
rect 28092 26166 28396 26194
rect 28000 25996 28304 26024
rect 28170 25936 28226 25945
rect 28170 25871 28226 25880
rect 27804 25764 27856 25770
rect 27804 25706 27856 25712
rect 27490 25622 27752 25650
rect 27434 25599 27490 25608
rect 27837 25596 28145 25605
rect 27837 25594 27843 25596
rect 27899 25594 27923 25596
rect 27979 25594 28003 25596
rect 28059 25594 28083 25596
rect 28139 25594 28145 25596
rect 27899 25542 27901 25594
rect 28081 25542 28083 25594
rect 27837 25540 27843 25542
rect 27899 25540 27923 25542
rect 27979 25540 28003 25542
rect 28059 25540 28083 25542
rect 28139 25540 28145 25542
rect 27434 25528 27490 25537
rect 27434 25463 27490 25472
rect 27618 25528 27674 25537
rect 27837 25531 28145 25540
rect 27618 25463 27674 25472
rect 27988 25492 28040 25498
rect 27448 25140 27476 25463
rect 27632 25412 27660 25463
rect 27988 25434 28040 25440
rect 27632 25384 27752 25412
rect 27724 25294 27752 25384
rect 27804 25356 27856 25362
rect 27804 25298 27856 25304
rect 27712 25288 27764 25294
rect 27712 25230 27764 25236
rect 27448 25112 27752 25140
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27434 24848 27490 24857
rect 27632 24834 27660 24890
rect 27490 24806 27660 24834
rect 27724 24818 27752 25112
rect 27712 24812 27764 24818
rect 27434 24783 27490 24792
rect 27712 24754 27764 24760
rect 27816 24698 27844 25298
rect 28000 24750 28028 25434
rect 28184 25294 28212 25871
rect 28276 25537 28304 25996
rect 28368 25770 28396 26166
rect 28356 25764 28408 25770
rect 28356 25706 28408 25712
rect 28262 25528 28318 25537
rect 28262 25463 28318 25472
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28264 25220 28316 25226
rect 28264 25162 28316 25168
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 27632 24670 27844 24698
rect 27988 24744 28040 24750
rect 27988 24686 28040 24692
rect 27528 24608 27580 24614
rect 27528 24550 27580 24556
rect 27540 23866 27568 24550
rect 27632 24410 27660 24670
rect 27712 24608 27764 24614
rect 27712 24550 27764 24556
rect 27620 24404 27672 24410
rect 27620 24346 27672 24352
rect 27724 24154 27752 24550
rect 27837 24508 28145 24517
rect 27837 24506 27843 24508
rect 27899 24506 27923 24508
rect 27979 24506 28003 24508
rect 28059 24506 28083 24508
rect 28139 24506 28145 24508
rect 27899 24454 27901 24506
rect 28081 24454 28083 24506
rect 27837 24452 27843 24454
rect 27899 24452 27923 24454
rect 27979 24452 28003 24454
rect 28059 24452 28083 24454
rect 28139 24452 28145 24454
rect 27837 24443 28145 24452
rect 28184 24290 28212 24754
rect 28276 24410 28304 25162
rect 28460 24818 28488 27814
rect 28552 26994 28580 27934
rect 28630 27840 28686 27849
rect 28630 27775 28686 27784
rect 28540 26988 28592 26994
rect 28540 26930 28592 26936
rect 28538 26480 28594 26489
rect 28538 26415 28594 26424
rect 28448 24812 28500 24818
rect 28368 24772 28448 24800
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28184 24262 28304 24290
rect 27724 24126 28120 24154
rect 27804 24064 27856 24070
rect 27724 24024 27804 24052
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 27356 23752 27476 23780
rect 27172 23684 27384 23712
rect 27158 23624 27214 23633
rect 27158 23559 27214 23568
rect 27028 23208 27108 23236
rect 26976 23190 27028 23196
rect 26988 22642 27016 23190
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 27172 23066 27200 23559
rect 27356 23168 27384 23684
rect 27448 23497 27476 23752
rect 27724 23730 27752 24024
rect 27804 24006 27856 24012
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 28000 23508 28028 23666
rect 27434 23488 27490 23497
rect 27434 23423 27490 23432
rect 27632 23480 28028 23508
rect 28092 23508 28120 24126
rect 28092 23480 28212 23508
rect 27356 23140 27568 23168
rect 27080 22982 27108 23054
rect 27172 23038 27384 23066
rect 27068 22976 27120 22982
rect 27252 22976 27304 22982
rect 27068 22918 27120 22924
rect 27158 22944 27214 22953
rect 27252 22918 27304 22924
rect 27158 22879 27214 22888
rect 27172 22760 27200 22879
rect 27080 22732 27200 22760
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 26988 22137 27016 22170
rect 26974 22128 27030 22137
rect 26974 22063 27030 22072
rect 26974 21720 27030 21729
rect 26974 21655 27030 21664
rect 26988 21622 27016 21655
rect 26976 21616 27028 21622
rect 26976 21558 27028 21564
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 26988 21350 27016 21422
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26788 20686 26924 20714
rect 26700 20460 26752 20466
rect 26788 20448 26816 20686
rect 26976 20460 27028 20466
rect 26788 20420 26832 20448
rect 26700 20402 26752 20408
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26698 20360 26754 20369
rect 26146 20023 26202 20032
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26148 19984 26200 19990
rect 26148 19926 26200 19932
rect 26160 18698 26188 19926
rect 26424 19916 26476 19922
rect 26424 19858 26476 19864
rect 26332 19440 26384 19446
rect 26332 19382 26384 19388
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 25976 18414 26096 18442
rect 25976 18222 26004 18414
rect 26252 18358 26280 19110
rect 26344 18970 26372 19382
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 26436 18884 26464 19858
rect 26516 19780 26568 19786
rect 26516 19722 26568 19728
rect 26528 19009 26556 19722
rect 26620 19514 26648 20334
rect 26698 20295 26754 20304
rect 26712 19514 26740 20295
rect 26804 20058 26832 20420
rect 26976 20402 27028 20408
rect 26882 20360 26938 20369
rect 26882 20295 26938 20304
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26896 19922 26924 20295
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26882 19816 26938 19825
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 26514 19000 26570 19009
rect 26514 18935 26570 18944
rect 26436 18856 26556 18884
rect 26332 18828 26384 18834
rect 26332 18770 26384 18776
rect 26344 18680 26372 18770
rect 26528 18714 26556 18856
rect 26620 18834 26648 19450
rect 26700 19236 26752 19242
rect 26700 19178 26752 19184
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26712 18737 26740 19178
rect 26804 18834 26832 19790
rect 26882 19751 26938 19760
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 26698 18728 26754 18737
rect 26528 18686 26648 18714
rect 26344 18652 26464 18680
rect 26148 18352 26200 18358
rect 26148 18294 26200 18300
rect 26240 18352 26292 18358
rect 26240 18294 26292 18300
rect 25964 18216 26016 18222
rect 25962 18184 25964 18193
rect 26016 18184 26018 18193
rect 25962 18119 26018 18128
rect 26160 17746 26188 18294
rect 26252 17785 26280 18294
rect 26330 18184 26386 18193
rect 26330 18119 26386 18128
rect 26238 17776 26294 17785
rect 26148 17740 26200 17746
rect 26238 17711 26294 17720
rect 26148 17682 26200 17688
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25976 16590 26004 17478
rect 26068 17134 26096 17614
rect 26148 17604 26200 17610
rect 26148 17546 26200 17552
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 26068 16658 26096 17070
rect 26160 16658 26188 17546
rect 26252 17241 26280 17546
rect 26238 17232 26294 17241
rect 26238 17167 26294 17176
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 25976 15706 26004 16526
rect 26068 16250 26096 16594
rect 26056 16244 26108 16250
rect 26056 16186 26108 16192
rect 26160 16182 26188 16594
rect 26148 16176 26200 16182
rect 26148 16118 26200 16124
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 26054 15464 26110 15473
rect 26054 15399 26110 15408
rect 25962 15328 26018 15337
rect 25962 15263 26018 15272
rect 25976 15094 26004 15263
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 25964 14952 26016 14958
rect 26068 14929 26096 15399
rect 26160 15366 26188 16118
rect 26252 15910 26280 17167
rect 26344 16726 26372 18119
rect 26436 16794 26464 18652
rect 26620 18340 26648 18686
rect 26698 18663 26754 18672
rect 26792 18624 26844 18630
rect 26896 18612 26924 19751
rect 26988 19378 27016 20402
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 26988 19145 27016 19314
rect 26974 19136 27030 19145
rect 26974 19071 27030 19080
rect 26976 18964 27028 18970
rect 26976 18906 27028 18912
rect 26988 18698 27016 18906
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26844 18584 26924 18612
rect 26792 18566 26844 18572
rect 26700 18352 26752 18358
rect 26514 18320 26570 18329
rect 26620 18312 26700 18340
rect 26700 18294 26752 18300
rect 26514 18255 26570 18264
rect 26528 18154 26556 18255
rect 26804 18204 26832 18566
rect 26884 18420 26936 18426
rect 26884 18362 26936 18368
rect 26896 18329 26924 18362
rect 26882 18320 26938 18329
rect 26882 18255 26938 18264
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26620 18176 26832 18204
rect 26988 18193 27016 18226
rect 26974 18184 27030 18193
rect 26516 18148 26568 18154
rect 26516 18090 26568 18096
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26528 17270 26556 17682
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 26516 17060 26568 17066
rect 26516 17002 26568 17008
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26332 16720 26384 16726
rect 26332 16662 26384 16668
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26344 15722 26372 16662
rect 26252 15694 26372 15722
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 26252 15178 26280 15694
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26160 15150 26280 15178
rect 25964 14894 26016 14900
rect 26054 14920 26110 14929
rect 25976 13841 26004 14894
rect 26054 14855 26110 14864
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 26068 14521 26096 14758
rect 26054 14512 26110 14521
rect 26054 14447 26110 14456
rect 26068 14414 26096 14447
rect 26056 14408 26108 14414
rect 26056 14350 26108 14356
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 25962 13832 26018 13841
rect 25962 13767 26018 13776
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25976 13326 26004 13670
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25872 12368 25924 12374
rect 25870 12336 25872 12345
rect 25924 12336 25926 12345
rect 25870 12271 25926 12280
rect 26068 12238 26096 14214
rect 26160 13938 26188 15150
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 26252 14464 26280 15030
rect 26344 14657 26372 15302
rect 26330 14648 26386 14657
rect 26330 14583 26386 14592
rect 26252 14436 26372 14464
rect 26238 13968 26294 13977
rect 26148 13932 26200 13938
rect 26238 13903 26294 13912
rect 26148 13874 26200 13880
rect 26252 13802 26280 13903
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26344 13433 26372 14436
rect 26436 14006 26464 16730
rect 26528 16697 26556 17002
rect 26514 16688 26570 16697
rect 26514 16623 26570 16632
rect 26620 16590 26648 18176
rect 26974 18119 27030 18128
rect 26804 18006 27016 18034
rect 26698 17912 26754 17921
rect 26698 17847 26754 17856
rect 26712 17542 26740 17847
rect 26804 17610 26832 18006
rect 26988 17921 27016 18006
rect 26974 17912 27030 17921
rect 26884 17876 26936 17882
rect 26974 17847 27030 17856
rect 26884 17818 26936 17824
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26790 17504 26846 17513
rect 26790 17439 26846 17448
rect 26700 17264 26752 17270
rect 26700 17206 26752 17212
rect 26712 17134 26740 17206
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 26698 16960 26754 16969
rect 26698 16895 26754 16904
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26712 16153 26740 16895
rect 26698 16144 26754 16153
rect 26516 16108 26568 16114
rect 26698 16079 26754 16088
rect 26516 16050 26568 16056
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26330 13424 26386 13433
rect 26330 13359 26386 13368
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 26160 12084 26188 13194
rect 26240 12844 26292 12850
rect 26528 12832 26556 16050
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 26620 13977 26648 15982
rect 26606 13968 26662 13977
rect 26712 13938 26740 16079
rect 26804 16017 26832 17439
rect 26896 17241 26924 17818
rect 26974 17640 27030 17649
rect 26974 17575 26976 17584
rect 27028 17575 27030 17584
rect 26976 17546 27028 17552
rect 26882 17232 26938 17241
rect 26882 17167 26938 17176
rect 26988 16833 27016 17546
rect 26974 16824 27030 16833
rect 26884 16788 26936 16794
rect 26974 16759 27030 16768
rect 26884 16730 26936 16736
rect 26896 16640 26924 16730
rect 26976 16652 27028 16658
rect 26896 16612 26976 16640
rect 26976 16594 27028 16600
rect 26884 16448 26936 16454
rect 26882 16416 26884 16425
rect 26936 16416 26938 16425
rect 26882 16351 26938 16360
rect 26790 16008 26846 16017
rect 26790 15943 26846 15952
rect 26804 15570 26832 15943
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26884 15496 26936 15502
rect 26882 15464 26884 15473
rect 26936 15464 26938 15473
rect 26882 15399 26938 15408
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26804 14618 26832 15302
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26896 14550 26924 14826
rect 26884 14544 26936 14550
rect 26884 14486 26936 14492
rect 26896 14346 26924 14486
rect 26988 14482 27016 16594
rect 27080 16454 27108 22732
rect 27264 22642 27292 22918
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27250 22536 27306 22545
rect 27250 22471 27306 22480
rect 27264 22438 27292 22471
rect 27252 22432 27304 22438
rect 27252 22374 27304 22380
rect 27264 22094 27292 22374
rect 27172 22066 27292 22094
rect 27356 22080 27384 23038
rect 27540 22964 27568 23140
rect 27632 23118 27660 23480
rect 27837 23420 28145 23429
rect 27837 23418 27843 23420
rect 27899 23418 27923 23420
rect 27979 23418 28003 23420
rect 28059 23418 28083 23420
rect 28139 23418 28145 23420
rect 27899 23366 27901 23418
rect 28081 23366 28083 23418
rect 27837 23364 27843 23366
rect 27899 23364 27923 23366
rect 27979 23364 28003 23366
rect 28059 23364 28083 23366
rect 28139 23364 28145 23366
rect 27710 23352 27766 23361
rect 27837 23355 28145 23364
rect 27710 23287 27712 23296
rect 27764 23287 27766 23296
rect 27712 23258 27764 23264
rect 27804 23248 27856 23254
rect 27804 23190 27856 23196
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27724 22964 27752 23054
rect 27540 22936 27752 22964
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27526 22536 27582 22545
rect 27526 22471 27582 22480
rect 27540 22438 27568 22471
rect 27528 22432 27580 22438
rect 27632 22409 27660 22578
rect 27816 22420 27844 23190
rect 28078 22808 28134 22817
rect 28078 22743 28134 22752
rect 28092 22574 28120 22743
rect 28080 22568 28132 22574
rect 28080 22510 28132 22516
rect 27528 22374 27580 22380
rect 27618 22400 27674 22409
rect 27618 22335 27674 22344
rect 27724 22392 27844 22420
rect 27528 22092 27580 22098
rect 27172 21894 27200 22066
rect 27356 22052 27476 22080
rect 27252 22024 27304 22030
rect 27252 21966 27304 21972
rect 27448 21978 27476 22052
rect 27724 22080 27752 22392
rect 28184 22386 28212 23480
rect 28276 22817 28304 24262
rect 28368 23730 28396 24772
rect 28448 24754 28500 24760
rect 28448 24608 28500 24614
rect 28448 24550 28500 24556
rect 28460 23798 28488 24550
rect 28552 24138 28580 26415
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28448 23792 28500 23798
rect 28448 23734 28500 23740
rect 28356 23724 28408 23730
rect 28356 23666 28408 23672
rect 28460 23361 28488 23734
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28552 23594 28580 23666
rect 28540 23588 28592 23594
rect 28540 23530 28592 23536
rect 28538 23488 28594 23497
rect 28538 23423 28594 23432
rect 28446 23352 28502 23361
rect 28552 23322 28580 23423
rect 28446 23287 28502 23296
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28644 23202 28672 27775
rect 28736 27538 28764 30874
rect 28828 29730 28856 30874
rect 28908 30660 28960 30666
rect 28908 30602 28960 30608
rect 28920 30258 28948 30602
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 28828 29702 28948 29730
rect 28816 29640 28868 29646
rect 28816 29582 28868 29588
rect 28828 29073 28856 29582
rect 28920 29152 28948 29702
rect 29012 29646 29040 30534
rect 29000 29640 29052 29646
rect 29000 29582 29052 29588
rect 29000 29504 29052 29510
rect 29000 29446 29052 29452
rect 29012 29345 29040 29446
rect 28998 29336 29054 29345
rect 28998 29271 29054 29280
rect 28920 29124 29040 29152
rect 28814 29064 28870 29073
rect 28814 28999 28870 29008
rect 28908 29028 28960 29034
rect 28908 28970 28960 28976
rect 28816 28960 28868 28966
rect 28920 28937 28948 28970
rect 28816 28902 28868 28908
rect 28906 28928 28962 28937
rect 28828 28150 28856 28902
rect 28906 28863 28962 28872
rect 28906 28656 28962 28665
rect 28906 28591 28962 28600
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 28816 28008 28868 28014
rect 28816 27950 28868 27956
rect 28828 27538 28856 27950
rect 28724 27532 28776 27538
rect 28724 27474 28776 27480
rect 28816 27532 28868 27538
rect 28816 27474 28868 27480
rect 28736 27418 28764 27474
rect 28920 27418 28948 28591
rect 29012 28422 29040 29124
rect 29104 28626 29132 34303
rect 29656 32434 29684 34350
rect 30378 33960 30434 33969
rect 30378 33895 30434 33904
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 30288 32224 30340 32230
rect 30288 32166 30340 32172
rect 29276 31952 29328 31958
rect 29276 31894 29328 31900
rect 29642 31920 29698 31929
rect 29184 29844 29236 29850
rect 29184 29786 29236 29792
rect 29196 28966 29224 29786
rect 29184 28960 29236 28966
rect 29184 28902 29236 28908
rect 29092 28620 29144 28626
rect 29092 28562 29144 28568
rect 29104 28422 29132 28562
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29092 28416 29144 28422
rect 29092 28358 29144 28364
rect 29012 27538 29040 28358
rect 29090 27704 29146 27713
rect 29090 27639 29092 27648
rect 29144 27639 29146 27648
rect 29092 27610 29144 27616
rect 29000 27532 29052 27538
rect 29000 27474 29052 27480
rect 28736 27390 28856 27418
rect 28920 27390 29040 27418
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28736 26874 28764 27270
rect 28828 27062 28856 27390
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28920 27169 28948 27270
rect 28906 27160 28962 27169
rect 28906 27095 28962 27104
rect 28816 27056 28868 27062
rect 28816 26998 28868 27004
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 28736 26846 28856 26874
rect 28724 26784 28776 26790
rect 28828 26761 28856 26846
rect 28724 26726 28776 26732
rect 28814 26752 28870 26761
rect 28736 26602 28764 26726
rect 28814 26687 28870 26696
rect 28736 26574 28856 26602
rect 28920 26586 28948 26930
rect 28828 26466 28856 26574
rect 28908 26580 28960 26586
rect 28908 26522 28960 26528
rect 29012 26518 29040 27390
rect 29092 27396 29144 27402
rect 29092 27338 29144 27344
rect 29000 26512 29052 26518
rect 28906 26480 28962 26489
rect 28828 26438 28906 26466
rect 29104 26489 29132 27338
rect 29000 26454 29052 26460
rect 29090 26480 29146 26489
rect 28906 26415 28962 26424
rect 29090 26415 29146 26424
rect 28724 26376 28776 26382
rect 28722 26344 28724 26353
rect 29000 26376 29052 26382
rect 28776 26344 28778 26353
rect 29092 26376 29144 26382
rect 29000 26318 29052 26324
rect 29090 26344 29092 26353
rect 29144 26344 29146 26353
rect 28722 26279 28778 26288
rect 28908 26036 28960 26042
rect 28908 25978 28960 25984
rect 28816 25900 28868 25906
rect 28816 25842 28868 25848
rect 28828 25294 28856 25842
rect 28816 25288 28868 25294
rect 28816 25230 28868 25236
rect 28816 24948 28868 24954
rect 28816 24890 28868 24896
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28736 24274 28764 24754
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28724 24064 28776 24070
rect 28724 24006 28776 24012
rect 28736 23594 28764 24006
rect 28828 23610 28856 24890
rect 28920 24410 28948 25978
rect 29012 24449 29040 26318
rect 29090 26279 29146 26288
rect 29092 26240 29144 26246
rect 29092 26182 29144 26188
rect 29104 24954 29132 26182
rect 29196 26042 29224 28426
rect 29288 28393 29316 31894
rect 29642 31855 29698 31864
rect 29368 31136 29420 31142
rect 29368 31078 29420 31084
rect 29380 29034 29408 31078
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29472 29170 29500 29990
rect 29460 29164 29512 29170
rect 29460 29106 29512 29112
rect 29368 29028 29420 29034
rect 29368 28970 29420 28976
rect 29274 28384 29330 28393
rect 29274 28319 29330 28328
rect 29276 28144 29328 28150
rect 29276 28086 29328 28092
rect 29288 27849 29316 28086
rect 29274 27840 29330 27849
rect 29274 27775 29330 27784
rect 29274 27704 29330 27713
rect 29274 27639 29330 27648
rect 29288 27062 29316 27639
rect 29276 27056 29328 27062
rect 29276 26998 29328 27004
rect 29380 26994 29408 28970
rect 29458 28656 29514 28665
rect 29458 28591 29514 28600
rect 29472 28558 29500 28591
rect 29460 28552 29512 28558
rect 29460 28494 29512 28500
rect 29460 28416 29512 28422
rect 29460 28358 29512 28364
rect 29472 28150 29500 28358
rect 29460 28144 29512 28150
rect 29460 28086 29512 28092
rect 29472 27985 29500 28086
rect 29564 28082 29592 30126
rect 29552 28076 29604 28082
rect 29552 28018 29604 28024
rect 29458 27976 29514 27985
rect 29458 27911 29514 27920
rect 29460 27872 29512 27878
rect 29460 27814 29512 27820
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29368 26852 29420 26858
rect 29368 26794 29420 26800
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 29288 26081 29316 26726
rect 29380 26586 29408 26794
rect 29368 26580 29420 26586
rect 29368 26522 29420 26528
rect 29368 26376 29420 26382
rect 29368 26318 29420 26324
rect 29274 26072 29330 26081
rect 29184 26036 29236 26042
rect 29274 26007 29330 26016
rect 29184 25978 29236 25984
rect 29380 25956 29408 26318
rect 29182 25936 29238 25945
rect 29182 25871 29238 25880
rect 29288 25928 29408 25956
rect 29196 25838 29224 25871
rect 29184 25832 29236 25838
rect 29184 25774 29236 25780
rect 29196 25650 29224 25774
rect 29288 25770 29316 25928
rect 29366 25800 29422 25809
rect 29276 25764 29328 25770
rect 29366 25735 29422 25744
rect 29276 25706 29328 25712
rect 29196 25622 29316 25650
rect 29184 25220 29236 25226
rect 29184 25162 29236 25168
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29090 24848 29146 24857
rect 29090 24783 29146 24792
rect 28998 24440 29054 24449
rect 28908 24404 28960 24410
rect 28998 24375 29054 24384
rect 28908 24346 28960 24352
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28920 23730 28948 24210
rect 28998 24168 29054 24177
rect 28998 24103 29054 24112
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28724 23588 28776 23594
rect 28828 23582 28948 23610
rect 28724 23530 28776 23536
rect 28722 23488 28778 23497
rect 28722 23423 28778 23432
rect 28552 23174 28672 23202
rect 28262 22808 28318 22817
rect 28262 22743 28318 22752
rect 28264 22636 28316 22642
rect 28448 22636 28500 22642
rect 28316 22596 28396 22624
rect 28264 22578 28316 22584
rect 28368 22409 28396 22596
rect 28448 22578 28500 22584
rect 28460 22545 28488 22578
rect 28446 22536 28502 22545
rect 28446 22471 28502 22480
rect 28354 22400 28410 22409
rect 28184 22358 28304 22386
rect 27837 22332 28145 22341
rect 27837 22330 27843 22332
rect 27899 22330 27923 22332
rect 27979 22330 28003 22332
rect 28059 22330 28083 22332
rect 28139 22330 28145 22332
rect 27899 22278 27901 22330
rect 28081 22278 28083 22330
rect 27837 22276 27843 22278
rect 27899 22276 27923 22278
rect 27979 22276 28003 22278
rect 28059 22276 28083 22278
rect 28139 22276 28145 22278
rect 27837 22267 28145 22276
rect 27580 22052 27752 22080
rect 27908 22052 28212 22080
rect 27528 22034 27580 22040
rect 27908 21978 27936 22052
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27160 21616 27212 21622
rect 27160 21558 27212 21564
rect 27172 20584 27200 21558
rect 27264 21049 27292 21966
rect 27344 21956 27396 21962
rect 27448 21950 27936 21978
rect 27988 22018 28040 22024
rect 27988 21960 28040 21966
rect 28184 21962 28212 22052
rect 27344 21898 27396 21904
rect 27250 21040 27306 21049
rect 27356 21010 27384 21898
rect 27436 21888 27488 21894
rect 28000 21876 28028 21960
rect 28172 21956 28224 21962
rect 28172 21898 28224 21904
rect 27436 21830 27488 21836
rect 27724 21848 28028 21876
rect 27448 21049 27476 21830
rect 27618 21312 27674 21321
rect 27618 21247 27674 21256
rect 27434 21040 27490 21049
rect 27250 20975 27306 20984
rect 27344 21004 27396 21010
rect 27632 21010 27660 21247
rect 27724 21128 27752 21848
rect 28276 21706 28304 22358
rect 28354 22335 28410 22344
rect 28354 22264 28410 22273
rect 28354 22199 28410 22208
rect 28448 22228 28500 22234
rect 28092 21678 28304 21706
rect 28092 21332 28120 21678
rect 28172 21616 28224 21622
rect 28224 21576 28304 21604
rect 28172 21558 28224 21564
rect 28092 21304 28212 21332
rect 27837 21244 28145 21253
rect 27837 21242 27843 21244
rect 27899 21242 27923 21244
rect 27979 21242 28003 21244
rect 28059 21242 28083 21244
rect 28139 21242 28145 21244
rect 27899 21190 27901 21242
rect 28081 21190 28083 21242
rect 27837 21188 27843 21190
rect 27899 21188 27923 21190
rect 27979 21188 28003 21190
rect 28059 21188 28083 21190
rect 28139 21188 28145 21190
rect 27837 21179 28145 21188
rect 27724 21100 27844 21128
rect 27434 20975 27490 20984
rect 27620 21004 27672 21010
rect 27344 20946 27396 20952
rect 27620 20946 27672 20952
rect 27252 20868 27304 20874
rect 27252 20810 27304 20816
rect 27264 20584 27292 20810
rect 27526 20632 27582 20641
rect 27172 20556 27203 20584
rect 27264 20556 27384 20584
rect 27526 20567 27582 20576
rect 27175 20516 27203 20556
rect 27175 20488 27292 20516
rect 27264 20244 27292 20488
rect 27175 20216 27292 20244
rect 27175 20210 27203 20216
rect 27172 20182 27203 20210
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27068 15972 27120 15978
rect 27068 15914 27120 15920
rect 27080 15706 27108 15914
rect 27068 15700 27120 15706
rect 27068 15642 27120 15648
rect 26976 14476 27028 14482
rect 26976 14418 27028 14424
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26884 14340 26936 14346
rect 26884 14282 26936 14288
rect 26804 14249 26832 14282
rect 26790 14240 26846 14249
rect 26790 14175 26846 14184
rect 26606 13903 26662 13912
rect 26700 13932 26752 13938
rect 26292 12804 26556 12832
rect 26240 12786 26292 12792
rect 26068 12056 26188 12084
rect 25872 11756 25924 11762
rect 25872 11698 25924 11704
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25884 10826 25912 11698
rect 25792 10798 25912 10826
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 24950 7440 25006 7449
rect 24860 7404 24912 7410
rect 25792 7426 25820 10798
rect 26068 9518 26096 12056
rect 26146 11928 26202 11937
rect 26146 11863 26148 11872
rect 26200 11863 26202 11872
rect 26148 11834 26200 11840
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 26148 9104 26200 9110
rect 26148 9046 26200 9052
rect 26056 8288 26108 8294
rect 26056 8230 26108 8236
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 24950 7375 25006 7384
rect 25700 7398 25820 7426
rect 24860 7346 24912 7352
rect 24964 7206 24992 7375
rect 25700 7206 25728 7398
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 25688 7200 25740 7206
rect 25688 7142 25740 7148
rect 25700 6662 25728 7142
rect 25884 6934 25912 8026
rect 26068 7478 26096 8230
rect 26056 7472 26108 7478
rect 26056 7414 26108 7420
rect 25872 6928 25924 6934
rect 25872 6870 25924 6876
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25700 6254 25728 6598
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 5170 5199 5226 5208
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 4791 4924 5099 4933
rect 4791 4922 4797 4924
rect 4853 4922 4877 4924
rect 4933 4922 4957 4924
rect 5013 4922 5037 4924
rect 5093 4922 5099 4924
rect 4853 4870 4855 4922
rect 5035 4870 5037 4922
rect 4791 4868 4797 4870
rect 4853 4868 4877 4870
rect 4933 4868 4957 4870
rect 5013 4868 5037 4870
rect 5093 4868 5099 4870
rect 4791 4859 5099 4868
rect 12473 4924 12781 4933
rect 12473 4922 12479 4924
rect 12535 4922 12559 4924
rect 12615 4922 12639 4924
rect 12695 4922 12719 4924
rect 12775 4922 12781 4924
rect 12535 4870 12537 4922
rect 12717 4870 12719 4922
rect 12473 4868 12479 4870
rect 12535 4868 12559 4870
rect 12615 4868 12639 4870
rect 12695 4868 12719 4870
rect 12775 4868 12781 4870
rect 12473 4859 12781 4868
rect 20155 4924 20463 4933
rect 20155 4922 20161 4924
rect 20217 4922 20241 4924
rect 20297 4922 20321 4924
rect 20377 4922 20401 4924
rect 20457 4922 20463 4924
rect 20217 4870 20219 4922
rect 20399 4870 20401 4922
rect 20155 4868 20161 4870
rect 20217 4868 20241 4870
rect 20297 4868 20321 4870
rect 20377 4868 20401 4870
rect 20457 4868 20463 4870
rect 20155 4859 20463 4868
rect 26160 4758 26188 9046
rect 26252 8634 26280 12786
rect 26620 12782 26648 13903
rect 26700 13874 26752 13880
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26608 12776 26660 12782
rect 26608 12718 26660 12724
rect 26712 12434 26740 13874
rect 26896 13841 26924 13874
rect 26882 13832 26938 13841
rect 26792 13796 26844 13802
rect 26882 13767 26938 13776
rect 26792 13738 26844 13744
rect 26804 12850 26832 13738
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26712 12406 26832 12434
rect 26700 12368 26752 12374
rect 26700 12310 26752 12316
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 26344 11762 26372 12174
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 26606 11384 26662 11393
rect 26606 11319 26608 11328
rect 26660 11319 26662 11328
rect 26608 11290 26660 11296
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26344 10674 26372 10950
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26608 10464 26660 10470
rect 26606 10432 26608 10441
rect 26660 10432 26662 10441
rect 26606 10367 26662 10376
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 26436 9761 26464 9862
rect 26422 9752 26478 9761
rect 26422 9687 26478 9696
rect 26608 9580 26660 9586
rect 26608 9522 26660 9528
rect 26424 9376 26476 9382
rect 26422 9344 26424 9353
rect 26476 9344 26478 9353
rect 26422 9279 26478 9288
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26252 8362 26280 8570
rect 26240 8356 26292 8362
rect 26240 8298 26292 8304
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26344 7290 26372 7686
rect 26252 7262 26372 7290
rect 26252 6662 26280 7262
rect 26436 6798 26464 9279
rect 26620 7478 26648 9522
rect 26712 7750 26740 12310
rect 26804 11626 26832 12406
rect 26896 12238 26924 13767
rect 26988 13530 27016 14418
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 26988 12442 27016 12786
rect 27080 12782 27108 15642
rect 27172 14618 27200 20182
rect 27250 20088 27306 20097
rect 27240 20032 27250 20074
rect 27240 20023 27306 20032
rect 27240 19972 27268 20023
rect 27240 19944 27292 19972
rect 27264 19718 27292 19944
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27250 19408 27306 19417
rect 27250 19343 27252 19352
rect 27304 19343 27306 19352
rect 27252 19314 27304 19320
rect 27252 19236 27304 19242
rect 27252 19178 27304 19184
rect 27264 18737 27292 19178
rect 27250 18728 27306 18737
rect 27250 18663 27306 18672
rect 27160 14612 27212 14618
rect 27160 14554 27212 14560
rect 27264 14498 27292 18663
rect 27172 14470 27292 14498
rect 27172 12986 27200 14470
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26974 11928 27030 11937
rect 26974 11863 27030 11872
rect 26792 11620 26844 11626
rect 26792 11562 26844 11568
rect 26804 10130 26832 11562
rect 26884 11348 26936 11354
rect 26884 11290 26936 11296
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26804 8090 26832 10066
rect 26896 9994 26924 11290
rect 26988 10062 27016 11863
rect 27080 11014 27108 12718
rect 27264 12306 27292 13806
rect 27356 13530 27384 20556
rect 27540 20516 27568 20567
rect 27712 20528 27764 20534
rect 27448 20488 27568 20516
rect 27632 20488 27712 20516
rect 27448 20380 27476 20488
rect 27447 20352 27476 20380
rect 27528 20392 27580 20398
rect 27447 20244 27475 20352
rect 27528 20334 27580 20340
rect 27447 20216 27476 20244
rect 27448 20176 27476 20216
rect 27447 20148 27476 20176
rect 27447 20097 27475 20148
rect 27434 20088 27490 20097
rect 27434 20023 27490 20032
rect 27448 19990 27476 20023
rect 27436 19984 27488 19990
rect 27436 19926 27488 19932
rect 27540 19768 27568 20334
rect 27632 19938 27660 20488
rect 27712 20470 27764 20476
rect 27816 20369 27844 21100
rect 27896 20392 27948 20398
rect 27802 20360 27858 20369
rect 27896 20334 27948 20340
rect 27802 20295 27858 20304
rect 27908 20244 27936 20334
rect 27724 20216 27936 20244
rect 27724 20058 27752 20216
rect 27837 20156 28145 20165
rect 27837 20154 27843 20156
rect 27899 20154 27923 20156
rect 27979 20154 28003 20156
rect 28059 20154 28083 20156
rect 28139 20154 28145 20156
rect 27899 20102 27901 20154
rect 28081 20102 28083 20154
rect 27837 20100 27843 20102
rect 27899 20100 27923 20102
rect 27979 20100 28003 20102
rect 28059 20100 28083 20102
rect 28139 20100 28145 20102
rect 27837 20091 28145 20100
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 27632 19922 27752 19938
rect 27632 19916 27764 19922
rect 27632 19910 27712 19916
rect 27712 19858 27764 19864
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27540 19740 27660 19768
rect 27436 19508 27488 19514
rect 27436 19450 27488 19456
rect 27528 19508 27580 19514
rect 27528 19450 27580 19456
rect 27448 19378 27476 19450
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27434 19000 27490 19009
rect 27434 18935 27490 18944
rect 27448 18902 27476 18935
rect 27436 18896 27488 18902
rect 27436 18838 27488 18844
rect 27436 18760 27488 18766
rect 27434 18728 27436 18737
rect 27488 18728 27490 18737
rect 27434 18663 27490 18672
rect 27436 18284 27488 18290
rect 27540 18272 27568 19450
rect 27632 19242 27660 19740
rect 27710 19680 27766 19689
rect 27710 19615 27766 19624
rect 27724 19417 27752 19615
rect 27804 19508 27856 19514
rect 27804 19450 27856 19456
rect 27710 19408 27766 19417
rect 27816 19378 27844 19450
rect 27710 19343 27766 19352
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27908 19310 27936 19790
rect 28184 19496 28212 21304
rect 28276 21185 28304 21576
rect 28262 21176 28318 21185
rect 28262 21111 28318 21120
rect 28262 20088 28318 20097
rect 28262 20023 28318 20032
rect 28276 19718 28304 20023
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 28092 19468 28212 19496
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27620 19236 27672 19242
rect 27620 19178 27672 19184
rect 28092 19156 28120 19468
rect 28172 19372 28224 19378
rect 28224 19332 28304 19360
rect 28172 19314 28224 19320
rect 28172 19236 28224 19242
rect 28172 19178 28224 19184
rect 27724 19128 28120 19156
rect 27724 18970 27752 19128
rect 28184 19122 28212 19178
rect 28276 19145 28304 19332
rect 28368 19174 28396 22199
rect 28448 22170 28500 22176
rect 28460 21418 28488 22170
rect 28552 22098 28580 23174
rect 28736 23100 28764 23423
rect 28814 23352 28870 23361
rect 28814 23287 28816 23296
rect 28868 23287 28870 23296
rect 28816 23258 28868 23264
rect 28644 23089 28764 23100
rect 28816 23112 28868 23118
rect 28630 23080 28764 23089
rect 28686 23072 28764 23080
rect 28814 23080 28816 23089
rect 28868 23080 28870 23089
rect 28630 23015 28686 23024
rect 28814 23015 28870 23024
rect 28724 22500 28776 22506
rect 28920 22488 28948 23582
rect 28776 22460 28948 22488
rect 28724 22442 28776 22448
rect 29012 22438 29040 24103
rect 29104 23866 29132 24783
rect 29196 24342 29224 25162
rect 29288 24818 29316 25622
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29288 24614 29316 24754
rect 29276 24608 29328 24614
rect 29276 24550 29328 24556
rect 29184 24336 29236 24342
rect 29184 24278 29236 24284
rect 29274 24168 29330 24177
rect 29184 24132 29236 24138
rect 29274 24103 29330 24112
rect 29184 24074 29236 24080
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 29090 23488 29146 23497
rect 29090 23423 29146 23432
rect 28632 22432 28684 22438
rect 29000 22432 29052 22438
rect 28684 22380 28856 22386
rect 28632 22374 28856 22380
rect 29000 22374 29052 22380
rect 28644 22358 28856 22374
rect 28632 22228 28684 22234
rect 28632 22170 28684 22176
rect 28644 22098 28672 22170
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 28632 22092 28684 22098
rect 28828 22094 28856 22358
rect 29104 22234 29132 23423
rect 29196 22642 29224 24074
rect 29288 23186 29316 24103
rect 29380 23526 29408 25735
rect 29472 24138 29500 27814
rect 29656 27674 29684 31855
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 29748 31521 29776 31758
rect 29734 31512 29790 31521
rect 29734 31447 29790 31456
rect 29736 30864 29788 30870
rect 29736 30806 29788 30812
rect 29748 30258 29776 30806
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29840 30122 29868 31758
rect 30012 31136 30064 31142
rect 30012 31078 30064 31084
rect 30024 30705 30052 31078
rect 30010 30696 30066 30705
rect 30010 30631 30066 30640
rect 30104 30592 30156 30598
rect 30104 30534 30156 30540
rect 30116 30326 30144 30534
rect 30012 30320 30064 30326
rect 30012 30262 30064 30268
rect 30104 30320 30156 30326
rect 30104 30262 30156 30268
rect 29828 30116 29880 30122
rect 29828 30058 29880 30064
rect 29920 29640 29972 29646
rect 29918 29608 29920 29617
rect 29972 29608 29974 29617
rect 29918 29543 29974 29552
rect 30024 29492 30052 30262
rect 30196 30252 30248 30258
rect 30196 30194 30248 30200
rect 30104 29776 30156 29782
rect 30104 29718 30156 29724
rect 29932 29464 30052 29492
rect 29828 29164 29880 29170
rect 29828 29106 29880 29112
rect 29840 29073 29868 29106
rect 29826 29064 29882 29073
rect 29736 29028 29788 29034
rect 29826 28999 29882 29008
rect 29736 28970 29788 28976
rect 29644 27668 29696 27674
rect 29644 27610 29696 27616
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 29564 27305 29592 27474
rect 29550 27296 29606 27305
rect 29550 27231 29606 27240
rect 29564 26994 29592 27231
rect 29552 26988 29604 26994
rect 29552 26930 29604 26936
rect 29552 26512 29604 26518
rect 29552 26454 29604 26460
rect 29460 24132 29512 24138
rect 29460 24074 29512 24080
rect 29564 23730 29592 26454
rect 29656 25974 29684 27610
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29748 25838 29776 28970
rect 29828 28416 29880 28422
rect 29828 28358 29880 28364
rect 29840 28121 29868 28358
rect 29826 28112 29882 28121
rect 29826 28047 29882 28056
rect 29828 27940 29880 27946
rect 29828 27882 29880 27888
rect 29840 27713 29868 27882
rect 29826 27704 29882 27713
rect 29826 27639 29882 27648
rect 29828 27396 29880 27402
rect 29828 27338 29880 27344
rect 29840 27305 29868 27338
rect 29826 27296 29882 27305
rect 29826 27231 29882 27240
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 29840 26790 29868 27066
rect 29828 26784 29880 26790
rect 29828 26726 29880 26732
rect 29828 26512 29880 26518
rect 29828 26454 29880 26460
rect 29840 26314 29868 26454
rect 29828 26308 29880 26314
rect 29828 26250 29880 26256
rect 29826 26072 29882 26081
rect 29826 26007 29882 26016
rect 29840 25906 29868 26007
rect 29828 25900 29880 25906
rect 29828 25842 29880 25848
rect 29736 25832 29788 25838
rect 29736 25774 29788 25780
rect 29644 25764 29696 25770
rect 29644 25706 29696 25712
rect 29656 25673 29684 25706
rect 29642 25664 29698 25673
rect 29826 25664 29882 25673
rect 29698 25622 29776 25650
rect 29642 25599 29698 25608
rect 29642 25528 29698 25537
rect 29748 25498 29776 25622
rect 29826 25599 29882 25608
rect 29642 25463 29644 25472
rect 29696 25463 29698 25472
rect 29736 25492 29788 25498
rect 29644 25434 29696 25440
rect 29736 25434 29788 25440
rect 29656 24274 29684 25434
rect 29840 25294 29868 25599
rect 29828 25288 29880 25294
rect 29734 25256 29790 25265
rect 29828 25230 29880 25236
rect 29734 25191 29790 25200
rect 29748 25158 29776 25191
rect 29736 25152 29788 25158
rect 29736 25094 29788 25100
rect 29932 24970 29960 29464
rect 30012 29164 30064 29170
rect 30012 29106 30064 29112
rect 30024 28694 30052 29106
rect 30012 28688 30064 28694
rect 30012 28630 30064 28636
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 30024 28393 30052 28494
rect 30010 28384 30066 28393
rect 30010 28319 30066 28328
rect 30116 28082 30144 29718
rect 30208 29306 30236 30194
rect 30196 29300 30248 29306
rect 30196 29242 30248 29248
rect 30196 28960 30248 28966
rect 30196 28902 30248 28908
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 30104 28076 30156 28082
rect 30104 28018 30156 28024
rect 29748 24942 29960 24970
rect 29748 24818 29776 24942
rect 29826 24848 29882 24857
rect 29736 24812 29788 24818
rect 29826 24783 29828 24792
rect 29736 24754 29788 24760
rect 29880 24783 29882 24792
rect 29828 24754 29880 24760
rect 30024 24750 30052 28018
rect 30208 27946 30236 28902
rect 30300 28014 30328 32166
rect 30392 31754 30420 33895
rect 30562 32464 30618 32473
rect 30944 32434 30972 34462
rect 32034 34350 32090 35150
rect 31678 32668 31986 32677
rect 31678 32666 31684 32668
rect 31740 32666 31764 32668
rect 31820 32666 31844 32668
rect 31900 32666 31924 32668
rect 31980 32666 31986 32668
rect 31740 32614 31742 32666
rect 31922 32614 31924 32666
rect 31678 32612 31684 32614
rect 31740 32612 31764 32614
rect 31820 32612 31844 32614
rect 31900 32612 31924 32614
rect 31980 32612 31986 32614
rect 31678 32603 31986 32612
rect 30562 32399 30618 32408
rect 30932 32428 30984 32434
rect 30576 32026 30604 32399
rect 30932 32370 30984 32376
rect 32220 32360 32272 32366
rect 32220 32302 32272 32308
rect 30840 32224 30892 32230
rect 30840 32166 30892 32172
rect 30564 32020 30616 32026
rect 30564 31962 30616 31968
rect 30392 31726 30604 31754
rect 30472 30728 30524 30734
rect 30472 30670 30524 30676
rect 30380 30048 30432 30054
rect 30380 29990 30432 29996
rect 30392 29170 30420 29990
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30378 28520 30434 28529
rect 30378 28455 30434 28464
rect 30392 28422 30420 28455
rect 30380 28416 30432 28422
rect 30380 28358 30432 28364
rect 30288 28008 30340 28014
rect 30288 27950 30340 27956
rect 30196 27940 30248 27946
rect 30196 27882 30248 27888
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30196 27464 30248 27470
rect 30196 27406 30248 27412
rect 30102 27160 30158 27169
rect 30208 27130 30236 27406
rect 30102 27095 30158 27104
rect 30196 27124 30248 27130
rect 30116 27062 30144 27095
rect 30196 27066 30248 27072
rect 30104 27056 30156 27062
rect 30104 26998 30156 27004
rect 30196 26988 30248 26994
rect 30196 26930 30248 26936
rect 30104 26512 30156 26518
rect 30102 26480 30104 26489
rect 30156 26480 30158 26489
rect 30102 26415 30158 26424
rect 30116 25294 30144 26415
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 29736 24676 29788 24682
rect 29736 24618 29788 24624
rect 29644 24268 29696 24274
rect 29644 24210 29696 24216
rect 29748 24070 29776 24618
rect 29920 24336 29972 24342
rect 29826 24304 29882 24313
rect 29920 24278 29972 24284
rect 29826 24239 29882 24248
rect 29840 24206 29868 24239
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 29736 24064 29788 24070
rect 29736 24006 29788 24012
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29644 23860 29696 23866
rect 29644 23802 29696 23808
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29460 23588 29512 23594
rect 29460 23530 29512 23536
rect 29368 23520 29420 23526
rect 29368 23462 29420 23468
rect 29276 23180 29328 23186
rect 29276 23122 29328 23128
rect 29184 22636 29236 22642
rect 29184 22578 29236 22584
rect 29092 22228 29144 22234
rect 29092 22170 29144 22176
rect 28828 22066 28948 22094
rect 28632 22034 28684 22040
rect 28552 21978 28580 22034
rect 28920 22030 28948 22066
rect 28908 22024 28960 22030
rect 28552 21950 28764 21978
rect 28908 21966 28960 21972
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 28448 21412 28500 21418
rect 28448 21354 28500 21360
rect 28630 21176 28686 21185
rect 28630 21111 28686 21120
rect 28540 21004 28592 21010
rect 28460 20964 28540 20992
rect 28460 19514 28488 20964
rect 28540 20946 28592 20952
rect 28540 20868 28592 20874
rect 28540 20810 28592 20816
rect 28552 20584 28580 20810
rect 28644 20806 28672 21111
rect 28632 20800 28684 20806
rect 28632 20742 28684 20748
rect 28552 20556 28672 20584
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28448 19508 28500 19514
rect 28448 19450 28500 19456
rect 28552 19258 28580 20402
rect 28644 20233 28672 20556
rect 28736 20398 28764 21950
rect 28908 21888 28960 21894
rect 29012 21865 29040 21966
rect 29092 21956 29144 21962
rect 29092 21898 29144 21904
rect 28908 21830 28960 21836
rect 28998 21856 29054 21865
rect 28816 21616 28868 21622
rect 28816 21558 28868 21564
rect 28828 21457 28856 21558
rect 28920 21554 28948 21830
rect 28998 21791 29054 21800
rect 28908 21548 28960 21554
rect 28908 21490 28960 21496
rect 29012 21457 29040 21791
rect 28814 21448 28870 21457
rect 28814 21383 28870 21392
rect 28998 21448 29054 21457
rect 28998 21383 29054 21392
rect 28816 21344 28868 21350
rect 28816 21286 28868 21292
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28998 21312 29054 21321
rect 28828 20466 28856 21286
rect 28816 20460 28868 20466
rect 28816 20402 28868 20408
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28814 20360 28870 20369
rect 28814 20295 28870 20304
rect 28724 20256 28776 20262
rect 28630 20224 28686 20233
rect 28724 20198 28776 20204
rect 28630 20159 28686 20168
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 28644 19417 28672 19450
rect 28630 19408 28686 19417
rect 28630 19343 28686 19352
rect 28552 19230 28672 19258
rect 28356 19168 28408 19174
rect 28177 19094 28212 19122
rect 28262 19136 28318 19145
rect 27837 19068 28145 19077
rect 27837 19066 27843 19068
rect 27899 19066 27923 19068
rect 27979 19066 28003 19068
rect 28059 19066 28083 19068
rect 28139 19066 28145 19068
rect 27899 19014 27901 19066
rect 28081 19014 28083 19066
rect 27837 19012 27843 19014
rect 27899 19012 27923 19014
rect 27979 19012 28003 19014
rect 28059 19012 28083 19014
rect 28139 19012 28145 19014
rect 27837 19003 28145 19012
rect 27712 18964 27764 18970
rect 27488 18244 27568 18272
rect 27632 18924 27712 18952
rect 27436 18226 27488 18232
rect 27448 18057 27476 18226
rect 27526 18184 27582 18193
rect 27526 18119 27582 18128
rect 27434 18048 27490 18057
rect 27434 17983 27490 17992
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27448 17513 27476 17614
rect 27540 17610 27568 18119
rect 27632 17746 27660 18924
rect 27712 18906 27764 18912
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 27896 18828 27948 18834
rect 27896 18770 27948 18776
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 27802 18728 27858 18737
rect 27802 18663 27858 18672
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27724 17921 27752 18362
rect 27816 18154 27844 18663
rect 27908 18358 27936 18770
rect 27896 18352 27948 18358
rect 27896 18294 27948 18300
rect 28000 18290 28028 18770
rect 28092 18698 28120 18906
rect 28177 18884 28205 19094
rect 28356 19110 28408 19116
rect 28262 19071 28318 19080
rect 28446 19000 28502 19009
rect 28356 18964 28408 18970
rect 28446 18935 28448 18944
rect 28356 18906 28408 18912
rect 28500 18935 28502 18944
rect 28448 18906 28500 18912
rect 28177 18856 28212 18884
rect 28080 18692 28132 18698
rect 28080 18634 28132 18640
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 28184 18222 28212 18856
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28080 18216 28132 18222
rect 28078 18184 28080 18193
rect 28172 18216 28224 18222
rect 28132 18184 28134 18193
rect 27804 18148 27856 18154
rect 28172 18158 28224 18164
rect 28078 18119 28134 18128
rect 27804 18090 27856 18096
rect 27837 17980 28145 17989
rect 27837 17978 27843 17980
rect 27899 17978 27923 17980
rect 27979 17978 28003 17980
rect 28059 17978 28083 17980
rect 28139 17978 28145 17980
rect 27899 17926 27901 17978
rect 28081 17926 28083 17978
rect 27837 17924 27843 17926
rect 27899 17924 27923 17926
rect 27979 17924 28003 17926
rect 28059 17924 28083 17926
rect 28139 17924 28145 17926
rect 27710 17912 27766 17921
rect 27837 17915 28145 17924
rect 28276 17921 28304 18226
rect 28262 17912 28318 17921
rect 27710 17847 27766 17856
rect 28172 17876 28224 17882
rect 28262 17847 28318 17856
rect 28172 17818 28224 17824
rect 27710 17776 27766 17785
rect 27620 17740 27672 17746
rect 27710 17711 27712 17720
rect 27620 17682 27672 17688
rect 27764 17711 27766 17720
rect 27712 17682 27764 17688
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 27528 17604 27580 17610
rect 27528 17546 27580 17552
rect 28092 17513 28120 17614
rect 27434 17504 27490 17513
rect 27434 17439 27490 17448
rect 28078 17504 28134 17513
rect 28078 17439 28134 17448
rect 28184 17338 28212 17818
rect 28368 17814 28396 18906
rect 28540 18828 28592 18834
rect 28540 18770 28592 18776
rect 28448 18624 28500 18630
rect 28448 18566 28500 18572
rect 28460 18290 28488 18566
rect 28552 18329 28580 18770
rect 28538 18320 28594 18329
rect 28448 18284 28500 18290
rect 28538 18255 28594 18264
rect 28448 18226 28500 18232
rect 28356 17808 28408 17814
rect 28356 17750 28408 17756
rect 28264 17536 28316 17542
rect 28262 17504 28264 17513
rect 28316 17504 28318 17513
rect 28262 17439 28318 17448
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 27436 17264 27488 17270
rect 27712 17264 27764 17270
rect 27436 17206 27488 17212
rect 27632 17224 27712 17252
rect 27448 16833 27476 17206
rect 27528 17060 27580 17066
rect 27528 17002 27580 17008
rect 27434 16824 27490 16833
rect 27434 16759 27490 16768
rect 27434 16688 27490 16697
rect 27434 16623 27436 16632
rect 27488 16623 27490 16632
rect 27436 16594 27488 16600
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27448 16114 27476 16390
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27436 15632 27488 15638
rect 27436 15574 27488 15580
rect 27448 14414 27476 15574
rect 27540 15570 27568 17002
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27632 15450 27660 17224
rect 27712 17206 27764 17212
rect 27837 16892 28145 16901
rect 27837 16890 27843 16892
rect 27899 16890 27923 16892
rect 27979 16890 28003 16892
rect 28059 16890 28083 16892
rect 28139 16890 28145 16892
rect 27899 16838 27901 16890
rect 28081 16838 28083 16890
rect 27837 16836 27843 16838
rect 27899 16836 27923 16838
rect 27979 16836 28003 16838
rect 28059 16836 28083 16838
rect 28139 16836 28145 16838
rect 27837 16827 28145 16836
rect 28184 16697 28212 17274
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28264 17060 28316 17066
rect 28264 17002 28316 17008
rect 28276 16726 28304 17002
rect 28264 16720 28316 16726
rect 28170 16688 28226 16697
rect 28264 16662 28316 16668
rect 28170 16623 28226 16632
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27540 15422 27660 15450
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27448 13326 27476 14350
rect 27540 13954 27568 15422
rect 27724 15416 27752 16526
rect 28368 16402 28396 17138
rect 28460 16794 28488 18226
rect 28644 18193 28672 19230
rect 28630 18184 28686 18193
rect 28630 18119 28686 18128
rect 28630 17776 28686 17785
rect 28630 17711 28686 17720
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28552 17338 28580 17478
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 28552 17241 28580 17274
rect 28538 17232 28594 17241
rect 28538 17167 28594 17176
rect 28538 16824 28594 16833
rect 28448 16788 28500 16794
rect 28538 16759 28594 16768
rect 28448 16730 28500 16736
rect 28276 16374 28396 16402
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28078 16280 28134 16289
rect 28078 16215 28134 16224
rect 27896 16176 27948 16182
rect 27896 16118 27948 16124
rect 27908 15978 27936 16118
rect 28092 15978 28120 16215
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 28080 15972 28132 15978
rect 28080 15914 28132 15920
rect 27837 15804 28145 15813
rect 27837 15802 27843 15804
rect 27899 15802 27923 15804
rect 27979 15802 28003 15804
rect 28059 15802 28083 15804
rect 28139 15802 28145 15804
rect 27899 15750 27901 15802
rect 28081 15750 28083 15802
rect 27837 15748 27843 15750
rect 27899 15748 27923 15750
rect 27979 15748 28003 15750
rect 28059 15748 28083 15750
rect 28139 15748 28145 15750
rect 27837 15739 28145 15748
rect 28276 15722 28304 16374
rect 28460 16289 28488 16390
rect 28446 16280 28502 16289
rect 28356 16244 28408 16250
rect 28446 16215 28502 16224
rect 28356 16186 28408 16192
rect 28368 16096 28396 16186
rect 28368 16068 28488 16096
rect 27896 15700 27948 15706
rect 28184 15694 28304 15722
rect 28184 15688 28212 15694
rect 27948 15660 28212 15688
rect 27896 15642 27948 15648
rect 27804 15428 27856 15434
rect 27724 15388 27804 15416
rect 27804 15370 27856 15376
rect 27816 15094 27844 15370
rect 27894 15328 27950 15337
rect 27894 15263 27950 15272
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27632 14074 27660 14758
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27540 13926 27660 13954
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 27342 13016 27398 13025
rect 27342 12951 27344 12960
rect 27396 12951 27398 12960
rect 27344 12922 27396 12928
rect 27540 12850 27568 13262
rect 27632 13258 27660 13926
rect 27724 13462 27752 14962
rect 27908 14958 27936 15263
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27896 14952 27948 14958
rect 27896 14894 27948 14900
rect 28000 14804 28028 14962
rect 28184 14906 28212 15660
rect 28264 15632 28316 15638
rect 28264 15574 28316 15580
rect 28276 15502 28304 15574
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28356 15428 28408 15434
rect 28356 15370 28408 15376
rect 28184 14878 28304 14906
rect 28172 14816 28224 14822
rect 28000 14776 28172 14804
rect 28172 14758 28224 14764
rect 27837 14716 28145 14725
rect 27837 14714 27843 14716
rect 27899 14714 27923 14716
rect 27979 14714 28003 14716
rect 28059 14714 28083 14716
rect 28139 14714 28145 14716
rect 27899 14662 27901 14714
rect 28081 14662 28083 14714
rect 27837 14660 27843 14662
rect 27899 14660 27923 14662
rect 27979 14660 28003 14662
rect 28059 14660 28083 14662
rect 28139 14660 28145 14662
rect 27837 14651 28145 14660
rect 27804 14544 27856 14550
rect 27804 14486 27856 14492
rect 27896 14544 27948 14550
rect 27896 14486 27948 14492
rect 28078 14512 28134 14521
rect 27816 13938 27844 14486
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27908 13734 27936 14486
rect 28078 14447 28134 14456
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 28000 13802 28028 14214
rect 28092 13938 28120 14447
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28170 13832 28226 13841
rect 27988 13796 28040 13802
rect 28170 13767 28226 13776
rect 27988 13738 28040 13744
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27837 13628 28145 13637
rect 27837 13626 27843 13628
rect 27899 13626 27923 13628
rect 27979 13626 28003 13628
rect 28059 13626 28083 13628
rect 28139 13626 28145 13628
rect 27899 13574 27901 13626
rect 28081 13574 28083 13626
rect 27837 13572 27843 13574
rect 27899 13572 27923 13574
rect 27979 13572 28003 13574
rect 28059 13572 28083 13574
rect 28139 13572 28145 13574
rect 27837 13563 28145 13572
rect 28184 13530 28212 13767
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 27712 13456 27764 13462
rect 27712 13398 27764 13404
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 28276 13190 28304 14878
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 27710 12880 27766 12889
rect 27528 12844 27580 12850
rect 27710 12815 27766 12824
rect 27528 12786 27580 12792
rect 27252 12300 27304 12306
rect 27252 12242 27304 12248
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27068 11008 27120 11014
rect 27068 10950 27120 10956
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26884 9988 26936 9994
rect 26884 9930 26936 9936
rect 27080 8634 27108 10950
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26608 7472 26660 7478
rect 26608 7414 26660 7420
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26252 5166 26280 6598
rect 26620 5778 26648 7414
rect 26792 7404 26844 7410
rect 26792 7346 26844 7352
rect 26804 6662 26832 7346
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 26608 5772 26660 5778
rect 26608 5714 26660 5720
rect 26240 5160 26292 5166
rect 26240 5102 26292 5108
rect 26148 4752 26200 4758
rect 26148 4694 26200 4700
rect 26804 4622 26832 6598
rect 27172 5302 27200 12038
rect 27540 11830 27568 12786
rect 27618 12472 27674 12481
rect 27618 12407 27674 12416
rect 27632 11830 27660 12407
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 27620 11824 27672 11830
rect 27620 11766 27672 11772
rect 27724 11558 27752 12815
rect 27837 12540 28145 12549
rect 27837 12538 27843 12540
rect 27899 12538 27923 12540
rect 27979 12538 28003 12540
rect 28059 12538 28083 12540
rect 28139 12538 28145 12540
rect 27899 12486 27901 12538
rect 28081 12486 28083 12538
rect 27837 12484 27843 12486
rect 27899 12484 27923 12486
rect 27979 12484 28003 12486
rect 28059 12484 28083 12486
rect 28139 12484 28145 12486
rect 27837 12475 28145 12484
rect 28172 12436 28224 12442
rect 28172 12378 28224 12384
rect 28080 12368 28132 12374
rect 28080 12310 28132 12316
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 28000 11626 28028 12038
rect 28092 11898 28120 12310
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 27988 11620 28040 11626
rect 27988 11562 28040 11568
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27620 11212 27672 11218
rect 27620 11154 27672 11160
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27264 7886 27292 10950
rect 27436 9104 27488 9110
rect 27436 9046 27488 9052
rect 27448 8090 27476 9046
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 27448 6914 27476 8026
rect 27540 7478 27568 11018
rect 27632 10985 27660 11154
rect 27724 11014 27752 11494
rect 27837 11452 28145 11461
rect 27837 11450 27843 11452
rect 27899 11450 27923 11452
rect 27979 11450 28003 11452
rect 28059 11450 28083 11452
rect 28139 11450 28145 11452
rect 27899 11398 27901 11450
rect 28081 11398 28083 11450
rect 27837 11396 27843 11398
rect 27899 11396 27923 11398
rect 27979 11396 28003 11398
rect 28059 11396 28083 11398
rect 28139 11396 28145 11398
rect 27837 11387 28145 11396
rect 27988 11348 28040 11354
rect 27988 11290 28040 11296
rect 28000 11082 28028 11290
rect 28184 11286 28212 12378
rect 28276 11898 28304 13126
rect 28368 12714 28396 15370
rect 28460 15366 28488 16068
rect 28448 15360 28500 15366
rect 28448 15302 28500 15308
rect 28460 14958 28488 15302
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28460 14550 28488 14894
rect 28448 14544 28500 14550
rect 28448 14486 28500 14492
rect 28446 14376 28502 14385
rect 28446 14311 28448 14320
rect 28500 14311 28502 14320
rect 28448 14282 28500 14288
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 28356 12708 28408 12714
rect 28356 12650 28408 12656
rect 28460 12442 28488 13874
rect 28552 13530 28580 16759
rect 28644 15609 28672 17711
rect 28630 15600 28686 15609
rect 28630 15535 28632 15544
rect 28684 15535 28686 15544
rect 28632 15506 28684 15512
rect 28632 15360 28684 15366
rect 28632 15302 28684 15308
rect 28644 15162 28672 15302
rect 28632 15156 28684 15162
rect 28632 15098 28684 15104
rect 28630 15056 28686 15065
rect 28630 14991 28632 15000
rect 28684 14991 28686 15000
rect 28632 14962 28684 14968
rect 28632 14884 28684 14890
rect 28632 14826 28684 14832
rect 28644 14793 28672 14826
rect 28630 14784 28686 14793
rect 28630 14719 28686 14728
rect 28630 14648 28686 14657
rect 28630 14583 28686 14592
rect 28644 14482 28672 14583
rect 28632 14476 28684 14482
rect 28632 14418 28684 14424
rect 28736 14226 28764 20198
rect 28828 19145 28856 20295
rect 28814 19136 28870 19145
rect 28920 19122 28948 21286
rect 28998 21247 29054 21256
rect 29012 21146 29040 21247
rect 29000 21140 29052 21146
rect 29000 21082 29052 21088
rect 29104 20913 29132 21898
rect 29090 20904 29146 20913
rect 29090 20839 29146 20848
rect 29092 20528 29144 20534
rect 29092 20470 29144 20476
rect 28998 20360 29054 20369
rect 28998 20295 29054 20304
rect 29012 20058 29040 20295
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 28998 19408 29054 19417
rect 28998 19343 29000 19352
rect 29052 19343 29054 19352
rect 29000 19314 29052 19320
rect 28814 19071 28870 19080
rect 28904 19094 28948 19122
rect 28904 18986 28932 19094
rect 28828 18958 28932 18986
rect 28828 18884 28856 18958
rect 28828 18856 28932 18884
rect 28904 18748 28932 18856
rect 28904 18720 28948 18748
rect 28816 18216 28868 18222
rect 28816 18158 28868 18164
rect 28828 16522 28856 18158
rect 28920 17338 28948 18720
rect 29012 18442 29040 19314
rect 29104 18601 29132 20470
rect 29196 19310 29224 22578
rect 29276 22500 29328 22506
rect 29276 22442 29328 22448
rect 29288 22234 29316 22442
rect 29276 22228 29328 22234
rect 29276 22170 29328 22176
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29184 19304 29236 19310
rect 29184 19246 29236 19252
rect 29184 19168 29236 19174
rect 29182 19136 29184 19145
rect 29236 19136 29238 19145
rect 29182 19071 29238 19080
rect 29182 19000 29238 19009
rect 29182 18935 29238 18944
rect 29196 18630 29224 18935
rect 29184 18624 29236 18630
rect 29090 18592 29146 18601
rect 29184 18566 29236 18572
rect 29090 18527 29146 18536
rect 29012 18414 29224 18442
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 28906 17232 28962 17241
rect 28906 17167 28962 17176
rect 28816 16516 28868 16522
rect 28816 16458 28868 16464
rect 28828 15706 28856 16458
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 28816 15156 28868 15162
rect 28816 15098 28868 15104
rect 28828 14278 28856 15098
rect 28644 14198 28764 14226
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28644 14074 28672 14198
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28724 14068 28776 14074
rect 28724 14010 28776 14016
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28736 13297 28764 14010
rect 28722 13288 28778 13297
rect 28722 13223 28778 13232
rect 28538 12880 28594 12889
rect 28538 12815 28594 12824
rect 28552 12714 28580 12815
rect 28540 12708 28592 12714
rect 28540 12650 28592 12656
rect 28448 12436 28500 12442
rect 28448 12378 28500 12384
rect 28552 12322 28580 12650
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28356 12300 28408 12306
rect 28356 12242 28408 12248
rect 28460 12294 28580 12322
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28172 11280 28224 11286
rect 28172 11222 28224 11228
rect 28276 11150 28304 11834
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 27988 11076 28040 11082
rect 27988 11018 28040 11024
rect 27712 11008 27764 11014
rect 27618 10976 27674 10985
rect 27712 10950 27764 10956
rect 27618 10911 27674 10920
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27724 9042 27752 10406
rect 27837 10364 28145 10373
rect 27837 10362 27843 10364
rect 27899 10362 27923 10364
rect 27979 10362 28003 10364
rect 28059 10362 28083 10364
rect 28139 10362 28145 10364
rect 27899 10310 27901 10362
rect 28081 10310 28083 10362
rect 27837 10308 27843 10310
rect 27899 10308 27923 10310
rect 27979 10308 28003 10310
rect 28059 10308 28083 10310
rect 28139 10308 28145 10310
rect 27837 10299 28145 10308
rect 28276 10266 28304 11086
rect 28368 10538 28396 12242
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28264 10260 28316 10266
rect 28184 10220 28264 10248
rect 27837 9276 28145 9285
rect 27837 9274 27843 9276
rect 27899 9274 27923 9276
rect 27979 9274 28003 9276
rect 28059 9274 28083 9276
rect 28139 9274 28145 9276
rect 27899 9222 27901 9274
rect 28081 9222 28083 9274
rect 27837 9220 27843 9222
rect 27899 9220 27923 9222
rect 27979 9220 28003 9222
rect 28059 9220 28083 9222
rect 28139 9220 28145 9222
rect 27837 9211 28145 9220
rect 28184 9110 28212 10220
rect 28264 10202 28316 10208
rect 28368 10146 28396 10474
rect 28276 10118 28396 10146
rect 28172 9104 28224 9110
rect 28172 9046 28224 9052
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27837 8188 28145 8197
rect 27837 8186 27843 8188
rect 27899 8186 27923 8188
rect 27979 8186 28003 8188
rect 28059 8186 28083 8188
rect 28139 8186 28145 8188
rect 27899 8134 27901 8186
rect 28081 8134 28083 8186
rect 27837 8132 27843 8134
rect 27899 8132 27923 8134
rect 27979 8132 28003 8134
rect 28059 8132 28083 8134
rect 28139 8132 28145 8134
rect 27837 8123 28145 8132
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27632 7857 27660 7890
rect 27618 7848 27674 7857
rect 27618 7783 27674 7792
rect 27528 7472 27580 7478
rect 27528 7414 27580 7420
rect 27264 6886 27476 6914
rect 27160 5296 27212 5302
rect 27160 5238 27212 5244
rect 27264 4690 27292 6886
rect 27632 6730 27660 7783
rect 27837 7100 28145 7109
rect 27837 7098 27843 7100
rect 27899 7098 27923 7100
rect 27979 7098 28003 7100
rect 28059 7098 28083 7100
rect 28139 7098 28145 7100
rect 27899 7046 27901 7098
rect 28081 7046 28083 7098
rect 27837 7044 27843 7046
rect 27899 7044 27923 7046
rect 27979 7044 28003 7046
rect 28059 7044 28083 7046
rect 28139 7044 28145 7046
rect 27837 7035 28145 7044
rect 27620 6724 27672 6730
rect 27620 6666 27672 6672
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27632 5574 27660 6190
rect 27712 6112 27764 6118
rect 27712 6054 27764 6060
rect 27724 5846 27752 6054
rect 27837 6012 28145 6021
rect 27837 6010 27843 6012
rect 27899 6010 27923 6012
rect 27979 6010 28003 6012
rect 28059 6010 28083 6012
rect 28139 6010 28145 6012
rect 27899 5958 27901 6010
rect 28081 5958 28083 6010
rect 27837 5956 27843 5958
rect 27899 5956 27923 5958
rect 27979 5956 28003 5958
rect 28059 5956 28083 5958
rect 28139 5956 28145 5958
rect 27837 5947 28145 5956
rect 28276 5846 28304 10118
rect 28460 9926 28488 12294
rect 28538 11112 28594 11121
rect 28538 11047 28594 11056
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28552 9042 28580 11047
rect 28540 9036 28592 9042
rect 28540 8978 28592 8984
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28368 8090 28396 8910
rect 28448 8424 28500 8430
rect 28448 8366 28500 8372
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28368 7818 28396 8026
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 27712 5840 27764 5846
rect 27712 5782 27764 5788
rect 28264 5840 28316 5846
rect 28264 5782 28316 5788
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 28356 5568 28408 5574
rect 28356 5510 28408 5516
rect 28368 5030 28396 5510
rect 28460 5030 28488 8366
rect 28552 7478 28580 8978
rect 28540 7472 28592 7478
rect 28540 7414 28592 7420
rect 28644 5137 28672 12582
rect 28828 12374 28856 14214
rect 28920 13938 28948 17167
rect 29012 17066 29040 18226
rect 29196 18222 29224 18414
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 29000 17060 29052 17066
rect 29000 17002 29052 17008
rect 28998 16688 29054 16697
rect 28998 16623 29054 16632
rect 29012 16590 29040 16623
rect 29000 16584 29052 16590
rect 29000 16526 29052 16532
rect 29104 16436 29132 17614
rect 29196 17338 29224 18158
rect 29288 18086 29316 21966
rect 29472 21468 29500 23530
rect 29564 23118 29592 23666
rect 29656 23118 29684 23802
rect 29840 23633 29868 24006
rect 29826 23624 29882 23633
rect 29736 23588 29788 23594
rect 29826 23559 29882 23568
rect 29736 23530 29788 23536
rect 29748 23322 29776 23530
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29736 23180 29788 23186
rect 29736 23122 29788 23128
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29644 23112 29696 23118
rect 29644 23054 29696 23060
rect 29656 22953 29684 23054
rect 29642 22944 29698 22953
rect 29642 22879 29698 22888
rect 29748 22817 29776 23122
rect 29826 23080 29882 23089
rect 29826 23015 29882 23024
rect 29734 22808 29790 22817
rect 29734 22743 29790 22752
rect 29644 22704 29696 22710
rect 29644 22646 29696 22652
rect 29552 22636 29604 22642
rect 29552 22578 29604 22584
rect 29564 22030 29592 22578
rect 29656 22506 29684 22646
rect 29840 22574 29868 23015
rect 29828 22568 29880 22574
rect 29828 22510 29880 22516
rect 29644 22500 29696 22506
rect 29644 22442 29696 22448
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29550 21856 29606 21865
rect 29550 21791 29606 21800
rect 29564 21622 29592 21791
rect 29552 21616 29604 21622
rect 29552 21558 29604 21564
rect 29472 21440 29592 21468
rect 29368 21412 29420 21418
rect 29368 21354 29420 21360
rect 29380 21146 29408 21354
rect 29460 21344 29512 21350
rect 29460 21286 29512 21292
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29368 20800 29420 20806
rect 29472 20777 29500 21286
rect 29368 20742 29420 20748
rect 29458 20768 29514 20777
rect 29380 18748 29408 20742
rect 29458 20703 29514 20712
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29472 19310 29500 20402
rect 29460 19304 29512 19310
rect 29460 19246 29512 19252
rect 29564 18970 29592 21440
rect 29656 21049 29684 21966
rect 29828 21956 29880 21962
rect 29828 21898 29880 21904
rect 29734 21720 29790 21729
rect 29840 21690 29868 21898
rect 29932 21865 29960 24278
rect 30010 23760 30066 23769
rect 30010 23695 30012 23704
rect 30064 23695 30066 23704
rect 30012 23666 30064 23672
rect 30116 23610 30144 25230
rect 30208 23866 30236 26930
rect 30196 23860 30248 23866
rect 30196 23802 30248 23808
rect 30194 23760 30250 23769
rect 30194 23695 30250 23704
rect 30024 23582 30144 23610
rect 30024 23202 30052 23582
rect 30102 23352 30158 23361
rect 30208 23322 30236 23695
rect 30300 23633 30328 27814
rect 30484 27418 30512 30670
rect 30576 30598 30604 31726
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30656 31136 30708 31142
rect 30656 31078 30708 31084
rect 30564 30592 30616 30598
rect 30564 30534 30616 30540
rect 30576 30433 30604 30534
rect 30562 30424 30618 30433
rect 30562 30359 30618 30368
rect 30564 30048 30616 30054
rect 30564 29990 30616 29996
rect 30576 28558 30604 29990
rect 30564 28552 30616 28558
rect 30668 28529 30696 31078
rect 30564 28494 30616 28500
rect 30654 28520 30710 28529
rect 30654 28455 30710 28464
rect 30760 28234 30788 31282
rect 30576 28206 30788 28234
rect 30576 27674 30604 28206
rect 30748 28144 30800 28150
rect 30748 28086 30800 28092
rect 30654 27704 30710 27713
rect 30564 27668 30616 27674
rect 30654 27639 30710 27648
rect 30564 27610 30616 27616
rect 30564 27532 30616 27538
rect 30564 27474 30616 27480
rect 30392 27390 30512 27418
rect 30392 26042 30420 27390
rect 30470 27296 30526 27305
rect 30470 27231 30526 27240
rect 30484 27130 30512 27231
rect 30472 27124 30524 27130
rect 30472 27066 30524 27072
rect 30380 26036 30432 26042
rect 30380 25978 30432 25984
rect 30378 25936 30434 25945
rect 30378 25871 30380 25880
rect 30432 25871 30434 25880
rect 30380 25842 30432 25848
rect 30484 25702 30512 27066
rect 30472 25696 30524 25702
rect 30472 25638 30524 25644
rect 30380 25356 30432 25362
rect 30380 25298 30432 25304
rect 30392 24818 30420 25298
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30286 23624 30342 23633
rect 30286 23559 30342 23568
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30102 23287 30104 23296
rect 30156 23287 30158 23296
rect 30196 23316 30248 23322
rect 30104 23258 30156 23264
rect 30196 23258 30248 23264
rect 30024 23174 30236 23202
rect 30300 23186 30328 23462
rect 30104 22432 30156 22438
rect 30104 22374 30156 22380
rect 30010 22128 30066 22137
rect 30010 22063 30066 22072
rect 29918 21856 29974 21865
rect 29918 21791 29974 21800
rect 29918 21720 29974 21729
rect 29734 21655 29790 21664
rect 29828 21684 29880 21690
rect 29748 21078 29776 21655
rect 29918 21655 29974 21664
rect 29828 21626 29880 21632
rect 29932 21622 29960 21655
rect 29920 21616 29972 21622
rect 29920 21558 29972 21564
rect 30024 21078 30052 22063
rect 30116 22030 30144 22374
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30104 21888 30156 21894
rect 30104 21830 30156 21836
rect 29736 21072 29788 21078
rect 29642 21040 29698 21049
rect 30012 21072 30064 21078
rect 29736 21014 29788 21020
rect 29826 21040 29882 21049
rect 29642 20975 29698 20984
rect 30012 21014 30064 21020
rect 29826 20975 29828 20984
rect 29880 20975 29882 20984
rect 29828 20946 29880 20952
rect 30010 20904 30066 20913
rect 29644 20868 29696 20874
rect 30010 20839 30066 20848
rect 29644 20810 29696 20816
rect 29656 20777 29684 20810
rect 29736 20800 29788 20806
rect 29642 20768 29698 20777
rect 29918 20768 29974 20777
rect 29736 20742 29788 20748
rect 29642 20703 29698 20712
rect 29748 20602 29776 20742
rect 29840 20726 29918 20754
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29734 20496 29790 20505
rect 29734 20431 29790 20440
rect 29644 20392 29696 20398
rect 29644 20334 29696 20340
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29380 18720 29500 18748
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29380 18329 29408 18566
rect 29366 18320 29422 18329
rect 29472 18290 29500 18720
rect 29656 18290 29684 20334
rect 29748 19786 29776 20431
rect 29736 19780 29788 19786
rect 29736 19722 29788 19728
rect 29366 18255 29422 18264
rect 29460 18284 29512 18290
rect 29276 18080 29328 18086
rect 29276 18022 29328 18028
rect 29380 17785 29408 18255
rect 29460 18226 29512 18232
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29366 17776 29422 17785
rect 29366 17711 29422 17720
rect 29380 17610 29408 17711
rect 29368 17604 29420 17610
rect 29368 17546 29420 17552
rect 29276 17536 29328 17542
rect 29276 17478 29328 17484
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 29196 17202 29224 17274
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29182 17096 29238 17105
rect 29182 17031 29184 17040
rect 29236 17031 29238 17040
rect 29184 17002 29236 17008
rect 29288 16969 29316 17478
rect 29368 17196 29420 17202
rect 29368 17138 29420 17144
rect 29274 16960 29330 16969
rect 29274 16895 29330 16904
rect 29380 16640 29408 17138
rect 29472 17134 29500 18226
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29460 17128 29512 17134
rect 29460 17070 29512 17076
rect 29288 16612 29408 16640
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29012 16408 29132 16436
rect 29012 16289 29040 16408
rect 28998 16280 29054 16289
rect 29196 16266 29224 16526
rect 29288 16425 29316 16612
rect 29366 16552 29422 16561
rect 29366 16487 29422 16496
rect 29274 16416 29330 16425
rect 29274 16351 29330 16360
rect 28998 16215 29054 16224
rect 29104 16238 29224 16266
rect 29012 15706 29040 16215
rect 29104 16017 29132 16238
rect 29184 16108 29236 16114
rect 29184 16050 29236 16056
rect 29276 16108 29328 16114
rect 29276 16050 29328 16056
rect 29090 16008 29146 16017
rect 29090 15943 29146 15952
rect 29092 15904 29144 15910
rect 29196 15881 29224 16050
rect 29092 15846 29144 15852
rect 29182 15872 29238 15881
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 29104 15638 29132 15846
rect 29182 15807 29238 15816
rect 29092 15632 29144 15638
rect 29092 15574 29144 15580
rect 29104 14940 29132 15574
rect 29196 15366 29224 15807
rect 29288 15473 29316 16050
rect 29380 16046 29408 16487
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 29274 15464 29330 15473
rect 29274 15399 29330 15408
rect 29184 15360 29236 15366
rect 29184 15302 29236 15308
rect 29182 15192 29238 15201
rect 29182 15127 29238 15136
rect 29012 14912 29132 14940
rect 29012 14521 29040 14912
rect 29196 14890 29224 15127
rect 29184 14884 29236 14890
rect 29184 14826 29236 14832
rect 29092 14816 29144 14822
rect 29092 14758 29144 14764
rect 28998 14512 29054 14521
rect 28998 14447 29054 14456
rect 29000 14408 29052 14414
rect 29000 14350 29052 14356
rect 29012 14006 29040 14350
rect 29104 14113 29132 14758
rect 29276 14340 29328 14346
rect 29276 14282 29328 14288
rect 29090 14104 29146 14113
rect 29288 14090 29316 14282
rect 29380 14249 29408 15846
rect 29472 15502 29500 17070
rect 29564 16833 29592 17682
rect 29550 16824 29606 16833
rect 29550 16759 29606 16768
rect 29656 16454 29684 18226
rect 29734 18184 29790 18193
rect 29840 18154 29868 20726
rect 29918 20703 29974 20712
rect 29920 20528 29972 20534
rect 29918 20496 29920 20505
rect 29972 20496 29974 20505
rect 29918 20431 29974 20440
rect 30024 20330 30052 20839
rect 30116 20380 30144 21830
rect 30208 21010 30236 23174
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30288 23044 30340 23050
rect 30288 22986 30340 22992
rect 30300 22778 30328 22986
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30392 22642 30420 24754
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30288 22432 30340 22438
rect 30288 22374 30340 22380
rect 30300 22166 30328 22374
rect 30288 22160 30340 22166
rect 30288 22102 30340 22108
rect 30380 22024 30432 22030
rect 30286 21992 30342 22001
rect 30380 21966 30432 21972
rect 30286 21927 30342 21936
rect 30300 21894 30328 21927
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 30288 21548 30340 21554
rect 30288 21490 30340 21496
rect 30300 21026 30328 21490
rect 30392 21486 30420 21966
rect 30380 21480 30432 21486
rect 30380 21422 30432 21428
rect 30196 21004 30248 21010
rect 30300 20998 30420 21026
rect 30196 20946 30248 20952
rect 30288 20936 30340 20942
rect 30194 20904 30250 20913
rect 30288 20878 30340 20884
rect 30194 20839 30250 20848
rect 30208 20806 30236 20839
rect 30196 20800 30248 20806
rect 30196 20742 30248 20748
rect 30300 20641 30328 20878
rect 30392 20777 30420 20998
rect 30378 20768 30434 20777
rect 30378 20703 30434 20712
rect 30286 20632 30342 20641
rect 30286 20567 30342 20576
rect 30116 20352 30420 20380
rect 30484 20369 30512 25638
rect 30576 25430 30604 27474
rect 30564 25424 30616 25430
rect 30564 25366 30616 25372
rect 30564 25288 30616 25294
rect 30564 25230 30616 25236
rect 30576 23730 30604 25230
rect 30668 23866 30696 27639
rect 30760 26042 30788 28086
rect 30852 26602 30880 32166
rect 31208 31952 31260 31958
rect 31208 31894 31260 31900
rect 31220 31793 31248 31894
rect 31206 31784 31262 31793
rect 31206 31719 31262 31728
rect 31678 31580 31986 31589
rect 31678 31578 31684 31580
rect 31740 31578 31764 31580
rect 31820 31578 31844 31580
rect 31900 31578 31924 31580
rect 31980 31578 31986 31580
rect 31740 31526 31742 31578
rect 31922 31526 31924 31578
rect 31678 31524 31684 31526
rect 31740 31524 31764 31526
rect 31820 31524 31844 31526
rect 31900 31524 31924 31526
rect 31980 31524 31986 31526
rect 31678 31515 31986 31524
rect 32128 31272 32180 31278
rect 32128 31214 32180 31220
rect 32036 31136 32088 31142
rect 32036 31078 32088 31084
rect 31576 30728 31628 30734
rect 31576 30670 31628 30676
rect 30930 30560 30986 30569
rect 30930 30495 30986 30504
rect 30944 26858 30972 30495
rect 31482 30152 31538 30161
rect 31482 30087 31538 30096
rect 31208 30048 31260 30054
rect 31208 29990 31260 29996
rect 31220 29753 31248 29990
rect 31206 29744 31262 29753
rect 31206 29679 31262 29688
rect 31116 29640 31168 29646
rect 31116 29582 31168 29588
rect 31024 29504 31076 29510
rect 31024 29446 31076 29452
rect 31036 28082 31064 29446
rect 31024 28076 31076 28082
rect 31024 28018 31076 28024
rect 31024 27940 31076 27946
rect 31024 27882 31076 27888
rect 31036 27062 31064 27882
rect 31024 27056 31076 27062
rect 31024 26998 31076 27004
rect 30932 26852 30984 26858
rect 30932 26794 30984 26800
rect 30852 26586 30972 26602
rect 30852 26580 30984 26586
rect 30852 26574 30932 26580
rect 30984 26540 31064 26568
rect 30932 26522 30984 26528
rect 30840 26512 30892 26518
rect 30838 26480 30840 26489
rect 30892 26480 30894 26489
rect 30838 26415 30894 26424
rect 30840 26376 30892 26382
rect 30838 26344 30840 26353
rect 30892 26344 30894 26353
rect 30838 26279 30894 26288
rect 30840 26240 30892 26246
rect 30840 26182 30892 26188
rect 30932 26240 30984 26246
rect 31036 26217 31064 26540
rect 30932 26182 30984 26188
rect 31022 26208 31078 26217
rect 30748 26036 30800 26042
rect 30748 25978 30800 25984
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30760 24818 30788 25638
rect 30852 25430 30880 26182
rect 30944 25906 30972 26182
rect 31022 26143 31078 26152
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 30932 25764 30984 25770
rect 30932 25706 30984 25712
rect 30944 25498 30972 25706
rect 30932 25492 30984 25498
rect 30932 25434 30984 25440
rect 30840 25424 30892 25430
rect 30944 25401 30972 25434
rect 30840 25366 30892 25372
rect 30930 25392 30986 25401
rect 30930 25327 30986 25336
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30930 25120 30986 25129
rect 30852 24954 30880 25094
rect 30930 25055 30986 25064
rect 30840 24948 30892 24954
rect 30840 24890 30892 24896
rect 30944 24818 30972 25055
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30930 24712 30986 24721
rect 30840 24676 30892 24682
rect 30930 24647 30986 24656
rect 30840 24618 30892 24624
rect 30852 24585 30880 24618
rect 30838 24576 30894 24585
rect 30838 24511 30894 24520
rect 30748 24200 30800 24206
rect 30748 24142 30800 24148
rect 30656 23860 30708 23866
rect 30656 23802 30708 23808
rect 30564 23724 30616 23730
rect 30564 23666 30616 23672
rect 30576 23594 30604 23666
rect 30564 23588 30616 23594
rect 30564 23530 30616 23536
rect 30760 22982 30788 24142
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30852 24041 30880 24074
rect 30838 24032 30894 24041
rect 30838 23967 30894 23976
rect 30944 23730 30972 24647
rect 31036 24410 31064 26143
rect 31128 24993 31156 29582
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31208 29028 31260 29034
rect 31208 28970 31260 28976
rect 31220 27713 31248 28970
rect 31312 28558 31340 29446
rect 31392 28756 31444 28762
rect 31392 28698 31444 28704
rect 31300 28552 31352 28558
rect 31300 28494 31352 28500
rect 31300 28416 31352 28422
rect 31300 28358 31352 28364
rect 31206 27704 31262 27713
rect 31206 27639 31262 27648
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31220 26450 31248 26930
rect 31208 26444 31260 26450
rect 31208 26386 31260 26392
rect 31220 25838 31248 26386
rect 31208 25832 31260 25838
rect 31208 25774 31260 25780
rect 31208 25696 31260 25702
rect 31312 25673 31340 28358
rect 31208 25638 31260 25644
rect 31298 25664 31354 25673
rect 31114 24984 31170 24993
rect 31114 24919 31170 24928
rect 31116 24880 31168 24886
rect 31116 24822 31168 24828
rect 31024 24404 31076 24410
rect 31024 24346 31076 24352
rect 31024 24268 31076 24274
rect 31128 24256 31156 24822
rect 31220 24342 31248 25638
rect 31298 25599 31354 25608
rect 31298 25392 31354 25401
rect 31298 25327 31354 25336
rect 31208 24336 31260 24342
rect 31208 24278 31260 24284
rect 31076 24228 31156 24256
rect 31024 24210 31076 24216
rect 31312 24188 31340 25327
rect 31220 24160 31340 24188
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 31116 23248 31168 23254
rect 31022 23216 31078 23225
rect 31116 23190 31168 23196
rect 31022 23151 31024 23160
rect 31076 23151 31078 23160
rect 31024 23122 31076 23128
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 30748 22976 30800 22982
rect 30800 22936 30880 22964
rect 30748 22918 30800 22924
rect 30852 22574 30880 22936
rect 30944 22642 30972 23054
rect 31024 23044 31076 23050
rect 31024 22986 31076 22992
rect 31036 22778 31064 22986
rect 31024 22772 31076 22778
rect 31024 22714 31076 22720
rect 31128 22710 31156 23190
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30748 22568 30800 22574
rect 30748 22510 30800 22516
rect 30840 22568 30892 22574
rect 30840 22510 30892 22516
rect 30760 22438 30788 22510
rect 30748 22432 30800 22438
rect 30748 22374 30800 22380
rect 30930 22400 30986 22409
rect 30930 22335 30986 22344
rect 30564 22092 30616 22098
rect 30564 22034 30616 22040
rect 30576 20534 30604 22034
rect 30654 21992 30710 22001
rect 30654 21927 30710 21936
rect 30668 21554 30696 21927
rect 30748 21684 30800 21690
rect 30748 21626 30800 21632
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30656 21412 30708 21418
rect 30656 21354 30708 21360
rect 30564 20528 30616 20534
rect 30564 20470 30616 20476
rect 30564 20392 30616 20398
rect 30012 20324 30064 20330
rect 30064 20284 30144 20312
rect 30012 20266 30064 20272
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 29918 19544 29974 19553
rect 29918 19479 29974 19488
rect 29932 19446 29960 19479
rect 29920 19440 29972 19446
rect 30024 19417 30052 19654
rect 29920 19382 29972 19388
rect 30010 19408 30066 19417
rect 30010 19343 30066 19352
rect 29920 19304 29972 19310
rect 29920 19246 29972 19252
rect 29734 18119 29790 18128
rect 29828 18148 29880 18154
rect 29748 17746 29776 18119
rect 29828 18090 29880 18096
rect 29826 17912 29882 17921
rect 29826 17847 29882 17856
rect 29736 17740 29788 17746
rect 29736 17682 29788 17688
rect 29736 17604 29788 17610
rect 29736 17546 29788 17552
rect 29748 16454 29776 17546
rect 29840 17202 29868 17847
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 29644 16448 29696 16454
rect 29550 16416 29606 16425
rect 29644 16390 29696 16396
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 29550 16351 29606 16360
rect 29460 15496 29512 15502
rect 29460 15438 29512 15444
rect 29564 15314 29592 16351
rect 29644 16176 29696 16182
rect 29748 16164 29776 16390
rect 29696 16136 29776 16164
rect 29644 16118 29696 16124
rect 29644 15972 29696 15978
rect 29644 15914 29696 15920
rect 29656 15337 29684 15914
rect 29472 15286 29592 15314
rect 29642 15328 29698 15337
rect 29366 14240 29422 14249
rect 29366 14175 29422 14184
rect 29288 14062 29408 14090
rect 29090 14039 29146 14048
rect 29000 14000 29052 14006
rect 29000 13942 29052 13948
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 29000 13728 29052 13734
rect 29000 13670 29052 13676
rect 28908 13184 28960 13190
rect 28906 13152 28908 13161
rect 28960 13152 28962 13161
rect 28906 13087 28962 13096
rect 28816 12368 28868 12374
rect 28816 12310 28868 12316
rect 28724 12232 28776 12238
rect 28724 12174 28776 12180
rect 28736 10996 28764 12174
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28828 11257 28856 12038
rect 28814 11248 28870 11257
rect 28814 11183 28870 11192
rect 28816 11008 28868 11014
rect 28736 10968 28816 10996
rect 28816 10950 28868 10956
rect 28828 9586 28856 10950
rect 28920 9654 28948 13087
rect 29012 10606 29040 13670
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 29104 9738 29132 14039
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29184 13728 29236 13734
rect 29184 13670 29236 13676
rect 29196 13433 29224 13670
rect 29182 13424 29238 13433
rect 29182 13359 29238 13368
rect 29288 13326 29316 13874
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 29380 13172 29408 14062
rect 29288 13144 29408 13172
rect 29288 12306 29316 13144
rect 29368 12640 29420 12646
rect 29368 12582 29420 12588
rect 29276 12300 29328 12306
rect 29276 12242 29328 12248
rect 29380 12170 29408 12582
rect 29368 12164 29420 12170
rect 29368 12106 29420 12112
rect 29472 11694 29500 15286
rect 29642 15263 29698 15272
rect 29656 15144 29684 15263
rect 29564 15116 29684 15144
rect 29564 12866 29592 15116
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29736 15020 29788 15026
rect 29736 14962 29788 14968
rect 29656 14414 29684 14962
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29656 13977 29684 14350
rect 29642 13968 29698 13977
rect 29748 13938 29776 14962
rect 29840 14414 29868 17138
rect 29932 16250 29960 19246
rect 30116 18850 30144 20284
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30024 18834 30144 18850
rect 30012 18828 30144 18834
rect 30064 18822 30144 18828
rect 30012 18770 30064 18776
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30116 18601 30144 18702
rect 30102 18592 30158 18601
rect 30102 18527 30158 18536
rect 30208 18426 30236 19858
rect 30300 19718 30328 20198
rect 30288 19712 30340 19718
rect 30288 19654 30340 19660
rect 30288 19440 30340 19446
rect 30286 19408 30288 19417
rect 30340 19408 30342 19417
rect 30286 19343 30342 19352
rect 30288 19304 30340 19310
rect 30288 19246 30340 19252
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30024 18068 30052 18226
rect 30208 18193 30236 18226
rect 30300 18222 30328 19246
rect 30288 18216 30340 18222
rect 30194 18184 30250 18193
rect 30288 18158 30340 18164
rect 30194 18119 30250 18128
rect 30024 18040 30236 18068
rect 30102 17776 30158 17785
rect 30102 17711 30158 17720
rect 30012 17536 30064 17542
rect 30012 17478 30064 17484
rect 30024 17270 30052 17478
rect 30012 17264 30064 17270
rect 30012 17206 30064 17212
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 29932 16017 29960 16050
rect 29918 16008 29974 16017
rect 29918 15943 29974 15952
rect 29920 15360 29972 15366
rect 29920 15302 29972 15308
rect 29932 14822 29960 15302
rect 30024 15162 30052 17206
rect 30116 16250 30144 17711
rect 30104 16244 30156 16250
rect 30104 16186 30156 16192
rect 30208 16046 30236 18040
rect 30286 17912 30342 17921
rect 30286 17847 30342 17856
rect 30196 16040 30248 16046
rect 30196 15982 30248 15988
rect 30196 15632 30248 15638
rect 30300 15620 30328 17847
rect 30392 16561 30420 20352
rect 30470 20360 30526 20369
rect 30564 20334 30616 20340
rect 30470 20295 30526 20304
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30484 19961 30512 20198
rect 30470 19952 30526 19961
rect 30470 19887 30526 19896
rect 30472 19848 30524 19854
rect 30470 19816 30472 19825
rect 30524 19816 30526 19825
rect 30470 19751 30526 19760
rect 30472 19712 30524 19718
rect 30472 19654 30524 19660
rect 30484 19378 30512 19654
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30484 19009 30512 19314
rect 30470 19000 30526 19009
rect 30470 18935 30526 18944
rect 30470 18864 30526 18873
rect 30470 18799 30526 18808
rect 30484 18290 30512 18799
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 30472 17876 30524 17882
rect 30472 17818 30524 17824
rect 30484 17678 30512 17818
rect 30472 17672 30524 17678
rect 30472 17614 30524 17620
rect 30470 17368 30526 17377
rect 30470 17303 30472 17312
rect 30524 17303 30526 17312
rect 30472 17274 30524 17280
rect 30472 17196 30524 17202
rect 30472 17138 30524 17144
rect 30484 17105 30512 17138
rect 30470 17096 30526 17105
rect 30470 17031 30526 17040
rect 30472 16992 30524 16998
rect 30472 16934 30524 16940
rect 30378 16552 30434 16561
rect 30378 16487 30434 16496
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 30248 15592 30328 15620
rect 30196 15574 30248 15580
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30010 15056 30066 15065
rect 30010 14991 30066 15000
rect 30024 14958 30052 14991
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 29920 14816 29972 14822
rect 29920 14758 29972 14764
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 29828 14272 29880 14278
rect 29828 14214 29880 14220
rect 29642 13903 29698 13912
rect 29736 13932 29788 13938
rect 29736 13874 29788 13880
rect 29734 13832 29790 13841
rect 29734 13767 29790 13776
rect 29564 12838 29684 12866
rect 29460 11688 29512 11694
rect 29460 11630 29512 11636
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 29184 9920 29236 9926
rect 29184 9862 29236 9868
rect 29012 9710 29132 9738
rect 28908 9648 28960 9654
rect 28908 9590 28960 9596
rect 28816 9580 28868 9586
rect 28816 9522 28868 9528
rect 28816 8356 28868 8362
rect 28816 8298 28868 8304
rect 28828 8090 28856 8298
rect 28816 8084 28868 8090
rect 28816 8026 28868 8032
rect 28724 6248 28776 6254
rect 28722 6216 28724 6225
rect 28776 6216 28778 6225
rect 28722 6151 28778 6160
rect 29012 5914 29040 9710
rect 29092 8832 29144 8838
rect 29090 8800 29092 8809
rect 29144 8800 29146 8809
rect 29090 8735 29146 8744
rect 29196 8634 29224 9862
rect 29184 8628 29236 8634
rect 29184 8570 29236 8576
rect 29184 7948 29236 7954
rect 29184 7890 29236 7896
rect 29092 7812 29144 7818
rect 29092 7754 29144 7760
rect 29104 6186 29132 7754
rect 29092 6180 29144 6186
rect 29092 6122 29144 6128
rect 29196 5914 29224 7890
rect 29380 6905 29408 11494
rect 29366 6896 29422 6905
rect 29472 6866 29500 11630
rect 29656 11354 29684 12838
rect 29748 12714 29776 13767
rect 29840 12918 29868 14214
rect 30024 14074 30052 14758
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 30010 13968 30066 13977
rect 30010 13903 30066 13912
rect 30024 13530 30052 13903
rect 30012 13524 30064 13530
rect 30012 13466 30064 13472
rect 29828 12912 29880 12918
rect 29828 12854 29880 12860
rect 29736 12708 29788 12714
rect 29736 12650 29788 12656
rect 29644 11348 29696 11354
rect 29644 11290 29696 11296
rect 29748 11014 29776 12650
rect 30116 11098 30144 15098
rect 30208 15094 30236 15574
rect 30196 15088 30248 15094
rect 30196 15030 30248 15036
rect 30208 12102 30236 15030
rect 30286 14648 30342 14657
rect 30286 14583 30342 14592
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 29932 11070 30144 11098
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29642 10840 29698 10849
rect 29642 10775 29698 10784
rect 29656 9722 29684 10775
rect 29748 10033 29776 10950
rect 29932 10606 29960 11070
rect 29920 10600 29972 10606
rect 29918 10568 29920 10577
rect 29972 10568 29974 10577
rect 29918 10503 29974 10512
rect 29734 10024 29790 10033
rect 29734 9959 29790 9968
rect 29644 9716 29696 9722
rect 29644 9658 29696 9664
rect 29656 8974 29684 9658
rect 30208 9518 30236 12038
rect 30300 10266 30328 14583
rect 30392 14498 30420 16390
rect 30484 15434 30512 16934
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30470 15328 30526 15337
rect 30470 15263 30526 15272
rect 30484 15094 30512 15263
rect 30576 15162 30604 20334
rect 30668 19174 30696 21354
rect 30760 20097 30788 21626
rect 30840 21548 30892 21554
rect 30840 21490 30892 21496
rect 30852 21457 30880 21490
rect 30838 21448 30894 21457
rect 30838 21383 30894 21392
rect 30838 21312 30894 21321
rect 30838 21247 30894 21256
rect 30852 20874 30880 21247
rect 30840 20868 30892 20874
rect 30840 20810 30892 20816
rect 30840 20460 30892 20466
rect 30840 20402 30892 20408
rect 30746 20088 30802 20097
rect 30852 20058 30880 20402
rect 30944 20398 30972 22335
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 30932 20392 30984 20398
rect 30932 20334 30984 20340
rect 30746 20023 30802 20032
rect 30840 20052 30892 20058
rect 30840 19994 30892 20000
rect 30748 19916 30800 19922
rect 30748 19858 30800 19864
rect 30760 19242 30788 19858
rect 30748 19236 30800 19242
rect 30748 19178 30800 19184
rect 30656 19168 30708 19174
rect 30656 19110 30708 19116
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 30668 17377 30696 18634
rect 30760 18154 30788 18702
rect 30852 18601 30880 19994
rect 31036 19281 31064 21966
rect 31116 21888 31168 21894
rect 31116 21830 31168 21836
rect 31128 21593 31156 21830
rect 31114 21584 31170 21593
rect 31114 21519 31170 21528
rect 31116 21344 31168 21350
rect 31116 21286 31168 21292
rect 31128 21185 31156 21286
rect 31114 21176 31170 21185
rect 31114 21111 31170 21120
rect 31220 21060 31248 24160
rect 31404 23798 31432 28698
rect 31496 27130 31524 30087
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31484 26376 31536 26382
rect 31484 26318 31536 26324
rect 31496 24886 31524 26318
rect 31484 24880 31536 24886
rect 31484 24822 31536 24828
rect 31482 24712 31538 24721
rect 31482 24647 31538 24656
rect 31392 23792 31444 23798
rect 31392 23734 31444 23740
rect 31300 23656 31352 23662
rect 31300 23598 31352 23604
rect 31392 23656 31444 23662
rect 31392 23598 31444 23604
rect 31312 22817 31340 23598
rect 31298 22808 31354 22817
rect 31298 22743 31354 22752
rect 31298 22672 31354 22681
rect 31298 22607 31354 22616
rect 31312 21146 31340 22607
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 31128 21032 31248 21060
rect 31128 19990 31156 21032
rect 31300 20936 31352 20942
rect 31206 20904 31262 20913
rect 31300 20878 31352 20884
rect 31206 20839 31262 20848
rect 31116 19984 31168 19990
rect 31116 19926 31168 19932
rect 31116 19848 31168 19854
rect 31116 19790 31168 19796
rect 31128 19689 31156 19790
rect 31114 19680 31170 19689
rect 31114 19615 31170 19624
rect 31022 19272 31078 19281
rect 31022 19207 31078 19216
rect 30932 19168 30984 19174
rect 30932 19110 30984 19116
rect 30944 18834 30972 19110
rect 31116 18896 31168 18902
rect 31022 18864 31078 18873
rect 30932 18828 30984 18834
rect 31116 18838 31168 18844
rect 31022 18799 31078 18808
rect 30932 18770 30984 18776
rect 30838 18592 30894 18601
rect 30838 18527 30894 18536
rect 30838 18456 30894 18465
rect 30838 18391 30840 18400
rect 30892 18391 30894 18400
rect 30840 18362 30892 18368
rect 30838 18184 30894 18193
rect 30748 18148 30800 18154
rect 30838 18119 30894 18128
rect 30748 18090 30800 18096
rect 30760 18057 30788 18090
rect 30746 18048 30802 18057
rect 30746 17983 30802 17992
rect 30748 17808 30800 17814
rect 30748 17750 30800 17756
rect 30760 17678 30788 17750
rect 30748 17672 30800 17678
rect 30748 17614 30800 17620
rect 30654 17368 30710 17377
rect 30654 17303 30710 17312
rect 30760 17252 30788 17614
rect 30668 17224 30788 17252
rect 30668 16590 30696 17224
rect 30746 17096 30802 17105
rect 30746 17031 30802 17040
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 30668 16153 30696 16390
rect 30760 16182 30788 17031
rect 30748 16176 30800 16182
rect 30654 16144 30710 16153
rect 30748 16118 30800 16124
rect 30654 16079 30710 16088
rect 30746 16008 30802 16017
rect 30746 15943 30748 15952
rect 30800 15943 30802 15952
rect 30748 15914 30800 15920
rect 30746 15464 30802 15473
rect 30656 15428 30708 15434
rect 30746 15399 30802 15408
rect 30656 15370 30708 15376
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30472 15088 30524 15094
rect 30472 15030 30524 15036
rect 30470 14920 30526 14929
rect 30470 14855 30526 14864
rect 30484 14618 30512 14855
rect 30472 14612 30524 14618
rect 30472 14554 30524 14560
rect 30392 14470 30512 14498
rect 30378 14376 30434 14385
rect 30378 14311 30434 14320
rect 30392 11558 30420 14311
rect 30484 12238 30512 14470
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30472 11824 30524 11830
rect 30472 11766 30524 11772
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30288 10260 30340 10266
rect 30288 10202 30340 10208
rect 30196 9512 30248 9518
rect 30196 9454 30248 9460
rect 30104 9376 30156 9382
rect 30104 9318 30156 9324
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29734 8664 29790 8673
rect 29734 8599 29736 8608
rect 29788 8599 29790 8608
rect 29736 8570 29788 8576
rect 30116 8537 30144 9318
rect 30208 9178 30236 9454
rect 30196 9172 30248 9178
rect 30196 9114 30248 9120
rect 30300 8616 30328 10202
rect 30208 8588 30328 8616
rect 30102 8528 30158 8537
rect 30102 8463 30158 8472
rect 29736 8084 29788 8090
rect 29736 8026 29788 8032
rect 29366 6831 29422 6840
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29368 6792 29420 6798
rect 29368 6734 29420 6740
rect 29000 5908 29052 5914
rect 29000 5850 29052 5856
rect 29184 5908 29236 5914
rect 29184 5850 29236 5856
rect 29380 5166 29408 6734
rect 29748 6458 29776 8026
rect 30208 7954 30236 8588
rect 30392 8548 30420 11494
rect 30300 8520 30420 8548
rect 30196 7948 30248 7954
rect 30196 7890 30248 7896
rect 30300 7342 30328 8520
rect 30378 8392 30434 8401
rect 30378 8327 30380 8336
rect 30432 8327 30434 8336
rect 30380 8298 30432 8304
rect 30484 7478 30512 11766
rect 30472 7472 30524 7478
rect 30472 7414 30524 7420
rect 29920 7336 29972 7342
rect 29918 7304 29920 7313
rect 30288 7336 30340 7342
rect 29972 7304 29974 7313
rect 30288 7278 30340 7284
rect 29918 7239 29974 7248
rect 30470 6760 30526 6769
rect 30470 6695 30472 6704
rect 30524 6695 30526 6704
rect 30472 6666 30524 6672
rect 29736 6452 29788 6458
rect 29736 6394 29788 6400
rect 29368 5160 29420 5166
rect 28630 5128 28686 5137
rect 29368 5102 29420 5108
rect 28630 5063 28686 5072
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 27837 4924 28145 4933
rect 27837 4922 27843 4924
rect 27899 4922 27923 4924
rect 27979 4922 28003 4924
rect 28059 4922 28083 4924
rect 28139 4922 28145 4924
rect 27899 4870 27901 4922
rect 28081 4870 28083 4922
rect 27837 4868 27843 4870
rect 27899 4868 27923 4870
rect 27979 4868 28003 4870
rect 28059 4868 28083 4870
rect 28139 4868 28145 4870
rect 27837 4859 28145 4868
rect 27252 4684 27304 4690
rect 27252 4626 27304 4632
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 8632 4380 8940 4389
rect 8632 4378 8638 4380
rect 8694 4378 8718 4380
rect 8774 4378 8798 4380
rect 8854 4378 8878 4380
rect 8934 4378 8940 4380
rect 8694 4326 8696 4378
rect 8876 4326 8878 4378
rect 8632 4324 8638 4326
rect 8694 4324 8718 4326
rect 8774 4324 8798 4326
rect 8854 4324 8878 4326
rect 8934 4324 8940 4326
rect 8632 4315 8940 4324
rect 16314 4380 16622 4389
rect 16314 4378 16320 4380
rect 16376 4378 16400 4380
rect 16456 4378 16480 4380
rect 16536 4378 16560 4380
rect 16616 4378 16622 4380
rect 16376 4326 16378 4378
rect 16558 4326 16560 4378
rect 16314 4324 16320 4326
rect 16376 4324 16400 4326
rect 16456 4324 16480 4326
rect 16536 4324 16560 4326
rect 16616 4324 16622 4326
rect 16314 4315 16622 4324
rect 23996 4380 24304 4389
rect 23996 4378 24002 4380
rect 24058 4378 24082 4380
rect 24138 4378 24162 4380
rect 24218 4378 24242 4380
rect 24298 4378 24304 4380
rect 24058 4326 24060 4378
rect 24240 4326 24242 4378
rect 23996 4324 24002 4326
rect 24058 4324 24082 4326
rect 24138 4324 24162 4326
rect 24218 4324 24242 4326
rect 24298 4324 24304 4326
rect 23996 4315 24304 4324
rect 1584 4072 1636 4078
rect 1582 4040 1584 4049
rect 1636 4040 1638 4049
rect 1582 3975 1638 3984
rect 28368 3942 28396 4966
rect 28920 4826 28948 4966
rect 28908 4820 28960 4826
rect 28908 4762 28960 4768
rect 30576 4146 30604 14350
rect 30668 13530 30696 15370
rect 30656 13524 30708 13530
rect 30656 13466 30708 13472
rect 30760 13394 30788 15399
rect 30852 13938 30880 18119
rect 30840 13932 30892 13938
rect 30840 13874 30892 13880
rect 30944 13818 30972 18770
rect 31036 14414 31064 18799
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 30852 13790 30972 13818
rect 30748 13388 30800 13394
rect 30748 13330 30800 13336
rect 30852 12434 30880 13790
rect 31128 13682 31156 18838
rect 30760 12406 30880 12434
rect 30944 13654 31156 13682
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30668 5302 30696 12038
rect 30760 8498 30788 12406
rect 30944 10169 30972 13654
rect 31114 13560 31170 13569
rect 31114 13495 31170 13504
rect 31022 10840 31078 10849
rect 31022 10775 31024 10784
rect 31076 10775 31078 10784
rect 31024 10746 31076 10752
rect 30930 10160 30986 10169
rect 30930 10095 30986 10104
rect 31024 10056 31076 10062
rect 31024 9998 31076 10004
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30760 8090 30788 8434
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 31036 6798 31064 9998
rect 31128 6866 31156 13495
rect 31220 13326 31248 20839
rect 31312 20777 31340 20878
rect 31298 20768 31354 20777
rect 31298 20703 31354 20712
rect 31404 20618 31432 23598
rect 31496 22982 31524 24647
rect 31588 24313 31616 30670
rect 31678 30492 31986 30501
rect 31678 30490 31684 30492
rect 31740 30490 31764 30492
rect 31820 30490 31844 30492
rect 31900 30490 31924 30492
rect 31980 30490 31986 30492
rect 31740 30438 31742 30490
rect 31922 30438 31924 30490
rect 31678 30436 31684 30438
rect 31740 30436 31764 30438
rect 31820 30436 31844 30438
rect 31900 30436 31924 30438
rect 31980 30436 31986 30438
rect 31678 30427 31986 30436
rect 31678 29404 31986 29413
rect 31678 29402 31684 29404
rect 31740 29402 31764 29404
rect 31820 29402 31844 29404
rect 31900 29402 31924 29404
rect 31980 29402 31986 29404
rect 31740 29350 31742 29402
rect 31922 29350 31924 29402
rect 31678 29348 31684 29350
rect 31740 29348 31764 29350
rect 31820 29348 31844 29350
rect 31900 29348 31924 29350
rect 31980 29348 31986 29350
rect 31678 29339 31986 29348
rect 31678 28316 31986 28325
rect 31678 28314 31684 28316
rect 31740 28314 31764 28316
rect 31820 28314 31844 28316
rect 31900 28314 31924 28316
rect 31980 28314 31986 28316
rect 31740 28262 31742 28314
rect 31922 28262 31924 28314
rect 31678 28260 31684 28262
rect 31740 28260 31764 28262
rect 31820 28260 31844 28262
rect 31900 28260 31924 28262
rect 31980 28260 31986 28262
rect 31678 28251 31986 28260
rect 31678 27228 31986 27237
rect 31678 27226 31684 27228
rect 31740 27226 31764 27228
rect 31820 27226 31844 27228
rect 31900 27226 31924 27228
rect 31980 27226 31986 27228
rect 31740 27174 31742 27226
rect 31922 27174 31924 27226
rect 31678 27172 31684 27174
rect 31740 27172 31764 27174
rect 31820 27172 31844 27174
rect 31900 27172 31924 27174
rect 31980 27172 31986 27174
rect 31678 27163 31986 27172
rect 31668 27056 31720 27062
rect 31668 26998 31720 27004
rect 31850 27024 31906 27033
rect 31680 26246 31708 26998
rect 31850 26959 31906 26968
rect 31760 26920 31812 26926
rect 31760 26862 31812 26868
rect 31772 26246 31800 26862
rect 31864 26314 31892 26959
rect 32048 26353 32076 31078
rect 32140 26625 32168 31214
rect 32126 26616 32182 26625
rect 32126 26551 32182 26560
rect 32034 26344 32090 26353
rect 31852 26308 31904 26314
rect 32034 26279 32090 26288
rect 31852 26250 31904 26256
rect 31668 26240 31720 26246
rect 31668 26182 31720 26188
rect 31760 26240 31812 26246
rect 32140 26234 32168 26551
rect 31760 26182 31812 26188
rect 32048 26206 32168 26234
rect 31678 26140 31986 26149
rect 31678 26138 31684 26140
rect 31740 26138 31764 26140
rect 31820 26138 31844 26140
rect 31900 26138 31924 26140
rect 31980 26138 31986 26140
rect 31740 26086 31742 26138
rect 31922 26086 31924 26138
rect 31678 26084 31684 26086
rect 31740 26084 31764 26086
rect 31820 26084 31844 26086
rect 31900 26084 31924 26086
rect 31980 26084 31986 26086
rect 31678 26075 31986 26084
rect 31678 25052 31986 25061
rect 31678 25050 31684 25052
rect 31740 25050 31764 25052
rect 31820 25050 31844 25052
rect 31900 25050 31924 25052
rect 31980 25050 31986 25052
rect 31740 24998 31742 25050
rect 31922 24998 31924 25050
rect 31678 24996 31684 24998
rect 31740 24996 31764 24998
rect 31820 24996 31844 24998
rect 31900 24996 31924 24998
rect 31980 24996 31986 24998
rect 31678 24987 31986 24996
rect 32048 24449 32076 26206
rect 32128 26172 32180 26178
rect 32128 26114 32180 26120
rect 32034 24440 32090 24449
rect 32034 24375 32090 24384
rect 31574 24304 31630 24313
rect 31574 24239 31630 24248
rect 31576 24064 31628 24070
rect 31576 24006 31628 24012
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31484 22024 31536 22030
rect 31484 21966 31536 21972
rect 31312 20590 31432 20618
rect 31312 17746 31340 20590
rect 31496 20516 31524 21966
rect 31404 20488 31524 20516
rect 31404 19825 31432 20488
rect 31588 20466 31616 24006
rect 31678 23964 31986 23973
rect 31678 23962 31684 23964
rect 31740 23962 31764 23964
rect 31820 23962 31844 23964
rect 31900 23962 31924 23964
rect 31980 23962 31986 23964
rect 31740 23910 31742 23962
rect 31922 23910 31924 23962
rect 31678 23908 31684 23910
rect 31740 23908 31764 23910
rect 31820 23908 31844 23910
rect 31900 23908 31924 23910
rect 31980 23908 31986 23910
rect 31678 23899 31986 23908
rect 31678 22876 31986 22885
rect 31678 22874 31684 22876
rect 31740 22874 31764 22876
rect 31820 22874 31844 22876
rect 31900 22874 31924 22876
rect 31980 22874 31986 22876
rect 31740 22822 31742 22874
rect 31922 22822 31924 22874
rect 31678 22820 31684 22822
rect 31740 22820 31764 22822
rect 31820 22820 31844 22822
rect 31900 22820 31924 22822
rect 31980 22820 31986 22822
rect 31678 22811 31986 22820
rect 32140 22438 32168 26114
rect 32232 24818 32260 32302
rect 32496 31884 32548 31890
rect 32496 31826 32548 31832
rect 32404 29232 32456 29238
rect 32404 29174 32456 29180
rect 32416 28676 32444 29174
rect 32324 28648 32444 28676
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 31678 21788 31986 21797
rect 31678 21786 31684 21788
rect 31740 21786 31764 21788
rect 31820 21786 31844 21788
rect 31900 21786 31924 21788
rect 31980 21786 31986 21788
rect 31740 21734 31742 21786
rect 31922 21734 31924 21786
rect 31678 21732 31684 21734
rect 31740 21732 31764 21734
rect 31820 21732 31844 21734
rect 31900 21732 31924 21734
rect 31980 21732 31986 21734
rect 31678 21723 31986 21732
rect 31678 20700 31986 20709
rect 31678 20698 31684 20700
rect 31740 20698 31764 20700
rect 31820 20698 31844 20700
rect 31900 20698 31924 20700
rect 31980 20698 31986 20700
rect 31740 20646 31742 20698
rect 31922 20646 31924 20698
rect 31678 20644 31684 20646
rect 31740 20644 31764 20646
rect 31820 20644 31844 20646
rect 31900 20644 31924 20646
rect 31980 20644 31986 20646
rect 31678 20635 31986 20644
rect 32036 20528 32088 20534
rect 32036 20470 32088 20476
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31482 20224 31538 20233
rect 31482 20159 31538 20168
rect 31390 19816 31446 19825
rect 31390 19751 31446 19760
rect 31390 19408 31446 19417
rect 31390 19343 31446 19352
rect 31300 17740 31352 17746
rect 31300 17682 31352 17688
rect 31300 17536 31352 17542
rect 31300 17478 31352 17484
rect 31312 16794 31340 17478
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 31298 16688 31354 16697
rect 31298 16623 31354 16632
rect 31312 16522 31340 16623
rect 31300 16516 31352 16522
rect 31300 16458 31352 16464
rect 31312 16250 31340 16458
rect 31300 16244 31352 16250
rect 31300 16186 31352 16192
rect 31298 16144 31354 16153
rect 31298 16079 31354 16088
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 31220 5370 31248 13262
rect 31312 12850 31340 16079
rect 31404 14618 31432 19343
rect 31392 14612 31444 14618
rect 31392 14554 31444 14560
rect 31496 13938 31524 20159
rect 31576 19916 31628 19922
rect 31576 19858 31628 19864
rect 31588 17610 31616 19858
rect 31678 19612 31986 19621
rect 31678 19610 31684 19612
rect 31740 19610 31764 19612
rect 31820 19610 31844 19612
rect 31900 19610 31924 19612
rect 31980 19610 31986 19612
rect 31740 19558 31742 19610
rect 31922 19558 31924 19610
rect 31678 19556 31684 19558
rect 31740 19556 31764 19558
rect 31820 19556 31844 19558
rect 31900 19556 31924 19558
rect 31980 19556 31986 19558
rect 31678 19547 31986 19556
rect 31668 18760 31720 18766
rect 31666 18728 31668 18737
rect 31720 18728 31722 18737
rect 31666 18663 31722 18672
rect 31678 18524 31986 18533
rect 31678 18522 31684 18524
rect 31740 18522 31764 18524
rect 31820 18522 31844 18524
rect 31900 18522 31924 18524
rect 31980 18522 31986 18524
rect 31740 18470 31742 18522
rect 31922 18470 31924 18522
rect 31678 18468 31684 18470
rect 31740 18468 31764 18470
rect 31820 18468 31844 18470
rect 31900 18468 31924 18470
rect 31980 18468 31986 18470
rect 31678 18459 31986 18468
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31576 17604 31628 17610
rect 31576 17546 31628 17552
rect 31680 17542 31708 18226
rect 32048 17649 32076 20470
rect 32034 17640 32090 17649
rect 32034 17575 32090 17584
rect 31668 17536 31720 17542
rect 31668 17478 31720 17484
rect 31678 17436 31986 17445
rect 31678 17434 31684 17436
rect 31740 17434 31764 17436
rect 31820 17434 31844 17436
rect 31900 17434 31924 17436
rect 31980 17434 31986 17436
rect 31740 17382 31742 17434
rect 31922 17382 31924 17434
rect 31678 17380 31684 17382
rect 31740 17380 31764 17382
rect 31820 17380 31844 17382
rect 31900 17380 31924 17382
rect 31980 17380 31986 17382
rect 31678 17371 31986 17380
rect 32140 17252 32168 22374
rect 32232 19446 32260 23666
rect 32324 19514 32352 28648
rect 32404 28484 32456 28490
rect 32404 28426 32456 28432
rect 32416 23662 32444 28426
rect 32508 25945 32536 31826
rect 32586 30152 32642 30161
rect 32586 30087 32642 30096
rect 32494 25936 32550 25945
rect 32494 25871 32550 25880
rect 32494 25392 32550 25401
rect 32494 25327 32550 25336
rect 32508 24750 32536 25327
rect 32496 24744 32548 24750
rect 32496 24686 32548 24692
rect 32600 24614 32628 30087
rect 32678 29336 32734 29345
rect 32678 29271 32734 29280
rect 32588 24608 32640 24614
rect 32588 24550 32640 24556
rect 32692 24426 32720 29271
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 32770 26752 32826 26761
rect 32770 26687 32826 26696
rect 32508 24398 32720 24426
rect 32404 23656 32456 23662
rect 32404 23598 32456 23604
rect 32402 23352 32458 23361
rect 32402 23287 32458 23296
rect 32312 19508 32364 19514
rect 32312 19450 32364 19456
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 32416 18222 32444 23287
rect 32508 18698 32536 24398
rect 32784 23118 32812 26687
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 32876 22964 32904 29038
rect 32784 22936 32904 22964
rect 32680 22568 32732 22574
rect 32680 22510 32732 22516
rect 32588 20256 32640 20262
rect 32588 20198 32640 20204
rect 32496 18692 32548 18698
rect 32496 18634 32548 18640
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32220 18148 32272 18154
rect 32220 18090 32272 18096
rect 31588 17224 32168 17252
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31390 13424 31446 13433
rect 31390 13359 31446 13368
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31404 12730 31432 13359
rect 31312 12702 31432 12730
rect 31312 12442 31340 12702
rect 31300 12436 31352 12442
rect 31300 12378 31352 12384
rect 31588 12209 31616 17224
rect 32128 17128 32180 17134
rect 31666 17096 31722 17105
rect 32128 17070 32180 17076
rect 31666 17031 31722 17040
rect 31680 16998 31708 17031
rect 31668 16992 31720 16998
rect 31668 16934 31720 16940
rect 32034 16960 32090 16969
rect 32034 16895 32090 16904
rect 31678 16348 31986 16357
rect 31678 16346 31684 16348
rect 31740 16346 31764 16348
rect 31820 16346 31844 16348
rect 31900 16346 31924 16348
rect 31980 16346 31986 16348
rect 31740 16294 31742 16346
rect 31922 16294 31924 16346
rect 31678 16292 31684 16294
rect 31740 16292 31764 16294
rect 31820 16292 31844 16294
rect 31900 16292 31924 16294
rect 31980 16292 31986 16294
rect 31678 16283 31986 16292
rect 31668 16244 31720 16250
rect 31668 16186 31720 16192
rect 31680 15366 31708 16186
rect 31668 15360 31720 15366
rect 31668 15302 31720 15308
rect 31678 15260 31986 15269
rect 31678 15258 31684 15260
rect 31740 15258 31764 15260
rect 31820 15258 31844 15260
rect 31900 15258 31924 15260
rect 31980 15258 31986 15260
rect 31740 15206 31742 15258
rect 31922 15206 31924 15258
rect 31678 15204 31684 15206
rect 31740 15204 31764 15206
rect 31820 15204 31844 15206
rect 31900 15204 31924 15206
rect 31980 15204 31986 15206
rect 31678 15195 31986 15204
rect 31678 14172 31986 14181
rect 31678 14170 31684 14172
rect 31740 14170 31764 14172
rect 31820 14170 31844 14172
rect 31900 14170 31924 14172
rect 31980 14170 31986 14172
rect 31740 14118 31742 14170
rect 31922 14118 31924 14170
rect 31678 14116 31684 14118
rect 31740 14116 31764 14118
rect 31820 14116 31844 14118
rect 31900 14116 31924 14118
rect 31980 14116 31986 14118
rect 31678 14107 31986 14116
rect 31678 13084 31986 13093
rect 31678 13082 31684 13084
rect 31740 13082 31764 13084
rect 31820 13082 31844 13084
rect 31900 13082 31924 13084
rect 31980 13082 31986 13084
rect 31740 13030 31742 13082
rect 31922 13030 31924 13082
rect 31678 13028 31684 13030
rect 31740 13028 31764 13030
rect 31820 13028 31844 13030
rect 31900 13028 31924 13030
rect 31980 13028 31986 13030
rect 31678 13019 31986 13028
rect 31574 12200 31630 12209
rect 31574 12135 31630 12144
rect 31678 11996 31986 12005
rect 31678 11994 31684 11996
rect 31740 11994 31764 11996
rect 31820 11994 31844 11996
rect 31900 11994 31924 11996
rect 31980 11994 31986 11996
rect 31740 11942 31742 11994
rect 31922 11942 31924 11994
rect 31678 11940 31684 11942
rect 31740 11940 31764 11942
rect 31820 11940 31844 11942
rect 31900 11940 31924 11942
rect 31980 11940 31986 11942
rect 31678 11931 31986 11940
rect 31298 11792 31354 11801
rect 31298 11727 31300 11736
rect 31352 11727 31354 11736
rect 31300 11698 31352 11704
rect 31298 11384 31354 11393
rect 31298 11319 31300 11328
rect 31352 11319 31354 11328
rect 31300 11290 31352 11296
rect 31390 10976 31446 10985
rect 31390 10911 31446 10920
rect 31404 10538 31432 10911
rect 31678 10908 31986 10917
rect 31678 10906 31684 10908
rect 31740 10906 31764 10908
rect 31820 10906 31844 10908
rect 31900 10906 31924 10908
rect 31980 10906 31986 10908
rect 31740 10854 31742 10906
rect 31922 10854 31924 10906
rect 31678 10852 31684 10854
rect 31740 10852 31764 10854
rect 31820 10852 31844 10854
rect 31900 10852 31924 10854
rect 31980 10852 31986 10854
rect 31678 10843 31986 10852
rect 31392 10532 31444 10538
rect 31392 10474 31444 10480
rect 31300 10056 31352 10062
rect 31298 10024 31300 10033
rect 31352 10024 31354 10033
rect 31298 9959 31354 9968
rect 31300 9376 31352 9382
rect 31298 9344 31300 9353
rect 31352 9344 31354 9353
rect 31298 9279 31354 9288
rect 31300 8356 31352 8362
rect 31300 8298 31352 8304
rect 31312 7993 31340 8298
rect 31404 8090 31432 10474
rect 31678 9820 31986 9829
rect 31678 9818 31684 9820
rect 31740 9818 31764 9820
rect 31820 9818 31844 9820
rect 31900 9818 31924 9820
rect 31980 9818 31986 9820
rect 31740 9766 31742 9818
rect 31922 9766 31924 9818
rect 31678 9764 31684 9766
rect 31740 9764 31764 9766
rect 31820 9764 31844 9766
rect 31900 9764 31924 9766
rect 31980 9764 31986 9766
rect 31678 9755 31986 9764
rect 31678 8732 31986 8741
rect 31678 8730 31684 8732
rect 31740 8730 31764 8732
rect 31820 8730 31844 8732
rect 31900 8730 31924 8732
rect 31980 8730 31986 8732
rect 31740 8678 31742 8730
rect 31922 8678 31924 8730
rect 31678 8676 31684 8678
rect 31740 8676 31764 8678
rect 31820 8676 31844 8678
rect 31900 8676 31924 8678
rect 31980 8676 31986 8678
rect 31678 8667 31986 8676
rect 32048 8566 32076 16895
rect 32140 15745 32168 17070
rect 32126 15736 32182 15745
rect 32126 15671 32182 15680
rect 32036 8560 32088 8566
rect 32036 8502 32088 8508
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 31298 7984 31354 7993
rect 31298 7919 31354 7928
rect 31678 7644 31986 7653
rect 31678 7642 31684 7644
rect 31740 7642 31764 7644
rect 31820 7642 31844 7644
rect 31900 7642 31924 7644
rect 31980 7642 31986 7644
rect 31740 7590 31742 7642
rect 31922 7590 31924 7642
rect 31678 7588 31684 7590
rect 31740 7588 31764 7590
rect 31820 7588 31844 7590
rect 31900 7588 31924 7590
rect 31980 7588 31986 7590
rect 31678 7579 31986 7588
rect 32140 7546 32168 15671
rect 32232 14385 32260 18090
rect 32312 18080 32364 18086
rect 32312 18022 32364 18028
rect 32218 14376 32274 14385
rect 32218 14311 32274 14320
rect 32324 8022 32352 18022
rect 32416 15026 32444 18158
rect 32404 15020 32456 15026
rect 32404 14962 32456 14968
rect 32600 10742 32628 20198
rect 32692 15881 32720 22510
rect 32784 18358 32812 22936
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 32876 20466 32904 22578
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 32864 20324 32916 20330
rect 32916 20284 32996 20312
rect 32864 20266 32916 20272
rect 32864 20188 32916 20194
rect 32864 20130 32916 20136
rect 32772 18352 32824 18358
rect 32772 18294 32824 18300
rect 32678 15872 32734 15881
rect 32678 15807 32734 15816
rect 32876 12434 32904 20130
rect 32784 12406 32904 12434
rect 32588 10736 32640 10742
rect 32588 10678 32640 10684
rect 32312 8016 32364 8022
rect 32312 7958 32364 7964
rect 32784 7886 32812 12406
rect 32968 10146 32996 20284
rect 32876 10118 32996 10146
rect 32876 9450 32904 10118
rect 32864 9444 32916 9450
rect 32864 9386 32916 9392
rect 32772 7880 32824 7886
rect 32772 7822 32824 7828
rect 32128 7540 32180 7546
rect 32128 7482 32180 7488
rect 31298 7304 31354 7313
rect 31298 7239 31300 7248
rect 31352 7239 31354 7248
rect 31300 7210 31352 7216
rect 31678 6556 31986 6565
rect 31678 6554 31684 6556
rect 31740 6554 31764 6556
rect 31820 6554 31844 6556
rect 31900 6554 31924 6556
rect 31980 6554 31986 6556
rect 31740 6502 31742 6554
rect 31922 6502 31924 6554
rect 31678 6500 31684 6502
rect 31740 6500 31764 6502
rect 31820 6500 31844 6502
rect 31900 6500 31924 6502
rect 31980 6500 31986 6502
rect 31678 6491 31986 6500
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31312 5953 31340 6054
rect 31298 5944 31354 5953
rect 31298 5879 31354 5888
rect 31300 5704 31352 5710
rect 31300 5646 31352 5652
rect 31208 5364 31260 5370
rect 31208 5306 31260 5312
rect 30656 5296 30708 5302
rect 31312 5273 31340 5646
rect 31678 5468 31986 5477
rect 31678 5466 31684 5468
rect 31740 5466 31764 5468
rect 31820 5466 31844 5468
rect 31900 5466 31924 5468
rect 31980 5466 31986 5468
rect 31740 5414 31742 5466
rect 31922 5414 31924 5466
rect 31678 5412 31684 5414
rect 31740 5412 31764 5414
rect 31820 5412 31844 5414
rect 31900 5412 31924 5414
rect 31980 5412 31986 5414
rect 31678 5403 31986 5412
rect 30656 5238 30708 5244
rect 31298 5264 31354 5273
rect 31298 5199 31354 5208
rect 31678 4380 31986 4389
rect 31678 4378 31684 4380
rect 31740 4378 31764 4380
rect 31820 4378 31844 4380
rect 31900 4378 31924 4380
rect 31980 4378 31986 4380
rect 31740 4326 31742 4378
rect 31922 4326 31924 4378
rect 31678 4324 31684 4326
rect 31740 4324 31764 4326
rect 31820 4324 31844 4326
rect 31900 4324 31924 4326
rect 31980 4324 31986 4326
rect 31678 4315 31986 4324
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 30472 3936 30524 3942
rect 31300 3936 31352 3942
rect 30472 3878 30524 3884
rect 31298 3904 31300 3913
rect 31352 3904 31354 3913
rect 4791 3836 5099 3845
rect 4791 3834 4797 3836
rect 4853 3834 4877 3836
rect 4933 3834 4957 3836
rect 5013 3834 5037 3836
rect 5093 3834 5099 3836
rect 4853 3782 4855 3834
rect 5035 3782 5037 3834
rect 4791 3780 4797 3782
rect 4853 3780 4877 3782
rect 4933 3780 4957 3782
rect 5013 3780 5037 3782
rect 5093 3780 5099 3782
rect 4791 3771 5099 3780
rect 12473 3836 12781 3845
rect 12473 3834 12479 3836
rect 12535 3834 12559 3836
rect 12615 3834 12639 3836
rect 12695 3834 12719 3836
rect 12775 3834 12781 3836
rect 12535 3782 12537 3834
rect 12717 3782 12719 3834
rect 12473 3780 12479 3782
rect 12535 3780 12559 3782
rect 12615 3780 12639 3782
rect 12695 3780 12719 3782
rect 12775 3780 12781 3782
rect 12473 3771 12781 3780
rect 20155 3836 20463 3845
rect 20155 3834 20161 3836
rect 20217 3834 20241 3836
rect 20297 3834 20321 3836
rect 20377 3834 20401 3836
rect 20457 3834 20463 3836
rect 20217 3782 20219 3834
rect 20399 3782 20401 3834
rect 20155 3780 20161 3782
rect 20217 3780 20241 3782
rect 20297 3780 20321 3782
rect 20377 3780 20401 3782
rect 20457 3780 20463 3782
rect 20155 3771 20463 3780
rect 27837 3836 28145 3845
rect 27837 3834 27843 3836
rect 27899 3834 27923 3836
rect 27979 3834 28003 3836
rect 28059 3834 28083 3836
rect 28139 3834 28145 3836
rect 27899 3782 27901 3834
rect 28081 3782 28083 3834
rect 27837 3780 27843 3782
rect 27899 3780 27923 3782
rect 27979 3780 28003 3782
rect 28059 3780 28083 3782
rect 28139 3780 28145 3782
rect 27837 3771 28145 3780
rect 30484 3738 30512 3878
rect 31298 3839 31354 3848
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 1584 3528 1636 3534
rect 31300 3528 31352 3534
rect 1584 3470 1636 3476
rect 31298 3496 31300 3505
rect 31352 3496 31354 3505
rect 1596 3233 1624 3470
rect 31298 3431 31354 3440
rect 8632 3292 8940 3301
rect 8632 3290 8638 3292
rect 8694 3290 8718 3292
rect 8774 3290 8798 3292
rect 8854 3290 8878 3292
rect 8934 3290 8940 3292
rect 8694 3238 8696 3290
rect 8876 3238 8878 3290
rect 8632 3236 8638 3238
rect 8694 3236 8718 3238
rect 8774 3236 8798 3238
rect 8854 3236 8878 3238
rect 8934 3236 8940 3238
rect 1582 3224 1638 3233
rect 8632 3227 8940 3236
rect 16314 3292 16622 3301
rect 16314 3290 16320 3292
rect 16376 3290 16400 3292
rect 16456 3290 16480 3292
rect 16536 3290 16560 3292
rect 16616 3290 16622 3292
rect 16376 3238 16378 3290
rect 16558 3238 16560 3290
rect 16314 3236 16320 3238
rect 16376 3236 16400 3238
rect 16456 3236 16480 3238
rect 16536 3236 16560 3238
rect 16616 3236 16622 3238
rect 16314 3227 16622 3236
rect 23996 3292 24304 3301
rect 23996 3290 24002 3292
rect 24058 3290 24082 3292
rect 24138 3290 24162 3292
rect 24218 3290 24242 3292
rect 24298 3290 24304 3292
rect 24058 3238 24060 3290
rect 24240 3238 24242 3290
rect 23996 3236 24002 3238
rect 24058 3236 24082 3238
rect 24138 3236 24162 3238
rect 24218 3236 24242 3238
rect 24298 3236 24304 3238
rect 23996 3227 24304 3236
rect 31678 3292 31986 3301
rect 31678 3290 31684 3292
rect 31740 3290 31764 3292
rect 31820 3290 31844 3292
rect 31900 3290 31924 3292
rect 31980 3290 31986 3292
rect 31740 3238 31742 3290
rect 31922 3238 31924 3290
rect 31678 3236 31684 3238
rect 31740 3236 31764 3238
rect 31820 3236 31844 3238
rect 31900 3236 31924 3238
rect 31980 3236 31986 3238
rect 31678 3227 31986 3236
rect 1582 3159 1638 3168
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 785 1440 2382
rect 1596 1601 1624 2790
rect 4791 2748 5099 2757
rect 4791 2746 4797 2748
rect 4853 2746 4877 2748
rect 4933 2746 4957 2748
rect 5013 2746 5037 2748
rect 5093 2746 5099 2748
rect 4853 2694 4855 2746
rect 5035 2694 5037 2746
rect 4791 2692 4797 2694
rect 4853 2692 4877 2694
rect 4933 2692 4957 2694
rect 5013 2692 5037 2694
rect 5093 2692 5099 2694
rect 4791 2683 5099 2692
rect 12473 2748 12781 2757
rect 12473 2746 12479 2748
rect 12535 2746 12559 2748
rect 12615 2746 12639 2748
rect 12695 2746 12719 2748
rect 12775 2746 12781 2748
rect 12535 2694 12537 2746
rect 12717 2694 12719 2746
rect 12473 2692 12479 2694
rect 12535 2692 12559 2694
rect 12615 2692 12639 2694
rect 12695 2692 12719 2694
rect 12775 2692 12781 2694
rect 12473 2683 12781 2692
rect 20155 2748 20463 2757
rect 20155 2746 20161 2748
rect 20217 2746 20241 2748
rect 20297 2746 20321 2748
rect 20377 2746 20401 2748
rect 20457 2746 20463 2748
rect 20217 2694 20219 2746
rect 20399 2694 20401 2746
rect 20155 2692 20161 2694
rect 20217 2692 20241 2694
rect 20297 2692 20321 2694
rect 20377 2692 20401 2694
rect 20457 2692 20463 2694
rect 20155 2683 20463 2692
rect 27837 2748 28145 2757
rect 27837 2746 27843 2748
rect 27899 2746 27923 2748
rect 27979 2746 28003 2748
rect 28059 2746 28083 2748
rect 28139 2746 28145 2748
rect 27899 2694 27901 2746
rect 28081 2694 28083 2746
rect 27837 2692 27843 2694
rect 27899 2692 27923 2694
rect 27979 2692 28003 2694
rect 28059 2692 28083 2694
rect 28139 2692 28145 2694
rect 27837 2683 28145 2692
rect 8632 2204 8940 2213
rect 8632 2202 8638 2204
rect 8694 2202 8718 2204
rect 8774 2202 8798 2204
rect 8854 2202 8878 2204
rect 8934 2202 8940 2204
rect 8694 2150 8696 2202
rect 8876 2150 8878 2202
rect 8632 2148 8638 2150
rect 8694 2148 8718 2150
rect 8774 2148 8798 2150
rect 8854 2148 8878 2150
rect 8934 2148 8940 2150
rect 8632 2139 8940 2148
rect 16314 2204 16622 2213
rect 16314 2202 16320 2204
rect 16376 2202 16400 2204
rect 16456 2202 16480 2204
rect 16536 2202 16560 2204
rect 16616 2202 16622 2204
rect 16376 2150 16378 2202
rect 16558 2150 16560 2202
rect 16314 2148 16320 2150
rect 16376 2148 16400 2150
rect 16456 2148 16480 2150
rect 16536 2148 16560 2150
rect 16616 2148 16622 2150
rect 16314 2139 16622 2148
rect 23996 2204 24304 2213
rect 23996 2202 24002 2204
rect 24058 2202 24082 2204
rect 24138 2202 24162 2204
rect 24218 2202 24242 2204
rect 24298 2202 24304 2204
rect 24058 2150 24060 2202
rect 24240 2150 24242 2202
rect 23996 2148 24002 2150
rect 24058 2148 24082 2150
rect 24138 2148 24162 2150
rect 24218 2148 24242 2150
rect 24298 2148 24304 2150
rect 23996 2139 24304 2148
rect 31678 2204 31986 2213
rect 31678 2202 31684 2204
rect 31740 2202 31764 2204
rect 31820 2202 31844 2204
rect 31900 2202 31924 2204
rect 31980 2202 31986 2204
rect 31740 2150 31742 2202
rect 31922 2150 31924 2202
rect 31678 2148 31684 2150
rect 31740 2148 31764 2150
rect 31820 2148 31844 2150
rect 31900 2148 31924 2150
rect 31980 2148 31986 2150
rect 31678 2139 31986 2148
rect 1582 1592 1638 1601
rect 1582 1527 1638 1536
rect 1398 776 1454 785
rect 1398 711 1454 720
<< via2 >>
rect 1582 32544 1638 32600
rect 3974 34720 4030 34776
rect 2870 33360 2926 33416
rect 1582 30912 1638 30968
rect 1582 30132 1584 30152
rect 1584 30132 1636 30152
rect 1636 30132 1638 30152
rect 1582 30096 1638 30132
rect 1582 28500 1584 28520
rect 1584 28500 1636 28520
rect 1636 28500 1638 28520
rect 1582 28464 1638 28500
rect 1582 27648 1638 27704
rect 1582 26016 1638 26072
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1582 23604 1584 23624
rect 1584 23604 1636 23624
rect 1636 23604 1638 23624
rect 1582 23568 1638 23604
rect 1582 22752 1638 22808
rect 1582 21120 1638 21176
rect 1582 20340 1584 20360
rect 1584 20340 1636 20360
rect 1636 20340 1638 20360
rect 1582 20304 1638 20340
rect 1582 18708 1584 18728
rect 1584 18708 1636 18728
rect 1636 18708 1638 18728
rect 1582 18672 1638 18708
rect 1582 17856 1638 17912
rect 1582 16224 1638 16280
rect 1582 15444 1584 15464
rect 1584 15444 1636 15464
rect 1636 15444 1638 15464
rect 1582 15408 1638 15444
rect 1582 13812 1584 13832
rect 1584 13812 1636 13832
rect 1636 13812 1638 13832
rect 1582 13776 1638 13812
rect 1582 12960 1638 13016
rect 1582 11328 1638 11384
rect 1582 10548 1584 10568
rect 1584 10548 1636 10568
rect 1636 10548 1638 10568
rect 1582 10512 1638 10548
rect 1582 8916 1584 8936
rect 1584 8916 1636 8936
rect 1636 8916 1638 8936
rect 1582 8880 1638 8916
rect 1582 8064 1638 8120
rect 1582 6432 1638 6488
rect 6642 34856 6698 34912
rect 4342 32408 4398 32464
rect 4797 32122 4853 32124
rect 4877 32122 4933 32124
rect 4957 32122 5013 32124
rect 5037 32122 5093 32124
rect 4797 32070 4843 32122
rect 4843 32070 4853 32122
rect 4877 32070 4907 32122
rect 4907 32070 4919 32122
rect 4919 32070 4933 32122
rect 4957 32070 4971 32122
rect 4971 32070 4983 32122
rect 4983 32070 5013 32122
rect 5037 32070 5047 32122
rect 5047 32070 5093 32122
rect 4797 32068 4853 32070
rect 4877 32068 4933 32070
rect 4957 32068 5013 32070
rect 5037 32068 5093 32070
rect 4797 31034 4853 31036
rect 4877 31034 4933 31036
rect 4957 31034 5013 31036
rect 5037 31034 5093 31036
rect 4797 30982 4843 31034
rect 4843 30982 4853 31034
rect 4877 30982 4907 31034
rect 4907 30982 4919 31034
rect 4919 30982 4933 31034
rect 4957 30982 4971 31034
rect 4971 30982 4983 31034
rect 4983 30982 5013 31034
rect 5037 30982 5047 31034
rect 5047 30982 5093 31034
rect 4797 30980 4853 30982
rect 4877 30980 4933 30982
rect 4957 30980 5013 30982
rect 5037 30980 5093 30982
rect 3974 20304 4030 20360
rect 3882 17720 3938 17776
rect 4797 29946 4853 29948
rect 4877 29946 4933 29948
rect 4957 29946 5013 29948
rect 5037 29946 5093 29948
rect 4797 29894 4843 29946
rect 4843 29894 4853 29946
rect 4877 29894 4907 29946
rect 4907 29894 4919 29946
rect 4919 29894 4933 29946
rect 4957 29894 4971 29946
rect 4971 29894 4983 29946
rect 4983 29894 5013 29946
rect 5037 29894 5047 29946
rect 5047 29894 5093 29946
rect 4797 29892 4853 29894
rect 4877 29892 4933 29894
rect 4957 29892 5013 29894
rect 5037 29892 5093 29894
rect 4526 29688 4582 29744
rect 4066 12688 4122 12744
rect 2686 6160 2742 6216
rect 4797 28858 4853 28860
rect 4877 28858 4933 28860
rect 4957 28858 5013 28860
rect 5037 28858 5093 28860
rect 4797 28806 4843 28858
rect 4843 28806 4853 28858
rect 4877 28806 4907 28858
rect 4907 28806 4919 28858
rect 4919 28806 4933 28858
rect 4957 28806 4971 28858
rect 4971 28806 4983 28858
rect 4983 28806 5013 28858
rect 5037 28806 5047 28858
rect 5047 28806 5093 28858
rect 4797 28804 4853 28806
rect 4877 28804 4933 28806
rect 4957 28804 5013 28806
rect 5037 28804 5093 28806
rect 4797 27770 4853 27772
rect 4877 27770 4933 27772
rect 4957 27770 5013 27772
rect 5037 27770 5093 27772
rect 4797 27718 4843 27770
rect 4843 27718 4853 27770
rect 4877 27718 4907 27770
rect 4907 27718 4919 27770
rect 4919 27718 4933 27770
rect 4957 27718 4971 27770
rect 4971 27718 4983 27770
rect 4983 27718 5013 27770
rect 5037 27718 5047 27770
rect 5047 27718 5093 27770
rect 4797 27716 4853 27718
rect 4877 27716 4933 27718
rect 4957 27716 5013 27718
rect 5037 27716 5093 27718
rect 5262 26832 5318 26888
rect 4797 26682 4853 26684
rect 4877 26682 4933 26684
rect 4957 26682 5013 26684
rect 5037 26682 5093 26684
rect 4797 26630 4843 26682
rect 4843 26630 4853 26682
rect 4877 26630 4907 26682
rect 4907 26630 4919 26682
rect 4919 26630 4933 26682
rect 4957 26630 4971 26682
rect 4971 26630 4983 26682
rect 4983 26630 5013 26682
rect 5037 26630 5047 26682
rect 5047 26630 5093 26682
rect 4797 26628 4853 26630
rect 4877 26628 4933 26630
rect 4957 26628 5013 26630
rect 5037 26628 5093 26630
rect 4797 25594 4853 25596
rect 4877 25594 4933 25596
rect 4957 25594 5013 25596
rect 5037 25594 5093 25596
rect 4797 25542 4843 25594
rect 4843 25542 4853 25594
rect 4877 25542 4907 25594
rect 4907 25542 4919 25594
rect 4919 25542 4933 25594
rect 4957 25542 4971 25594
rect 4971 25542 4983 25594
rect 4983 25542 5013 25594
rect 5037 25542 5047 25594
rect 5047 25542 5093 25594
rect 4797 25540 4853 25542
rect 4877 25540 4933 25542
rect 4957 25540 5013 25542
rect 5037 25540 5093 25542
rect 4797 24506 4853 24508
rect 4877 24506 4933 24508
rect 4957 24506 5013 24508
rect 5037 24506 5093 24508
rect 4797 24454 4843 24506
rect 4843 24454 4853 24506
rect 4877 24454 4907 24506
rect 4907 24454 4919 24506
rect 4919 24454 4933 24506
rect 4957 24454 4971 24506
rect 4971 24454 4983 24506
rect 4983 24454 5013 24506
rect 5037 24454 5047 24506
rect 5047 24454 5093 24506
rect 4797 24452 4853 24454
rect 4877 24452 4933 24454
rect 4957 24452 5013 24454
rect 5037 24452 5093 24454
rect 4797 23418 4853 23420
rect 4877 23418 4933 23420
rect 4957 23418 5013 23420
rect 5037 23418 5093 23420
rect 4797 23366 4843 23418
rect 4843 23366 4853 23418
rect 4877 23366 4907 23418
rect 4907 23366 4919 23418
rect 4919 23366 4933 23418
rect 4957 23366 4971 23418
rect 4971 23366 4983 23418
rect 4983 23366 5013 23418
rect 5037 23366 5047 23418
rect 5047 23366 5093 23418
rect 4797 23364 4853 23366
rect 4877 23364 4933 23366
rect 4957 23364 5013 23366
rect 5037 23364 5093 23366
rect 4797 22330 4853 22332
rect 4877 22330 4933 22332
rect 4957 22330 5013 22332
rect 5037 22330 5093 22332
rect 4797 22278 4843 22330
rect 4843 22278 4853 22330
rect 4877 22278 4907 22330
rect 4907 22278 4919 22330
rect 4919 22278 4933 22330
rect 4957 22278 4971 22330
rect 4971 22278 4983 22330
rect 4983 22278 5013 22330
rect 5037 22278 5047 22330
rect 5047 22278 5093 22330
rect 4797 22276 4853 22278
rect 4877 22276 4933 22278
rect 4957 22276 5013 22278
rect 5037 22276 5093 22278
rect 4710 21972 4712 21992
rect 4712 21972 4764 21992
rect 4764 21972 4766 21992
rect 4710 21936 4766 21972
rect 4797 21242 4853 21244
rect 4877 21242 4933 21244
rect 4957 21242 5013 21244
rect 5037 21242 5093 21244
rect 4797 21190 4843 21242
rect 4843 21190 4853 21242
rect 4877 21190 4907 21242
rect 4907 21190 4919 21242
rect 4919 21190 4933 21242
rect 4957 21190 4971 21242
rect 4971 21190 4983 21242
rect 4983 21190 5013 21242
rect 5037 21190 5047 21242
rect 5047 21190 5093 21242
rect 4797 21188 4853 21190
rect 4877 21188 4933 21190
rect 4957 21188 5013 21190
rect 5037 21188 5093 21190
rect 4797 20154 4853 20156
rect 4877 20154 4933 20156
rect 4957 20154 5013 20156
rect 5037 20154 5093 20156
rect 4797 20102 4843 20154
rect 4843 20102 4853 20154
rect 4877 20102 4907 20154
rect 4907 20102 4919 20154
rect 4919 20102 4933 20154
rect 4957 20102 4971 20154
rect 4971 20102 4983 20154
rect 4983 20102 5013 20154
rect 5037 20102 5047 20154
rect 5047 20102 5093 20154
rect 4797 20100 4853 20102
rect 4877 20100 4933 20102
rect 4957 20100 5013 20102
rect 5037 20100 5093 20102
rect 4797 19066 4853 19068
rect 4877 19066 4933 19068
rect 4957 19066 5013 19068
rect 5037 19066 5093 19068
rect 4797 19014 4843 19066
rect 4843 19014 4853 19066
rect 4877 19014 4907 19066
rect 4907 19014 4919 19066
rect 4919 19014 4933 19066
rect 4957 19014 4971 19066
rect 4971 19014 4983 19066
rect 4983 19014 5013 19066
rect 5037 19014 5047 19066
rect 5047 19014 5093 19066
rect 4797 19012 4853 19014
rect 4877 19012 4933 19014
rect 4957 19012 5013 19014
rect 5037 19012 5093 19014
rect 4797 17978 4853 17980
rect 4877 17978 4933 17980
rect 4957 17978 5013 17980
rect 5037 17978 5093 17980
rect 4797 17926 4843 17978
rect 4843 17926 4853 17978
rect 4877 17926 4907 17978
rect 4907 17926 4919 17978
rect 4919 17926 4933 17978
rect 4957 17926 4971 17978
rect 4971 17926 4983 17978
rect 4983 17926 5013 17978
rect 5037 17926 5047 17978
rect 5047 17926 5093 17978
rect 4797 17924 4853 17926
rect 4877 17924 4933 17926
rect 4957 17924 5013 17926
rect 5037 17924 5093 17926
rect 4797 16890 4853 16892
rect 4877 16890 4933 16892
rect 4957 16890 5013 16892
rect 5037 16890 5093 16892
rect 4797 16838 4843 16890
rect 4843 16838 4853 16890
rect 4877 16838 4907 16890
rect 4907 16838 4919 16890
rect 4919 16838 4933 16890
rect 4957 16838 4971 16890
rect 4971 16838 4983 16890
rect 4983 16838 5013 16890
rect 5037 16838 5047 16890
rect 5047 16838 5093 16890
rect 4797 16836 4853 16838
rect 4877 16836 4933 16838
rect 4957 16836 5013 16838
rect 5037 16836 5093 16838
rect 4797 15802 4853 15804
rect 4877 15802 4933 15804
rect 4957 15802 5013 15804
rect 5037 15802 5093 15804
rect 4797 15750 4843 15802
rect 4843 15750 4853 15802
rect 4877 15750 4907 15802
rect 4907 15750 4919 15802
rect 4919 15750 4933 15802
rect 4957 15750 4971 15802
rect 4971 15750 4983 15802
rect 4983 15750 5013 15802
rect 5037 15750 5047 15802
rect 5047 15750 5093 15802
rect 4797 15748 4853 15750
rect 4877 15748 4933 15750
rect 4957 15748 5013 15750
rect 5037 15748 5093 15750
rect 4797 14714 4853 14716
rect 4877 14714 4933 14716
rect 4957 14714 5013 14716
rect 5037 14714 5093 14716
rect 4797 14662 4843 14714
rect 4843 14662 4853 14714
rect 4877 14662 4907 14714
rect 4907 14662 4919 14714
rect 4919 14662 4933 14714
rect 4957 14662 4971 14714
rect 4971 14662 4983 14714
rect 4983 14662 5013 14714
rect 5037 14662 5047 14714
rect 5047 14662 5093 14714
rect 4797 14660 4853 14662
rect 4877 14660 4933 14662
rect 4957 14660 5013 14662
rect 5037 14660 5093 14662
rect 4797 13626 4853 13628
rect 4877 13626 4933 13628
rect 4957 13626 5013 13628
rect 5037 13626 5093 13628
rect 4797 13574 4843 13626
rect 4843 13574 4853 13626
rect 4877 13574 4907 13626
rect 4907 13574 4919 13626
rect 4919 13574 4933 13626
rect 4957 13574 4971 13626
rect 4971 13574 4983 13626
rect 4983 13574 5013 13626
rect 5037 13574 5047 13626
rect 5047 13574 5093 13626
rect 4797 13572 4853 13574
rect 4877 13572 4933 13574
rect 4957 13572 5013 13574
rect 5037 13572 5093 13574
rect 4797 12538 4853 12540
rect 4877 12538 4933 12540
rect 4957 12538 5013 12540
rect 5037 12538 5093 12540
rect 4797 12486 4843 12538
rect 4843 12486 4853 12538
rect 4877 12486 4907 12538
rect 4907 12486 4919 12538
rect 4919 12486 4933 12538
rect 4957 12486 4971 12538
rect 4971 12486 4983 12538
rect 4983 12486 5013 12538
rect 5037 12486 5047 12538
rect 5047 12486 5093 12538
rect 4797 12484 4853 12486
rect 4877 12484 4933 12486
rect 4957 12484 5013 12486
rect 5037 12484 5093 12486
rect 4797 11450 4853 11452
rect 4877 11450 4933 11452
rect 4957 11450 5013 11452
rect 5037 11450 5093 11452
rect 4797 11398 4843 11450
rect 4843 11398 4853 11450
rect 4877 11398 4907 11450
rect 4907 11398 4919 11450
rect 4919 11398 4933 11450
rect 4957 11398 4971 11450
rect 4971 11398 4983 11450
rect 4983 11398 5013 11450
rect 5037 11398 5047 11450
rect 5047 11398 5093 11450
rect 4797 11396 4853 11398
rect 4877 11396 4933 11398
rect 4957 11396 5013 11398
rect 5037 11396 5093 11398
rect 4797 10362 4853 10364
rect 4877 10362 4933 10364
rect 4957 10362 5013 10364
rect 5037 10362 5093 10364
rect 4797 10310 4843 10362
rect 4843 10310 4853 10362
rect 4877 10310 4907 10362
rect 4907 10310 4919 10362
rect 4919 10310 4933 10362
rect 4957 10310 4971 10362
rect 4971 10310 4983 10362
rect 4983 10310 5013 10362
rect 5037 10310 5047 10362
rect 5047 10310 5093 10362
rect 4797 10308 4853 10310
rect 4877 10308 4933 10310
rect 4957 10308 5013 10310
rect 5037 10308 5093 10310
rect 4797 9274 4853 9276
rect 4877 9274 4933 9276
rect 4957 9274 5013 9276
rect 5037 9274 5093 9276
rect 4797 9222 4843 9274
rect 4843 9222 4853 9274
rect 4877 9222 4907 9274
rect 4907 9222 4919 9274
rect 4919 9222 4933 9274
rect 4957 9222 4971 9274
rect 4971 9222 4983 9274
rect 4983 9222 5013 9274
rect 5037 9222 5047 9274
rect 5047 9222 5093 9274
rect 4797 9220 4853 9222
rect 4877 9220 4933 9222
rect 4957 9220 5013 9222
rect 5037 9220 5093 9222
rect 4797 8186 4853 8188
rect 4877 8186 4933 8188
rect 4957 8186 5013 8188
rect 5037 8186 5093 8188
rect 4797 8134 4843 8186
rect 4843 8134 4853 8186
rect 4877 8134 4907 8186
rect 4907 8134 4919 8186
rect 4919 8134 4933 8186
rect 4957 8134 4971 8186
rect 4971 8134 4983 8186
rect 4983 8134 5013 8186
rect 5037 8134 5047 8186
rect 5047 8134 5093 8186
rect 4797 8132 4853 8134
rect 4877 8132 4933 8134
rect 4957 8132 5013 8134
rect 5037 8132 5093 8134
rect 4797 7098 4853 7100
rect 4877 7098 4933 7100
rect 4957 7098 5013 7100
rect 5037 7098 5093 7100
rect 4797 7046 4843 7098
rect 4843 7046 4853 7098
rect 4877 7046 4907 7098
rect 4907 7046 4919 7098
rect 4919 7046 4933 7098
rect 4957 7046 4971 7098
rect 4971 7046 4983 7098
rect 4983 7046 5013 7098
rect 5037 7046 5047 7098
rect 5047 7046 5093 7098
rect 4797 7044 4853 7046
rect 4877 7044 4933 7046
rect 4957 7044 5013 7046
rect 5037 7044 5093 7046
rect 4797 6010 4853 6012
rect 4877 6010 4933 6012
rect 4957 6010 5013 6012
rect 5037 6010 5093 6012
rect 4797 5958 4843 6010
rect 4843 5958 4853 6010
rect 4877 5958 4907 6010
rect 4907 5958 4919 6010
rect 4919 5958 4933 6010
rect 4957 5958 4971 6010
rect 4971 5958 4983 6010
rect 4983 5958 5013 6010
rect 5037 5958 5047 6010
rect 5047 5958 5093 6010
rect 4797 5956 4853 5958
rect 4877 5956 4933 5958
rect 4957 5956 5013 5958
rect 5037 5956 5093 5958
rect 1582 5652 1584 5672
rect 1584 5652 1636 5672
rect 1636 5652 1638 5672
rect 1582 5616 1638 5652
rect 5998 24676 6054 24712
rect 5998 24656 6000 24676
rect 6000 24656 6052 24676
rect 6052 24656 6054 24676
rect 5814 24112 5870 24168
rect 5446 9560 5502 9616
rect 8638 32666 8694 32668
rect 8718 32666 8774 32668
rect 8798 32666 8854 32668
rect 8878 32666 8934 32668
rect 8638 32614 8684 32666
rect 8684 32614 8694 32666
rect 8718 32614 8748 32666
rect 8748 32614 8760 32666
rect 8760 32614 8774 32666
rect 8798 32614 8812 32666
rect 8812 32614 8824 32666
rect 8824 32614 8854 32666
rect 8878 32614 8888 32666
rect 8888 32614 8934 32666
rect 8638 32612 8694 32614
rect 8718 32612 8774 32614
rect 8798 32612 8854 32614
rect 8878 32612 8934 32614
rect 8638 31578 8694 31580
rect 8718 31578 8774 31580
rect 8798 31578 8854 31580
rect 8878 31578 8934 31580
rect 8638 31526 8684 31578
rect 8684 31526 8694 31578
rect 8718 31526 8748 31578
rect 8748 31526 8760 31578
rect 8760 31526 8774 31578
rect 8798 31526 8812 31578
rect 8812 31526 8824 31578
rect 8824 31526 8854 31578
rect 8878 31526 8888 31578
rect 8888 31526 8934 31578
rect 8638 31524 8694 31526
rect 8718 31524 8774 31526
rect 8798 31524 8854 31526
rect 8878 31524 8934 31526
rect 8206 31320 8262 31376
rect 7378 29144 7434 29200
rect 8022 27396 8078 27432
rect 8022 27376 8024 27396
rect 8024 27376 8076 27396
rect 8076 27376 8078 27396
rect 6918 24248 6974 24304
rect 6826 23432 6882 23488
rect 6734 21800 6790 21856
rect 6550 9560 6606 9616
rect 7838 22072 7894 22128
rect 8638 30490 8694 30492
rect 8718 30490 8774 30492
rect 8798 30490 8854 30492
rect 8878 30490 8934 30492
rect 8638 30438 8684 30490
rect 8684 30438 8694 30490
rect 8718 30438 8748 30490
rect 8748 30438 8760 30490
rect 8760 30438 8774 30490
rect 8798 30438 8812 30490
rect 8812 30438 8824 30490
rect 8824 30438 8854 30490
rect 8878 30438 8888 30490
rect 8888 30438 8934 30490
rect 8638 30436 8694 30438
rect 8718 30436 8774 30438
rect 8798 30436 8854 30438
rect 8878 30436 8934 30438
rect 8638 29402 8694 29404
rect 8718 29402 8774 29404
rect 8798 29402 8854 29404
rect 8878 29402 8934 29404
rect 8638 29350 8684 29402
rect 8684 29350 8694 29402
rect 8718 29350 8748 29402
rect 8748 29350 8760 29402
rect 8760 29350 8774 29402
rect 8798 29350 8812 29402
rect 8812 29350 8824 29402
rect 8824 29350 8854 29402
rect 8878 29350 8888 29402
rect 8888 29350 8934 29402
rect 8638 29348 8694 29350
rect 8718 29348 8774 29350
rect 8798 29348 8854 29350
rect 8878 29348 8934 29350
rect 8638 28314 8694 28316
rect 8718 28314 8774 28316
rect 8798 28314 8854 28316
rect 8878 28314 8934 28316
rect 8638 28262 8684 28314
rect 8684 28262 8694 28314
rect 8718 28262 8748 28314
rect 8748 28262 8760 28314
rect 8760 28262 8774 28314
rect 8798 28262 8812 28314
rect 8812 28262 8824 28314
rect 8824 28262 8854 28314
rect 8878 28262 8888 28314
rect 8888 28262 8934 28314
rect 8638 28260 8694 28262
rect 8718 28260 8774 28262
rect 8798 28260 8854 28262
rect 8878 28260 8934 28262
rect 8206 23024 8262 23080
rect 8206 22772 8262 22808
rect 8206 22752 8208 22772
rect 8208 22752 8260 22772
rect 8260 22752 8262 22772
rect 8206 22344 8262 22400
rect 7746 21120 7802 21176
rect 7654 19352 7710 19408
rect 7286 11192 7342 11248
rect 7378 11056 7434 11112
rect 5722 8336 5778 8392
rect 10046 31728 10102 31784
rect 8638 27226 8694 27228
rect 8718 27226 8774 27228
rect 8798 27226 8854 27228
rect 8878 27226 8934 27228
rect 8638 27174 8684 27226
rect 8684 27174 8694 27226
rect 8718 27174 8748 27226
rect 8748 27174 8760 27226
rect 8760 27174 8774 27226
rect 8798 27174 8812 27226
rect 8812 27174 8824 27226
rect 8824 27174 8854 27226
rect 8878 27174 8888 27226
rect 8888 27174 8934 27226
rect 8638 27172 8694 27174
rect 8718 27172 8774 27174
rect 8798 27172 8854 27174
rect 8878 27172 8934 27174
rect 8390 25744 8446 25800
rect 8638 26138 8694 26140
rect 8718 26138 8774 26140
rect 8798 26138 8854 26140
rect 8878 26138 8934 26140
rect 8638 26086 8684 26138
rect 8684 26086 8694 26138
rect 8718 26086 8748 26138
rect 8748 26086 8760 26138
rect 8760 26086 8774 26138
rect 8798 26086 8812 26138
rect 8812 26086 8824 26138
rect 8824 26086 8854 26138
rect 8878 26086 8888 26138
rect 8888 26086 8934 26138
rect 8638 26084 8694 26086
rect 8718 26084 8774 26086
rect 8798 26084 8854 26086
rect 8878 26084 8934 26086
rect 8638 25050 8694 25052
rect 8718 25050 8774 25052
rect 8798 25050 8854 25052
rect 8878 25050 8934 25052
rect 8638 24998 8684 25050
rect 8684 24998 8694 25050
rect 8718 24998 8748 25050
rect 8748 24998 8760 25050
rect 8760 24998 8774 25050
rect 8798 24998 8812 25050
rect 8812 24998 8824 25050
rect 8824 24998 8854 25050
rect 8878 24998 8888 25050
rect 8888 24998 8934 25050
rect 8638 24996 8694 24998
rect 8718 24996 8774 24998
rect 8798 24996 8854 24998
rect 8878 24996 8934 24998
rect 8298 21004 8354 21040
rect 8298 20984 8300 21004
rect 8300 20984 8352 21004
rect 8352 20984 8354 21004
rect 8638 23962 8694 23964
rect 8718 23962 8774 23964
rect 8798 23962 8854 23964
rect 8878 23962 8934 23964
rect 8638 23910 8684 23962
rect 8684 23910 8694 23962
rect 8718 23910 8748 23962
rect 8748 23910 8760 23962
rect 8760 23910 8774 23962
rect 8798 23910 8812 23962
rect 8812 23910 8824 23962
rect 8824 23910 8854 23962
rect 8878 23910 8888 23962
rect 8888 23910 8934 23962
rect 8638 23908 8694 23910
rect 8718 23908 8774 23910
rect 8798 23908 8854 23910
rect 8878 23908 8934 23910
rect 8482 23316 8538 23352
rect 8482 23296 8484 23316
rect 8484 23296 8536 23316
rect 8536 23296 8538 23316
rect 8850 23160 8906 23216
rect 8638 22874 8694 22876
rect 8718 22874 8774 22876
rect 8798 22874 8854 22876
rect 8878 22874 8934 22876
rect 8638 22822 8684 22874
rect 8684 22822 8694 22874
rect 8718 22822 8748 22874
rect 8748 22822 8760 22874
rect 8760 22822 8774 22874
rect 8798 22822 8812 22874
rect 8812 22822 8824 22874
rect 8824 22822 8854 22874
rect 8878 22822 8888 22874
rect 8888 22822 8934 22874
rect 8638 22820 8694 22822
rect 8718 22820 8774 22822
rect 8798 22820 8854 22822
rect 8878 22820 8934 22822
rect 8758 21936 8814 21992
rect 9954 30096 10010 30152
rect 9954 29028 10010 29064
rect 12070 33904 12126 33960
rect 9954 29008 9956 29028
rect 9956 29008 10008 29028
rect 10008 29008 10010 29028
rect 10322 27920 10378 27976
rect 9310 26324 9312 26344
rect 9312 26324 9364 26344
rect 9364 26324 9366 26344
rect 9310 26288 9366 26324
rect 9218 24792 9274 24848
rect 9494 25336 9550 25392
rect 8390 20576 8446 20632
rect 8390 9424 8446 9480
rect 9034 21800 9090 21856
rect 8638 21786 8694 21788
rect 8718 21786 8774 21788
rect 8798 21786 8854 21788
rect 8878 21786 8934 21788
rect 8638 21734 8684 21786
rect 8684 21734 8694 21786
rect 8718 21734 8748 21786
rect 8748 21734 8760 21786
rect 8760 21734 8774 21786
rect 8798 21734 8812 21786
rect 8812 21734 8824 21786
rect 8824 21734 8854 21786
rect 8878 21734 8888 21786
rect 8888 21734 8934 21786
rect 8638 21732 8694 21734
rect 8718 21732 8774 21734
rect 8798 21732 8854 21734
rect 8878 21732 8934 21734
rect 8638 20698 8694 20700
rect 8718 20698 8774 20700
rect 8798 20698 8854 20700
rect 8878 20698 8934 20700
rect 8638 20646 8684 20698
rect 8684 20646 8694 20698
rect 8718 20646 8748 20698
rect 8748 20646 8760 20698
rect 8760 20646 8774 20698
rect 8798 20646 8812 20698
rect 8812 20646 8824 20698
rect 8824 20646 8854 20698
rect 8878 20646 8888 20698
rect 8888 20646 8934 20698
rect 8638 20644 8694 20646
rect 8718 20644 8774 20646
rect 8798 20644 8854 20646
rect 8878 20644 8934 20646
rect 9034 20576 9090 20632
rect 8638 19610 8694 19612
rect 8718 19610 8774 19612
rect 8798 19610 8854 19612
rect 8878 19610 8934 19612
rect 8638 19558 8684 19610
rect 8684 19558 8694 19610
rect 8718 19558 8748 19610
rect 8748 19558 8760 19610
rect 8760 19558 8774 19610
rect 8798 19558 8812 19610
rect 8812 19558 8824 19610
rect 8824 19558 8854 19610
rect 8878 19558 8888 19610
rect 8888 19558 8934 19610
rect 8638 19556 8694 19558
rect 8718 19556 8774 19558
rect 8798 19556 8854 19558
rect 8878 19556 8934 19558
rect 8638 18522 8694 18524
rect 8718 18522 8774 18524
rect 8798 18522 8854 18524
rect 8878 18522 8934 18524
rect 8638 18470 8684 18522
rect 8684 18470 8694 18522
rect 8718 18470 8748 18522
rect 8748 18470 8760 18522
rect 8760 18470 8774 18522
rect 8798 18470 8812 18522
rect 8812 18470 8824 18522
rect 8824 18470 8854 18522
rect 8878 18470 8888 18522
rect 8888 18470 8934 18522
rect 8638 18468 8694 18470
rect 8718 18468 8774 18470
rect 8798 18468 8854 18470
rect 8878 18468 8934 18470
rect 8638 17434 8694 17436
rect 8718 17434 8774 17436
rect 8798 17434 8854 17436
rect 8878 17434 8934 17436
rect 8638 17382 8684 17434
rect 8684 17382 8694 17434
rect 8718 17382 8748 17434
rect 8748 17382 8760 17434
rect 8760 17382 8774 17434
rect 8798 17382 8812 17434
rect 8812 17382 8824 17434
rect 8824 17382 8854 17434
rect 8878 17382 8888 17434
rect 8888 17382 8934 17434
rect 8638 17380 8694 17382
rect 8718 17380 8774 17382
rect 8798 17380 8854 17382
rect 8878 17380 8934 17382
rect 8638 16346 8694 16348
rect 8718 16346 8774 16348
rect 8798 16346 8854 16348
rect 8878 16346 8934 16348
rect 8638 16294 8684 16346
rect 8684 16294 8694 16346
rect 8718 16294 8748 16346
rect 8748 16294 8760 16346
rect 8760 16294 8774 16346
rect 8798 16294 8812 16346
rect 8812 16294 8824 16346
rect 8824 16294 8854 16346
rect 8878 16294 8888 16346
rect 8888 16294 8934 16346
rect 8638 16292 8694 16294
rect 8718 16292 8774 16294
rect 8798 16292 8854 16294
rect 8878 16292 8934 16294
rect 8638 15258 8694 15260
rect 8718 15258 8774 15260
rect 8798 15258 8854 15260
rect 8878 15258 8934 15260
rect 8638 15206 8684 15258
rect 8684 15206 8694 15258
rect 8718 15206 8748 15258
rect 8748 15206 8760 15258
rect 8760 15206 8774 15258
rect 8798 15206 8812 15258
rect 8812 15206 8824 15258
rect 8824 15206 8854 15258
rect 8878 15206 8888 15258
rect 8888 15206 8934 15258
rect 8638 15204 8694 15206
rect 8718 15204 8774 15206
rect 8798 15204 8854 15206
rect 8878 15204 8934 15206
rect 8638 14170 8694 14172
rect 8718 14170 8774 14172
rect 8798 14170 8854 14172
rect 8878 14170 8934 14172
rect 8638 14118 8684 14170
rect 8684 14118 8694 14170
rect 8718 14118 8748 14170
rect 8748 14118 8760 14170
rect 8760 14118 8774 14170
rect 8798 14118 8812 14170
rect 8812 14118 8824 14170
rect 8824 14118 8854 14170
rect 8878 14118 8888 14170
rect 8888 14118 8934 14170
rect 8638 14116 8694 14118
rect 8718 14116 8774 14118
rect 8798 14116 8854 14118
rect 8878 14116 8934 14118
rect 8638 13082 8694 13084
rect 8718 13082 8774 13084
rect 8798 13082 8854 13084
rect 8878 13082 8934 13084
rect 8638 13030 8684 13082
rect 8684 13030 8694 13082
rect 8718 13030 8748 13082
rect 8748 13030 8760 13082
rect 8760 13030 8774 13082
rect 8798 13030 8812 13082
rect 8812 13030 8824 13082
rect 8824 13030 8854 13082
rect 8878 13030 8888 13082
rect 8888 13030 8934 13082
rect 8638 13028 8694 13030
rect 8718 13028 8774 13030
rect 8798 13028 8854 13030
rect 8878 13028 8934 13030
rect 8638 11994 8694 11996
rect 8718 11994 8774 11996
rect 8798 11994 8854 11996
rect 8878 11994 8934 11996
rect 8638 11942 8684 11994
rect 8684 11942 8694 11994
rect 8718 11942 8748 11994
rect 8748 11942 8760 11994
rect 8760 11942 8774 11994
rect 8798 11942 8812 11994
rect 8812 11942 8824 11994
rect 8824 11942 8854 11994
rect 8878 11942 8888 11994
rect 8888 11942 8934 11994
rect 8638 11940 8694 11942
rect 8718 11940 8774 11942
rect 8798 11940 8854 11942
rect 8878 11940 8934 11942
rect 8638 10906 8694 10908
rect 8718 10906 8774 10908
rect 8798 10906 8854 10908
rect 8878 10906 8934 10908
rect 8638 10854 8684 10906
rect 8684 10854 8694 10906
rect 8718 10854 8748 10906
rect 8748 10854 8760 10906
rect 8760 10854 8774 10906
rect 8798 10854 8812 10906
rect 8812 10854 8824 10906
rect 8824 10854 8854 10906
rect 8878 10854 8888 10906
rect 8888 10854 8934 10906
rect 8638 10852 8694 10854
rect 8718 10852 8774 10854
rect 8798 10852 8854 10854
rect 8878 10852 8934 10854
rect 8638 9818 8694 9820
rect 8718 9818 8774 9820
rect 8798 9818 8854 9820
rect 8878 9818 8934 9820
rect 8638 9766 8684 9818
rect 8684 9766 8694 9818
rect 8718 9766 8748 9818
rect 8748 9766 8760 9818
rect 8760 9766 8774 9818
rect 8798 9766 8812 9818
rect 8812 9766 8824 9818
rect 8824 9766 8854 9818
rect 8878 9766 8888 9818
rect 8888 9766 8934 9818
rect 8638 9764 8694 9766
rect 8718 9764 8774 9766
rect 8798 9764 8854 9766
rect 8878 9764 8934 9766
rect 8638 8730 8694 8732
rect 8718 8730 8774 8732
rect 8798 8730 8854 8732
rect 8878 8730 8934 8732
rect 8638 8678 8684 8730
rect 8684 8678 8694 8730
rect 8718 8678 8748 8730
rect 8748 8678 8760 8730
rect 8760 8678 8774 8730
rect 8798 8678 8812 8730
rect 8812 8678 8824 8730
rect 8824 8678 8854 8730
rect 8878 8678 8888 8730
rect 8888 8678 8934 8730
rect 8638 8676 8694 8678
rect 8718 8676 8774 8678
rect 8798 8676 8854 8678
rect 8878 8676 8934 8678
rect 9678 26152 9734 26208
rect 9678 23704 9734 23760
rect 9770 23568 9826 23624
rect 10230 25064 10286 25120
rect 11426 30796 11482 30832
rect 11426 30776 11428 30796
rect 11428 30776 11480 30796
rect 11480 30776 11482 30796
rect 10506 22636 10562 22672
rect 10506 22616 10508 22636
rect 10508 22616 10560 22636
rect 10560 22616 10562 22636
rect 10598 22480 10654 22536
rect 9770 21548 9826 21584
rect 9770 21528 9772 21548
rect 9772 21528 9824 21548
rect 9824 21528 9826 21548
rect 9678 21428 9680 21448
rect 9680 21428 9732 21448
rect 9732 21428 9734 21448
rect 9678 21392 9734 21428
rect 9678 20324 9734 20360
rect 9678 20304 9680 20324
rect 9680 20304 9732 20324
rect 9732 20304 9734 20324
rect 9678 19080 9734 19136
rect 10046 18420 10102 18456
rect 10046 18400 10048 18420
rect 10048 18400 10100 18420
rect 10100 18400 10102 18420
rect 10414 20440 10470 20496
rect 10598 20032 10654 20088
rect 10598 18400 10654 18456
rect 10414 17040 10470 17096
rect 10506 16940 10508 16960
rect 10508 16940 10560 16960
rect 10560 16940 10562 16960
rect 10506 16904 10562 16940
rect 10322 11736 10378 11792
rect 11058 23296 11114 23352
rect 11242 22752 11298 22808
rect 11150 22072 11206 22128
rect 11518 27104 11574 27160
rect 12479 32122 12535 32124
rect 12559 32122 12615 32124
rect 12639 32122 12695 32124
rect 12719 32122 12775 32124
rect 12479 32070 12525 32122
rect 12525 32070 12535 32122
rect 12559 32070 12589 32122
rect 12589 32070 12601 32122
rect 12601 32070 12615 32122
rect 12639 32070 12653 32122
rect 12653 32070 12665 32122
rect 12665 32070 12695 32122
rect 12719 32070 12729 32122
rect 12729 32070 12775 32122
rect 12479 32068 12535 32070
rect 12559 32068 12615 32070
rect 12639 32068 12695 32070
rect 12719 32068 12775 32070
rect 12479 31034 12535 31036
rect 12559 31034 12615 31036
rect 12639 31034 12695 31036
rect 12719 31034 12775 31036
rect 12479 30982 12525 31034
rect 12525 30982 12535 31034
rect 12559 30982 12589 31034
rect 12589 30982 12601 31034
rect 12601 30982 12615 31034
rect 12639 30982 12653 31034
rect 12653 30982 12665 31034
rect 12665 30982 12695 31034
rect 12719 30982 12729 31034
rect 12729 30982 12775 31034
rect 12479 30980 12535 30982
rect 12559 30980 12615 30982
rect 12639 30980 12695 30982
rect 12719 30980 12775 30982
rect 12806 30368 12862 30424
rect 14830 34448 14886 34504
rect 13266 34176 13322 34232
rect 13174 31184 13230 31240
rect 13358 30368 13414 30424
rect 13358 30232 13414 30288
rect 12479 29946 12535 29948
rect 12559 29946 12615 29948
rect 12639 29946 12695 29948
rect 12719 29946 12775 29948
rect 12479 29894 12525 29946
rect 12525 29894 12535 29946
rect 12559 29894 12589 29946
rect 12589 29894 12601 29946
rect 12601 29894 12615 29946
rect 12639 29894 12653 29946
rect 12653 29894 12665 29946
rect 12665 29894 12695 29946
rect 12719 29894 12729 29946
rect 12729 29894 12775 29946
rect 12479 29892 12535 29894
rect 12559 29892 12615 29894
rect 12639 29892 12695 29894
rect 12719 29892 12775 29894
rect 12806 29688 12862 29744
rect 11426 24112 11482 24168
rect 11426 22652 11428 22672
rect 11428 22652 11480 22672
rect 11480 22652 11482 22672
rect 11426 22616 11482 22652
rect 10874 20712 10930 20768
rect 10782 19488 10838 19544
rect 11426 20712 11482 20768
rect 11058 19896 11114 19952
rect 10966 19216 11022 19272
rect 11242 20168 11298 20224
rect 11610 23432 11666 23488
rect 11702 22616 11758 22672
rect 11886 23840 11942 23896
rect 12479 28858 12535 28860
rect 12559 28858 12615 28860
rect 12639 28858 12695 28860
rect 12719 28858 12775 28860
rect 12479 28806 12525 28858
rect 12525 28806 12535 28858
rect 12559 28806 12589 28858
rect 12589 28806 12601 28858
rect 12601 28806 12615 28858
rect 12639 28806 12653 28858
rect 12653 28806 12665 28858
rect 12665 28806 12695 28858
rect 12719 28806 12729 28858
rect 12729 28806 12775 28858
rect 12479 28804 12535 28806
rect 12559 28804 12615 28806
rect 12639 28804 12695 28806
rect 12719 28804 12775 28806
rect 12898 29144 12954 29200
rect 12479 27770 12535 27772
rect 12559 27770 12615 27772
rect 12639 27770 12695 27772
rect 12719 27770 12775 27772
rect 12479 27718 12525 27770
rect 12525 27718 12535 27770
rect 12559 27718 12589 27770
rect 12589 27718 12601 27770
rect 12601 27718 12615 27770
rect 12639 27718 12653 27770
rect 12653 27718 12665 27770
rect 12665 27718 12695 27770
rect 12719 27718 12729 27770
rect 12729 27718 12775 27770
rect 12479 27716 12535 27718
rect 12559 27716 12615 27718
rect 12639 27716 12695 27718
rect 12719 27716 12775 27718
rect 12254 27240 12310 27296
rect 12479 26682 12535 26684
rect 12559 26682 12615 26684
rect 12639 26682 12695 26684
rect 12719 26682 12775 26684
rect 12479 26630 12525 26682
rect 12525 26630 12535 26682
rect 12559 26630 12589 26682
rect 12589 26630 12601 26682
rect 12601 26630 12615 26682
rect 12639 26630 12653 26682
rect 12653 26630 12665 26682
rect 12665 26630 12695 26682
rect 12719 26630 12729 26682
rect 12729 26630 12775 26682
rect 12479 26628 12535 26630
rect 12559 26628 12615 26630
rect 12639 26628 12695 26630
rect 12719 26628 12775 26630
rect 12162 25200 12218 25256
rect 12346 26016 12402 26072
rect 12806 26424 12862 26480
rect 12162 24248 12218 24304
rect 12070 23704 12126 23760
rect 12162 23568 12218 23624
rect 11886 22888 11942 22944
rect 11794 19488 11850 19544
rect 11794 18808 11850 18864
rect 11610 18128 11666 18184
rect 11150 16496 11206 16552
rect 10690 12280 10746 12336
rect 11610 16088 11666 16144
rect 12162 22924 12164 22944
rect 12164 22924 12216 22944
rect 12216 22924 12218 22944
rect 11978 22228 12034 22264
rect 11978 22208 11980 22228
rect 11980 22208 12032 22228
rect 12032 22208 12034 22228
rect 12162 22888 12218 22924
rect 12162 22344 12218 22400
rect 12479 25594 12535 25596
rect 12559 25594 12615 25596
rect 12639 25594 12695 25596
rect 12719 25594 12775 25596
rect 12479 25542 12525 25594
rect 12525 25542 12535 25594
rect 12559 25542 12589 25594
rect 12589 25542 12601 25594
rect 12601 25542 12615 25594
rect 12639 25542 12653 25594
rect 12653 25542 12665 25594
rect 12665 25542 12695 25594
rect 12719 25542 12729 25594
rect 12729 25542 12775 25594
rect 12479 25540 12535 25542
rect 12559 25540 12615 25542
rect 12639 25540 12695 25542
rect 12719 25540 12775 25542
rect 12898 25472 12954 25528
rect 12806 24928 12862 24984
rect 13358 29008 13414 29064
rect 12479 24506 12535 24508
rect 12559 24506 12615 24508
rect 12639 24506 12695 24508
rect 12719 24506 12775 24508
rect 12479 24454 12525 24506
rect 12525 24454 12535 24506
rect 12559 24454 12589 24506
rect 12589 24454 12601 24506
rect 12601 24454 12615 24506
rect 12639 24454 12653 24506
rect 12653 24454 12665 24506
rect 12665 24454 12695 24506
rect 12719 24454 12729 24506
rect 12729 24454 12775 24506
rect 12479 24452 12535 24454
rect 12559 24452 12615 24454
rect 12639 24452 12695 24454
rect 12719 24452 12775 24454
rect 12438 24248 12494 24304
rect 12346 23724 12402 23760
rect 12346 23704 12348 23724
rect 12348 23704 12400 23724
rect 12400 23704 12402 23724
rect 12346 23432 12402 23488
rect 12479 23418 12535 23420
rect 12559 23418 12615 23420
rect 12639 23418 12695 23420
rect 12719 23418 12775 23420
rect 12479 23366 12525 23418
rect 12525 23366 12535 23418
rect 12559 23366 12589 23418
rect 12589 23366 12601 23418
rect 12601 23366 12615 23418
rect 12639 23366 12653 23418
rect 12653 23366 12665 23418
rect 12665 23366 12695 23418
rect 12719 23366 12729 23418
rect 12729 23366 12775 23418
rect 12479 23364 12535 23366
rect 12559 23364 12615 23366
rect 12639 23364 12695 23366
rect 12719 23364 12775 23366
rect 12714 23160 12770 23216
rect 12622 22888 12678 22944
rect 12806 23060 12808 23080
rect 12808 23060 12860 23080
rect 12860 23060 12862 23080
rect 12806 23024 12862 23060
rect 12990 23568 13046 23624
rect 13266 24928 13322 24984
rect 13542 31340 13598 31376
rect 13542 31320 13544 31340
rect 13544 31320 13596 31340
rect 13596 31320 13598 31340
rect 14370 32272 14426 32328
rect 17314 34312 17370 34368
rect 25318 34584 25374 34640
rect 24950 34448 25006 34504
rect 16320 32666 16376 32668
rect 16400 32666 16456 32668
rect 16480 32666 16536 32668
rect 16560 32666 16616 32668
rect 16320 32614 16366 32666
rect 16366 32614 16376 32666
rect 16400 32614 16430 32666
rect 16430 32614 16442 32666
rect 16442 32614 16456 32666
rect 16480 32614 16494 32666
rect 16494 32614 16506 32666
rect 16506 32614 16536 32666
rect 16560 32614 16570 32666
rect 16570 32614 16616 32666
rect 16320 32612 16376 32614
rect 16400 32612 16456 32614
rect 16480 32612 16536 32614
rect 16560 32612 16616 32614
rect 13634 26016 13690 26072
rect 13818 28756 13874 28792
rect 13818 28736 13820 28756
rect 13820 28736 13872 28756
rect 13872 28736 13874 28756
rect 13818 26968 13874 27024
rect 13266 24248 13322 24304
rect 13634 25744 13690 25800
rect 13726 25472 13782 25528
rect 13542 24112 13598 24168
rect 13266 23432 13322 23488
rect 13358 23296 13414 23352
rect 13542 23296 13598 23352
rect 12479 22330 12535 22332
rect 12559 22330 12615 22332
rect 12639 22330 12695 22332
rect 12719 22330 12775 22332
rect 12479 22278 12525 22330
rect 12525 22278 12535 22330
rect 12559 22278 12589 22330
rect 12589 22278 12601 22330
rect 12601 22278 12615 22330
rect 12639 22278 12653 22330
rect 12653 22278 12665 22330
rect 12665 22278 12695 22330
rect 12719 22278 12729 22330
rect 12729 22278 12775 22330
rect 12479 22276 12535 22278
rect 12559 22276 12615 22278
rect 12639 22276 12695 22278
rect 12719 22276 12775 22278
rect 12898 22208 12954 22264
rect 12622 21800 12678 21856
rect 12254 21664 12310 21720
rect 12438 21664 12494 21720
rect 12346 21392 12402 21448
rect 12806 22072 12862 22128
rect 12530 21412 12586 21448
rect 12530 21392 12532 21412
rect 12532 21392 12584 21412
rect 12584 21392 12586 21412
rect 12479 21242 12535 21244
rect 12559 21242 12615 21244
rect 12639 21242 12695 21244
rect 12719 21242 12775 21244
rect 12479 21190 12525 21242
rect 12525 21190 12535 21242
rect 12559 21190 12589 21242
rect 12589 21190 12601 21242
rect 12601 21190 12615 21242
rect 12639 21190 12653 21242
rect 12653 21190 12665 21242
rect 12665 21190 12695 21242
rect 12719 21190 12729 21242
rect 12729 21190 12775 21242
rect 12479 21188 12535 21190
rect 12559 21188 12615 21190
rect 12639 21188 12695 21190
rect 12719 21188 12775 21190
rect 12346 21120 12402 21176
rect 12070 20984 12126 21040
rect 12530 20884 12532 20904
rect 12532 20884 12584 20904
rect 12584 20884 12586 20904
rect 12530 20848 12586 20884
rect 12070 20712 12126 20768
rect 12346 20712 12402 20768
rect 12346 20576 12402 20632
rect 12254 20032 12310 20088
rect 12070 19624 12126 19680
rect 13450 23160 13506 23216
rect 13910 26152 13966 26208
rect 13910 24792 13966 24848
rect 13910 24148 13912 24168
rect 13912 24148 13964 24168
rect 13964 24148 13966 24168
rect 13910 24112 13966 24148
rect 14186 27412 14188 27432
rect 14188 27412 14240 27432
rect 14240 27412 14242 27432
rect 14186 27376 14242 27412
rect 14186 26696 14242 26752
rect 14094 25064 14150 25120
rect 14094 24248 14150 24304
rect 14002 23976 14058 24032
rect 13910 23296 13966 23352
rect 13450 22480 13506 22536
rect 13266 22344 13322 22400
rect 13726 22888 13782 22944
rect 13726 22208 13782 22264
rect 13358 21528 13414 21584
rect 13634 21120 13690 21176
rect 13266 20712 13322 20768
rect 12898 20596 12954 20632
rect 12898 20576 12900 20596
rect 12900 20576 12952 20596
rect 12952 20576 12954 20596
rect 12479 20154 12535 20156
rect 12559 20154 12615 20156
rect 12639 20154 12695 20156
rect 12719 20154 12775 20156
rect 12479 20102 12525 20154
rect 12525 20102 12535 20154
rect 12559 20102 12589 20154
rect 12589 20102 12601 20154
rect 12601 20102 12615 20154
rect 12639 20102 12653 20154
rect 12653 20102 12665 20154
rect 12665 20102 12695 20154
rect 12719 20102 12729 20154
rect 12729 20102 12775 20154
rect 12479 20100 12535 20102
rect 12559 20100 12615 20102
rect 12639 20100 12695 20102
rect 12719 20100 12775 20102
rect 12530 19488 12586 19544
rect 12806 19760 12862 19816
rect 12990 19488 13046 19544
rect 12806 19372 12862 19408
rect 12806 19352 12808 19372
rect 12808 19352 12860 19372
rect 12860 19352 12862 19372
rect 12346 19080 12402 19136
rect 12479 19066 12535 19068
rect 12559 19066 12615 19068
rect 12639 19066 12695 19068
rect 12719 19066 12775 19068
rect 12479 19014 12525 19066
rect 12525 19014 12535 19066
rect 12559 19014 12589 19066
rect 12589 19014 12601 19066
rect 12601 19014 12615 19066
rect 12639 19014 12653 19066
rect 12653 19014 12665 19066
rect 12665 19014 12695 19066
rect 12719 19014 12729 19066
rect 12729 19014 12775 19066
rect 12479 19012 12535 19014
rect 12559 19012 12615 19014
rect 12639 19012 12695 19014
rect 12719 19012 12775 19014
rect 12479 17978 12535 17980
rect 12559 17978 12615 17980
rect 12639 17978 12695 17980
rect 12719 17978 12775 17980
rect 12479 17926 12525 17978
rect 12525 17926 12535 17978
rect 12559 17926 12589 17978
rect 12589 17926 12601 17978
rect 12601 17926 12615 17978
rect 12639 17926 12653 17978
rect 12653 17926 12665 17978
rect 12665 17926 12695 17978
rect 12719 17926 12729 17978
rect 12729 17926 12775 17978
rect 12479 17924 12535 17926
rect 12559 17924 12615 17926
rect 12639 17924 12695 17926
rect 12719 17924 12775 17926
rect 13266 19352 13322 19408
rect 13450 20712 13506 20768
rect 13542 20576 13598 20632
rect 13450 19488 13506 19544
rect 13450 19216 13506 19272
rect 14738 31084 14740 31104
rect 14740 31084 14792 31104
rect 14792 31084 14794 31104
rect 14738 31048 14794 31084
rect 14370 29280 14426 29336
rect 14462 29008 14518 29064
rect 14554 28056 14610 28112
rect 14462 25880 14518 25936
rect 14278 25472 14334 25528
rect 14462 25236 14464 25256
rect 14464 25236 14516 25256
rect 14516 25236 14518 25256
rect 14462 25200 14518 25236
rect 14094 23296 14150 23352
rect 14922 30912 14978 30968
rect 15382 30096 15438 30152
rect 14922 27376 14978 27432
rect 14738 25472 14794 25528
rect 15106 26308 15162 26344
rect 15106 26288 15108 26308
rect 15108 26288 15160 26308
rect 15160 26288 15162 26308
rect 15474 28600 15530 28656
rect 15382 27512 15438 27568
rect 14922 24928 14978 24984
rect 14738 24792 14794 24848
rect 14830 24520 14886 24576
rect 14738 24404 14794 24440
rect 14738 24384 14740 24404
rect 14740 24384 14792 24404
rect 14792 24384 14794 24404
rect 14646 24112 14702 24168
rect 14554 23840 14610 23896
rect 14370 22072 14426 22128
rect 14922 23704 14978 23760
rect 15290 26016 15346 26072
rect 15290 25900 15346 25936
rect 15290 25880 15292 25900
rect 15292 25880 15344 25900
rect 15344 25880 15346 25900
rect 14922 23432 14978 23488
rect 14830 23316 14886 23352
rect 14830 23296 14832 23316
rect 14832 23296 14884 23316
rect 14884 23296 14886 23316
rect 14646 22752 14702 22808
rect 14646 21800 14702 21856
rect 14186 21664 14242 21720
rect 13818 20032 13874 20088
rect 14002 19624 14058 19680
rect 14462 21528 14518 21584
rect 14738 21392 14794 21448
rect 13174 18264 13230 18320
rect 13266 17856 13322 17912
rect 12898 17448 12954 17504
rect 12622 17312 12678 17368
rect 13082 17312 13138 17368
rect 12162 16496 12218 16552
rect 12479 16890 12535 16892
rect 12559 16890 12615 16892
rect 12639 16890 12695 16892
rect 12719 16890 12775 16892
rect 12479 16838 12525 16890
rect 12525 16838 12535 16890
rect 12559 16838 12589 16890
rect 12589 16838 12601 16890
rect 12601 16838 12615 16890
rect 12639 16838 12653 16890
rect 12653 16838 12665 16890
rect 12665 16838 12695 16890
rect 12719 16838 12729 16890
rect 12729 16838 12775 16890
rect 12479 16836 12535 16838
rect 12559 16836 12615 16838
rect 12639 16836 12695 16838
rect 12719 16836 12775 16838
rect 12714 16632 12770 16688
rect 12622 16360 12678 16416
rect 12254 15408 12310 15464
rect 12070 14864 12126 14920
rect 11978 14456 12034 14512
rect 12479 15802 12535 15804
rect 12559 15802 12615 15804
rect 12639 15802 12695 15804
rect 12719 15802 12775 15804
rect 12479 15750 12525 15802
rect 12525 15750 12535 15802
rect 12559 15750 12589 15802
rect 12589 15750 12601 15802
rect 12601 15750 12615 15802
rect 12639 15750 12653 15802
rect 12653 15750 12665 15802
rect 12665 15750 12695 15802
rect 12719 15750 12729 15802
rect 12729 15750 12775 15802
rect 12479 15748 12535 15750
rect 12559 15748 12615 15750
rect 12639 15748 12695 15750
rect 12719 15748 12775 15750
rect 12479 14714 12535 14716
rect 12559 14714 12615 14716
rect 12639 14714 12695 14716
rect 12719 14714 12775 14716
rect 12479 14662 12525 14714
rect 12525 14662 12535 14714
rect 12559 14662 12589 14714
rect 12589 14662 12601 14714
rect 12601 14662 12615 14714
rect 12639 14662 12653 14714
rect 12653 14662 12665 14714
rect 12665 14662 12695 14714
rect 12719 14662 12729 14714
rect 12729 14662 12775 14714
rect 12479 14660 12535 14662
rect 12559 14660 12615 14662
rect 12639 14660 12695 14662
rect 12719 14660 12775 14662
rect 12479 13626 12535 13628
rect 12559 13626 12615 13628
rect 12639 13626 12695 13628
rect 12719 13626 12775 13628
rect 12479 13574 12525 13626
rect 12525 13574 12535 13626
rect 12559 13574 12589 13626
rect 12589 13574 12601 13626
rect 12601 13574 12615 13626
rect 12639 13574 12653 13626
rect 12653 13574 12665 13626
rect 12665 13574 12695 13626
rect 12719 13574 12729 13626
rect 12729 13574 12775 13626
rect 12479 13572 12535 13574
rect 12559 13572 12615 13574
rect 12639 13572 12695 13574
rect 12719 13572 12775 13574
rect 12990 16496 13046 16552
rect 12898 12824 12954 12880
rect 12479 12538 12535 12540
rect 12559 12538 12615 12540
rect 12639 12538 12695 12540
rect 12719 12538 12775 12540
rect 12479 12486 12525 12538
rect 12525 12486 12535 12538
rect 12559 12486 12589 12538
rect 12589 12486 12601 12538
rect 12601 12486 12615 12538
rect 12639 12486 12653 12538
rect 12653 12486 12665 12538
rect 12665 12486 12695 12538
rect 12719 12486 12729 12538
rect 12729 12486 12775 12538
rect 12479 12484 12535 12486
rect 12559 12484 12615 12486
rect 12639 12484 12695 12486
rect 12719 12484 12775 12486
rect 11150 7928 11206 7984
rect 8638 7642 8694 7644
rect 8718 7642 8774 7644
rect 8798 7642 8854 7644
rect 8878 7642 8934 7644
rect 8638 7590 8684 7642
rect 8684 7590 8694 7642
rect 8718 7590 8748 7642
rect 8748 7590 8760 7642
rect 8760 7590 8774 7642
rect 8798 7590 8812 7642
rect 8812 7590 8824 7642
rect 8824 7590 8854 7642
rect 8878 7590 8888 7642
rect 8888 7590 8934 7642
rect 8638 7588 8694 7590
rect 8718 7588 8774 7590
rect 8798 7588 8854 7590
rect 8878 7588 8934 7590
rect 13450 18672 13506 18728
rect 13450 17604 13506 17640
rect 13450 17584 13452 17604
rect 13452 17584 13504 17604
rect 13504 17584 13506 17604
rect 13358 15852 13360 15872
rect 13360 15852 13412 15872
rect 13412 15852 13414 15872
rect 13358 15816 13414 15852
rect 13174 11600 13230 11656
rect 12990 11464 13046 11520
rect 12479 11450 12535 11452
rect 12559 11450 12615 11452
rect 12639 11450 12695 11452
rect 12719 11450 12775 11452
rect 12479 11398 12525 11450
rect 12525 11398 12535 11450
rect 12559 11398 12589 11450
rect 12589 11398 12601 11450
rect 12601 11398 12615 11450
rect 12639 11398 12653 11450
rect 12653 11398 12665 11450
rect 12665 11398 12695 11450
rect 12719 11398 12729 11450
rect 12729 11398 12775 11450
rect 12479 11396 12535 11398
rect 12559 11396 12615 11398
rect 12639 11396 12695 11398
rect 12719 11396 12775 11398
rect 12479 10362 12535 10364
rect 12559 10362 12615 10364
rect 12639 10362 12695 10364
rect 12719 10362 12775 10364
rect 12479 10310 12525 10362
rect 12525 10310 12535 10362
rect 12559 10310 12589 10362
rect 12589 10310 12601 10362
rect 12601 10310 12615 10362
rect 12639 10310 12653 10362
rect 12653 10310 12665 10362
rect 12665 10310 12695 10362
rect 12719 10310 12729 10362
rect 12729 10310 12775 10362
rect 12479 10308 12535 10310
rect 12559 10308 12615 10310
rect 12639 10308 12695 10310
rect 12719 10308 12775 10310
rect 13450 13640 13506 13696
rect 13726 19080 13782 19136
rect 15382 24692 15384 24712
rect 15384 24692 15436 24712
rect 15436 24692 15438 24712
rect 15382 24656 15438 24692
rect 15382 24520 15438 24576
rect 15290 23840 15346 23896
rect 15842 30096 15898 30152
rect 15750 29144 15806 29200
rect 15750 27512 15806 27568
rect 15658 27240 15714 27296
rect 15566 25880 15622 25936
rect 16118 31184 16174 31240
rect 16320 31578 16376 31580
rect 16400 31578 16456 31580
rect 16480 31578 16536 31580
rect 16560 31578 16616 31580
rect 16320 31526 16366 31578
rect 16366 31526 16376 31578
rect 16400 31526 16430 31578
rect 16430 31526 16442 31578
rect 16442 31526 16456 31578
rect 16480 31526 16494 31578
rect 16494 31526 16506 31578
rect 16506 31526 16536 31578
rect 16560 31526 16570 31578
rect 16570 31526 16616 31578
rect 16320 31524 16376 31526
rect 16400 31524 16456 31526
rect 16480 31524 16536 31526
rect 16560 31524 16616 31526
rect 16210 30912 16266 30968
rect 16118 30504 16174 30560
rect 16320 30490 16376 30492
rect 16400 30490 16456 30492
rect 16480 30490 16536 30492
rect 16560 30490 16616 30492
rect 16320 30438 16366 30490
rect 16366 30438 16376 30490
rect 16400 30438 16430 30490
rect 16430 30438 16442 30490
rect 16442 30438 16456 30490
rect 16480 30438 16494 30490
rect 16494 30438 16506 30490
rect 16506 30438 16536 30490
rect 16560 30438 16570 30490
rect 16570 30438 16616 30490
rect 16320 30436 16376 30438
rect 16400 30436 16456 30438
rect 16480 30436 16536 30438
rect 16560 30436 16616 30438
rect 15934 28212 15990 28248
rect 15934 28192 15936 28212
rect 15936 28192 15988 28212
rect 15988 28192 15990 28212
rect 15934 27512 15990 27568
rect 16320 29402 16376 29404
rect 16400 29402 16456 29404
rect 16480 29402 16536 29404
rect 16560 29402 16616 29404
rect 16320 29350 16366 29402
rect 16366 29350 16376 29402
rect 16400 29350 16430 29402
rect 16430 29350 16442 29402
rect 16442 29350 16456 29402
rect 16480 29350 16494 29402
rect 16494 29350 16506 29402
rect 16506 29350 16536 29402
rect 16560 29350 16570 29402
rect 16570 29350 16616 29402
rect 16320 29348 16376 29350
rect 16400 29348 16456 29350
rect 16480 29348 16536 29350
rect 16560 29348 16616 29350
rect 16210 29028 16266 29064
rect 16210 29008 16212 29028
rect 16212 29008 16264 29028
rect 16264 29008 16266 29028
rect 16854 30504 16910 30560
rect 17222 30776 17278 30832
rect 17130 30660 17186 30696
rect 17130 30640 17132 30660
rect 17132 30640 17184 30660
rect 17184 30640 17186 30660
rect 16762 29280 16818 29336
rect 16320 28314 16376 28316
rect 16400 28314 16456 28316
rect 16480 28314 16536 28316
rect 16560 28314 16616 28316
rect 16320 28262 16366 28314
rect 16366 28262 16376 28314
rect 16400 28262 16430 28314
rect 16430 28262 16442 28314
rect 16442 28262 16456 28314
rect 16480 28262 16494 28314
rect 16494 28262 16506 28314
rect 16506 28262 16536 28314
rect 16560 28262 16570 28314
rect 16570 28262 16616 28314
rect 16320 28260 16376 28262
rect 16400 28260 16456 28262
rect 16480 28260 16536 28262
rect 16560 28260 16616 28262
rect 16210 27512 16266 27568
rect 16026 26560 16082 26616
rect 15750 26016 15806 26072
rect 15566 24384 15622 24440
rect 15750 24248 15806 24304
rect 15014 20848 15070 20904
rect 15290 21936 15346 21992
rect 15750 23704 15806 23760
rect 15934 26152 15990 26208
rect 15934 25472 15990 25528
rect 15934 25200 15990 25256
rect 15934 25064 15990 25120
rect 15934 24676 15990 24712
rect 15934 24656 15936 24676
rect 15936 24656 15988 24676
rect 15988 24656 15990 24676
rect 16320 27226 16376 27228
rect 16400 27226 16456 27228
rect 16480 27226 16536 27228
rect 16560 27226 16616 27228
rect 16320 27174 16366 27226
rect 16366 27174 16376 27226
rect 16400 27174 16430 27226
rect 16430 27174 16442 27226
rect 16442 27174 16456 27226
rect 16480 27174 16494 27226
rect 16494 27174 16506 27226
rect 16506 27174 16536 27226
rect 16560 27174 16570 27226
rect 16570 27174 16616 27226
rect 16320 27172 16376 27174
rect 16400 27172 16456 27174
rect 16480 27172 16536 27174
rect 16560 27172 16616 27174
rect 16394 26324 16396 26344
rect 16396 26324 16448 26344
rect 16448 26324 16450 26344
rect 16394 26288 16450 26324
rect 16578 26832 16634 26888
rect 16854 28328 16910 28384
rect 17222 29452 17224 29472
rect 17224 29452 17276 29472
rect 17276 29452 17278 29472
rect 17222 29416 17278 29452
rect 16320 26138 16376 26140
rect 16400 26138 16456 26140
rect 16480 26138 16536 26140
rect 16560 26138 16616 26140
rect 16320 26086 16366 26138
rect 16366 26086 16376 26138
rect 16400 26086 16430 26138
rect 16430 26086 16442 26138
rect 16442 26086 16456 26138
rect 16480 26086 16494 26138
rect 16494 26086 16506 26138
rect 16506 26086 16536 26138
rect 16560 26086 16570 26138
rect 16570 26086 16616 26138
rect 16320 26084 16376 26086
rect 16400 26084 16456 26086
rect 16480 26084 16536 26086
rect 16560 26084 16616 26086
rect 16320 25050 16376 25052
rect 16400 25050 16456 25052
rect 16480 25050 16536 25052
rect 16560 25050 16616 25052
rect 16320 24998 16366 25050
rect 16366 24998 16376 25050
rect 16400 24998 16430 25050
rect 16430 24998 16442 25050
rect 16442 24998 16456 25050
rect 16480 24998 16494 25050
rect 16494 24998 16506 25050
rect 16506 24998 16536 25050
rect 16560 24998 16570 25050
rect 16570 24998 16616 25050
rect 16320 24996 16376 24998
rect 16400 24996 16456 24998
rect 16480 24996 16536 24998
rect 16560 24996 16616 24998
rect 15290 21548 15346 21584
rect 15290 21528 15292 21548
rect 15292 21528 15344 21548
rect 15344 21528 15346 21548
rect 15474 21800 15530 21856
rect 15290 20848 15346 20904
rect 16394 24656 16450 24712
rect 16578 24248 16634 24304
rect 16762 25492 16818 25528
rect 16762 25472 16764 25492
rect 16764 25472 16816 25492
rect 16816 25472 16818 25492
rect 16762 24928 16818 24984
rect 18050 32408 18106 32464
rect 19522 33088 19578 33144
rect 19246 32816 19302 32872
rect 17774 31456 17830 31512
rect 17498 27512 17554 27568
rect 17406 26832 17462 26888
rect 16854 24656 16910 24712
rect 16854 24248 16910 24304
rect 16118 23976 16174 24032
rect 16320 23962 16376 23964
rect 16400 23962 16456 23964
rect 16480 23962 16536 23964
rect 16560 23962 16616 23964
rect 16320 23910 16366 23962
rect 16366 23910 16376 23962
rect 16400 23910 16430 23962
rect 16430 23910 16442 23962
rect 16442 23910 16456 23962
rect 16480 23910 16494 23962
rect 16494 23910 16506 23962
rect 16506 23910 16536 23962
rect 16560 23910 16570 23962
rect 16570 23910 16616 23962
rect 16320 23908 16376 23910
rect 16400 23908 16456 23910
rect 16480 23908 16536 23910
rect 16560 23908 16616 23910
rect 16762 23976 16818 24032
rect 16210 23296 16266 23352
rect 15842 22752 15898 22808
rect 15842 22344 15898 22400
rect 16394 23296 16450 23352
rect 16026 22888 16082 22944
rect 16320 22874 16376 22876
rect 16400 22874 16456 22876
rect 16480 22874 16536 22876
rect 16560 22874 16616 22876
rect 16320 22822 16366 22874
rect 16366 22822 16376 22874
rect 16400 22822 16430 22874
rect 16430 22822 16442 22874
rect 16442 22822 16456 22874
rect 16480 22822 16494 22874
rect 16494 22822 16506 22874
rect 16506 22822 16536 22874
rect 16560 22822 16570 22874
rect 16570 22822 16616 22874
rect 16320 22820 16376 22822
rect 16400 22820 16456 22822
rect 16480 22820 16536 22822
rect 16560 22820 16616 22822
rect 16670 22208 16726 22264
rect 16118 21800 16174 21856
rect 16118 21684 16174 21720
rect 16118 21664 16120 21684
rect 16120 21664 16172 21684
rect 16172 21664 16174 21684
rect 16320 21786 16376 21788
rect 16400 21786 16456 21788
rect 16480 21786 16536 21788
rect 16560 21786 16616 21788
rect 16320 21734 16366 21786
rect 16366 21734 16376 21786
rect 16400 21734 16430 21786
rect 16430 21734 16442 21786
rect 16442 21734 16456 21786
rect 16480 21734 16494 21786
rect 16494 21734 16506 21786
rect 16506 21734 16536 21786
rect 16560 21734 16570 21786
rect 16570 21734 16616 21786
rect 16320 21732 16376 21734
rect 16400 21732 16456 21734
rect 16480 21732 16536 21734
rect 16560 21732 16616 21734
rect 16026 21120 16082 21176
rect 16394 21120 16450 21176
rect 17222 26152 17278 26208
rect 17498 26424 17554 26480
rect 17314 26016 17370 26072
rect 17130 25492 17186 25528
rect 17130 25472 17132 25492
rect 17132 25472 17184 25492
rect 17184 25472 17186 25492
rect 17774 29416 17830 29472
rect 17590 26288 17646 26344
rect 17682 25644 17684 25664
rect 17684 25644 17736 25664
rect 17736 25644 17738 25664
rect 17682 25608 17738 25644
rect 17498 25492 17554 25528
rect 17498 25472 17500 25492
rect 17500 25472 17552 25492
rect 17552 25472 17554 25492
rect 18142 30232 18198 30288
rect 17866 27512 17922 27568
rect 18050 27512 18106 27568
rect 18234 28872 18290 28928
rect 18970 30640 19026 30696
rect 18786 29724 18788 29744
rect 18788 29724 18840 29744
rect 18840 29724 18842 29744
rect 18786 29688 18842 29724
rect 18510 29552 18566 29608
rect 18694 29552 18750 29608
rect 18602 29280 18658 29336
rect 18510 28872 18566 28928
rect 18786 28600 18842 28656
rect 18602 28212 18658 28248
rect 18602 28192 18604 28212
rect 18604 28192 18656 28212
rect 18656 28192 18658 28212
rect 18418 27784 18474 27840
rect 18326 27104 18382 27160
rect 17866 26580 17922 26616
rect 17866 26560 17868 26580
rect 17868 26560 17920 26580
rect 17920 26560 17922 26580
rect 17958 26424 18014 26480
rect 17130 24792 17186 24848
rect 17314 24792 17370 24848
rect 17130 23296 17186 23352
rect 16946 22208 17002 22264
rect 17590 25200 17646 25256
rect 17498 24656 17554 24712
rect 17406 24384 17462 24440
rect 17498 24248 17554 24304
rect 17314 23840 17370 23896
rect 17590 23840 17646 23896
rect 18326 26696 18382 26752
rect 18142 26424 18198 26480
rect 18326 26288 18382 26344
rect 17774 25064 17830 25120
rect 17958 25064 18014 25120
rect 18326 26152 18382 26208
rect 18234 26016 18290 26072
rect 18418 26016 18474 26072
rect 18418 25900 18474 25936
rect 18418 25880 18420 25900
rect 18420 25880 18472 25900
rect 18472 25880 18474 25900
rect 18602 27784 18658 27840
rect 18970 28192 19026 28248
rect 18970 27920 19026 27976
rect 19246 30776 19302 30832
rect 20161 32122 20217 32124
rect 20241 32122 20297 32124
rect 20321 32122 20377 32124
rect 20401 32122 20457 32124
rect 20161 32070 20207 32122
rect 20207 32070 20217 32122
rect 20241 32070 20271 32122
rect 20271 32070 20283 32122
rect 20283 32070 20297 32122
rect 20321 32070 20335 32122
rect 20335 32070 20347 32122
rect 20347 32070 20377 32122
rect 20401 32070 20411 32122
rect 20411 32070 20457 32122
rect 20161 32068 20217 32070
rect 20241 32068 20297 32070
rect 20321 32068 20377 32070
rect 20401 32068 20457 32070
rect 19614 31592 19670 31648
rect 19338 30368 19394 30424
rect 19522 30232 19578 30288
rect 19430 29960 19486 30016
rect 19338 29552 19394 29608
rect 19246 29164 19302 29200
rect 19246 29144 19248 29164
rect 19248 29144 19300 29164
rect 19300 29144 19302 29164
rect 19246 28872 19302 28928
rect 19154 27920 19210 27976
rect 18878 27648 18934 27704
rect 18602 26288 18658 26344
rect 18602 26016 18658 26072
rect 17958 24656 18014 24712
rect 18142 24248 18198 24304
rect 17958 23976 18014 24032
rect 17774 23160 17830 23216
rect 18142 23976 18198 24032
rect 18142 23840 18198 23896
rect 17406 22888 17462 22944
rect 17314 22752 17370 22808
rect 17222 22616 17278 22672
rect 17222 22072 17278 22128
rect 17130 21936 17186 21992
rect 17314 21528 17370 21584
rect 16670 20984 16726 21040
rect 16302 20848 16358 20904
rect 15658 20748 15660 20768
rect 15660 20748 15712 20768
rect 15712 20748 15714 20768
rect 15658 20712 15714 20748
rect 15198 20168 15254 20224
rect 14830 20032 14886 20088
rect 14462 18944 14518 19000
rect 13910 18808 13966 18864
rect 13818 18264 13874 18320
rect 14462 18672 14518 18728
rect 14094 18300 14096 18320
rect 14096 18300 14148 18320
rect 14148 18300 14150 18320
rect 14094 18264 14150 18300
rect 13910 15036 13912 15056
rect 13912 15036 13964 15056
rect 13964 15036 13966 15056
rect 13910 15000 13966 15036
rect 14094 16768 14150 16824
rect 14186 16632 14242 16688
rect 14186 15972 14242 16008
rect 14186 15952 14188 15972
rect 14188 15952 14240 15972
rect 14240 15952 14242 15972
rect 14922 19116 14924 19136
rect 14924 19116 14976 19136
rect 14976 19116 14978 19136
rect 14922 19080 14978 19116
rect 14922 18400 14978 18456
rect 15382 20032 15438 20088
rect 14830 18028 14832 18048
rect 14832 18028 14884 18048
rect 14884 18028 14886 18048
rect 14830 17992 14886 18028
rect 14554 17876 14610 17912
rect 14554 17856 14556 17876
rect 14556 17856 14608 17876
rect 14608 17856 14610 17876
rect 15382 18808 15438 18864
rect 14922 17720 14978 17776
rect 15106 17756 15108 17776
rect 15108 17756 15160 17776
rect 15160 17756 15162 17776
rect 15106 17720 15162 17756
rect 14554 17040 14610 17096
rect 14462 16768 14518 16824
rect 14370 16632 14426 16688
rect 14462 16396 14464 16416
rect 14464 16396 14516 16416
rect 14516 16396 14518 16416
rect 14462 16360 14518 16396
rect 16320 20698 16376 20700
rect 16400 20698 16456 20700
rect 16480 20698 16536 20700
rect 16560 20698 16616 20700
rect 16320 20646 16366 20698
rect 16366 20646 16376 20698
rect 16400 20646 16430 20698
rect 16430 20646 16442 20698
rect 16442 20646 16456 20698
rect 16480 20646 16494 20698
rect 16494 20646 16506 20698
rect 16506 20646 16536 20698
rect 16560 20646 16570 20698
rect 16570 20646 16616 20698
rect 16320 20644 16376 20646
rect 16400 20644 16456 20646
rect 16480 20644 16536 20646
rect 16560 20644 16616 20646
rect 16118 20576 16174 20632
rect 16762 20576 16818 20632
rect 17774 22888 17830 22944
rect 17866 22752 17922 22808
rect 17682 22208 17738 22264
rect 17682 21936 17738 21992
rect 17774 21528 17830 21584
rect 18418 24248 18474 24304
rect 18326 23840 18382 23896
rect 18326 23296 18382 23352
rect 17958 21956 18014 21992
rect 18418 22888 18474 22944
rect 18418 22752 18474 22808
rect 18602 24520 18658 24576
rect 19062 27512 19118 27568
rect 18878 25608 18934 25664
rect 18786 24928 18842 24984
rect 19062 26016 19118 26072
rect 19430 28872 19486 28928
rect 19338 28600 19394 28656
rect 19430 28328 19486 28384
rect 19430 26560 19486 26616
rect 20534 32000 20590 32056
rect 19982 31048 20038 31104
rect 20161 31034 20217 31036
rect 20241 31034 20297 31036
rect 20321 31034 20377 31036
rect 20401 31034 20457 31036
rect 20161 30982 20207 31034
rect 20207 30982 20217 31034
rect 20241 30982 20271 31034
rect 20271 30982 20283 31034
rect 20283 30982 20297 31034
rect 20321 30982 20335 31034
rect 20335 30982 20347 31034
rect 20347 30982 20377 31034
rect 20401 30982 20411 31034
rect 20411 30982 20457 31034
rect 20161 30980 20217 30982
rect 20241 30980 20297 30982
rect 20321 30980 20377 30982
rect 20401 30980 20457 30982
rect 20534 30912 20590 30968
rect 20074 30640 20130 30696
rect 19614 27784 19670 27840
rect 19890 30232 19946 30288
rect 19890 29824 19946 29880
rect 19890 29416 19946 29472
rect 20350 30776 20406 30832
rect 20350 30540 20352 30560
rect 20352 30540 20404 30560
rect 20404 30540 20406 30560
rect 20350 30504 20406 30540
rect 20258 30368 20314 30424
rect 20442 30368 20498 30424
rect 20718 31048 20774 31104
rect 20718 30232 20774 30288
rect 20161 29946 20217 29948
rect 20241 29946 20297 29948
rect 20321 29946 20377 29948
rect 20401 29946 20457 29948
rect 20161 29894 20207 29946
rect 20207 29894 20217 29946
rect 20241 29894 20271 29946
rect 20271 29894 20283 29946
rect 20283 29894 20297 29946
rect 20321 29894 20335 29946
rect 20335 29894 20347 29946
rect 20347 29894 20377 29946
rect 20401 29894 20411 29946
rect 20411 29894 20457 29946
rect 20161 29892 20217 29894
rect 20241 29892 20297 29894
rect 20321 29892 20377 29894
rect 20401 29892 20457 29894
rect 19798 27648 19854 27704
rect 20161 28858 20217 28860
rect 20241 28858 20297 28860
rect 20321 28858 20377 28860
rect 20401 28858 20457 28860
rect 20161 28806 20207 28858
rect 20207 28806 20217 28858
rect 20241 28806 20271 28858
rect 20271 28806 20283 28858
rect 20283 28806 20297 28858
rect 20321 28806 20335 28858
rect 20335 28806 20347 28858
rect 20347 28806 20377 28858
rect 20401 28806 20411 28858
rect 20411 28806 20457 28858
rect 20161 28804 20217 28806
rect 20241 28804 20297 28806
rect 20321 28804 20377 28806
rect 20401 28804 20457 28806
rect 19982 28736 20038 28792
rect 20626 29960 20682 30016
rect 20994 30504 21050 30560
rect 20902 30232 20958 30288
rect 20810 29688 20866 29744
rect 20626 29552 20682 29608
rect 20810 29280 20866 29336
rect 20626 28872 20682 28928
rect 20350 28600 20406 28656
rect 20718 28736 20774 28792
rect 20994 29416 21050 29472
rect 20718 28464 20774 28520
rect 20902 28464 20958 28520
rect 21362 32408 21418 32464
rect 21546 30368 21602 30424
rect 21454 29688 21510 29744
rect 21454 29416 21510 29472
rect 19798 26832 19854 26888
rect 19614 26560 19670 26616
rect 20161 27770 20217 27772
rect 20241 27770 20297 27772
rect 20321 27770 20377 27772
rect 20401 27770 20457 27772
rect 20161 27718 20207 27770
rect 20207 27718 20217 27770
rect 20241 27718 20271 27770
rect 20271 27718 20283 27770
rect 20283 27718 20297 27770
rect 20321 27718 20335 27770
rect 20335 27718 20347 27770
rect 20347 27718 20377 27770
rect 20401 27718 20411 27770
rect 20411 27718 20457 27770
rect 20161 27716 20217 27718
rect 20241 27716 20297 27718
rect 20321 27716 20377 27718
rect 20401 27716 20457 27718
rect 20258 27512 20314 27568
rect 20994 27920 21050 27976
rect 20810 27784 20866 27840
rect 20534 26696 20590 26752
rect 20161 26682 20217 26684
rect 20241 26682 20297 26684
rect 20321 26682 20377 26684
rect 20401 26682 20457 26684
rect 20161 26630 20207 26682
rect 20207 26630 20217 26682
rect 20241 26630 20271 26682
rect 20271 26630 20283 26682
rect 20283 26630 20297 26682
rect 20321 26630 20335 26682
rect 20335 26630 20347 26682
rect 20347 26630 20377 26682
rect 20401 26630 20411 26682
rect 20411 26630 20457 26682
rect 20161 26628 20217 26630
rect 20241 26628 20297 26630
rect 20321 26628 20377 26630
rect 20401 26628 20457 26630
rect 19338 25356 19394 25392
rect 19338 25336 19340 25356
rect 19340 25336 19392 25356
rect 19392 25336 19394 25356
rect 19522 25336 19578 25392
rect 19062 24928 19118 24984
rect 18878 24520 18934 24576
rect 18878 24248 18934 24304
rect 18602 22344 18658 22400
rect 18786 22208 18842 22264
rect 18418 22108 18420 22128
rect 18420 22108 18472 22128
rect 18472 22108 18474 22128
rect 18418 22072 18474 22108
rect 19062 23976 19118 24032
rect 19798 25744 19854 25800
rect 19430 24928 19486 24984
rect 19430 24520 19486 24576
rect 20074 25744 20130 25800
rect 20258 26288 20314 26344
rect 20718 26560 20774 26616
rect 20161 25594 20217 25596
rect 20241 25594 20297 25596
rect 20321 25594 20377 25596
rect 20401 25594 20457 25596
rect 20161 25542 20207 25594
rect 20207 25542 20217 25594
rect 20241 25542 20271 25594
rect 20271 25542 20283 25594
rect 20283 25542 20297 25594
rect 20321 25542 20335 25594
rect 20335 25542 20347 25594
rect 20347 25542 20377 25594
rect 20401 25542 20411 25594
rect 20411 25542 20457 25594
rect 20161 25540 20217 25542
rect 20241 25540 20297 25542
rect 20321 25540 20377 25542
rect 20401 25540 20457 25542
rect 20074 25200 20130 25256
rect 19614 24520 19670 24576
rect 19522 24384 19578 24440
rect 19246 23704 19302 23760
rect 19062 23296 19118 23352
rect 19430 23432 19486 23488
rect 17958 21936 17960 21956
rect 17960 21936 18012 21956
rect 18012 21936 18014 21956
rect 18050 21800 18106 21856
rect 18234 21684 18290 21720
rect 18234 21664 18236 21684
rect 18236 21664 18288 21684
rect 18288 21664 18290 21684
rect 18510 21664 18566 21720
rect 17866 21392 17922 21448
rect 18694 21664 18750 21720
rect 18878 21664 18934 21720
rect 19338 22752 19394 22808
rect 19062 21664 19118 21720
rect 17314 20848 17370 20904
rect 17682 20868 17738 20904
rect 17682 20848 17684 20868
rect 17684 20848 17736 20868
rect 17736 20848 17738 20868
rect 18142 20712 18198 20768
rect 15842 19624 15898 19680
rect 15750 18808 15806 18864
rect 16118 19488 16174 19544
rect 17406 19896 17462 19952
rect 16762 19624 16818 19680
rect 16320 19610 16376 19612
rect 16400 19610 16456 19612
rect 16480 19610 16536 19612
rect 16560 19610 16616 19612
rect 16320 19558 16366 19610
rect 16366 19558 16376 19610
rect 16400 19558 16430 19610
rect 16430 19558 16442 19610
rect 16442 19558 16456 19610
rect 16480 19558 16494 19610
rect 16494 19558 16506 19610
rect 16506 19558 16536 19610
rect 16560 19558 16570 19610
rect 16570 19558 16616 19610
rect 16320 19556 16376 19558
rect 16400 19556 16456 19558
rect 16480 19556 16536 19558
rect 16560 19556 16616 19558
rect 16302 19372 16358 19408
rect 16302 19352 16304 19372
rect 16304 19352 16356 19372
rect 16356 19352 16358 19372
rect 16854 19488 16910 19544
rect 16578 18944 16634 19000
rect 16762 18944 16818 19000
rect 16026 18420 16082 18456
rect 16026 18400 16028 18420
rect 16028 18400 16080 18420
rect 16080 18400 16082 18420
rect 14738 16360 14794 16416
rect 14554 13912 14610 13968
rect 14738 13812 14740 13832
rect 14740 13812 14792 13832
rect 14792 13812 14794 13832
rect 14738 13776 14794 13812
rect 15198 16224 15254 16280
rect 16320 18522 16376 18524
rect 16400 18522 16456 18524
rect 16480 18522 16536 18524
rect 16560 18522 16616 18524
rect 16320 18470 16366 18522
rect 16366 18470 16376 18522
rect 16400 18470 16430 18522
rect 16430 18470 16442 18522
rect 16442 18470 16456 18522
rect 16480 18470 16494 18522
rect 16494 18470 16506 18522
rect 16506 18470 16536 18522
rect 16560 18470 16570 18522
rect 16570 18470 16616 18522
rect 16320 18468 16376 18470
rect 16400 18468 16456 18470
rect 16480 18468 16536 18470
rect 16560 18468 16616 18470
rect 16946 19080 17002 19136
rect 16762 18400 16818 18456
rect 15750 17856 15806 17912
rect 15842 17312 15898 17368
rect 15750 17040 15806 17096
rect 16394 17856 16450 17912
rect 17222 18808 17278 18864
rect 17038 18400 17094 18456
rect 16486 17720 16542 17776
rect 16026 17312 16082 17368
rect 15934 16904 15990 16960
rect 15382 16224 15438 16280
rect 15290 15680 15346 15736
rect 15198 15544 15254 15600
rect 12479 9274 12535 9276
rect 12559 9274 12615 9276
rect 12639 9274 12695 9276
rect 12719 9274 12775 9276
rect 12479 9222 12525 9274
rect 12525 9222 12535 9274
rect 12559 9222 12589 9274
rect 12589 9222 12601 9274
rect 12601 9222 12615 9274
rect 12639 9222 12653 9274
rect 12653 9222 12665 9274
rect 12665 9222 12695 9274
rect 12719 9222 12729 9274
rect 12729 9222 12775 9274
rect 12479 9220 12535 9222
rect 12559 9220 12615 9222
rect 12639 9220 12695 9222
rect 12719 9220 12775 9222
rect 15842 16360 15898 16416
rect 15014 14320 15070 14376
rect 15474 14612 15530 14648
rect 15474 14592 15476 14612
rect 15476 14592 15528 14612
rect 15528 14592 15530 14612
rect 15658 12552 15714 12608
rect 16026 16396 16028 16416
rect 16028 16396 16080 16416
rect 16080 16396 16082 16416
rect 16026 16360 16082 16396
rect 16320 17434 16376 17436
rect 16400 17434 16456 17436
rect 16480 17434 16536 17436
rect 16560 17434 16616 17436
rect 16320 17382 16366 17434
rect 16366 17382 16376 17434
rect 16400 17382 16430 17434
rect 16430 17382 16442 17434
rect 16442 17382 16456 17434
rect 16480 17382 16494 17434
rect 16494 17382 16506 17434
rect 16506 17382 16536 17434
rect 16560 17382 16570 17434
rect 16570 17382 16616 17434
rect 16320 17380 16376 17382
rect 16400 17380 16456 17382
rect 16480 17380 16536 17382
rect 16560 17380 16616 17382
rect 16578 17076 16580 17096
rect 16580 17076 16632 17096
rect 16632 17076 16634 17096
rect 16578 17040 16634 17076
rect 16320 16346 16376 16348
rect 16400 16346 16456 16348
rect 16480 16346 16536 16348
rect 16560 16346 16616 16348
rect 16320 16294 16366 16346
rect 16366 16294 16376 16346
rect 16400 16294 16430 16346
rect 16430 16294 16442 16346
rect 16442 16294 16456 16346
rect 16480 16294 16494 16346
rect 16494 16294 16506 16346
rect 16506 16294 16536 16346
rect 16560 16294 16570 16346
rect 16570 16294 16616 16346
rect 16320 16292 16376 16294
rect 16400 16292 16456 16294
rect 16480 16292 16536 16294
rect 16560 16292 16616 16294
rect 16762 16360 16818 16416
rect 16946 17448 17002 17504
rect 16946 17332 17002 17368
rect 16946 17312 16948 17332
rect 16948 17312 17000 17332
rect 17000 17312 17002 17332
rect 17222 18536 17278 18592
rect 18142 20168 18198 20224
rect 18050 20032 18106 20088
rect 18234 20052 18290 20088
rect 18234 20032 18236 20052
rect 18236 20032 18288 20052
rect 18288 20032 18290 20052
rect 18234 19896 18290 19952
rect 17590 19080 17646 19136
rect 17682 18944 17738 19000
rect 18050 19080 18106 19136
rect 18418 20168 18474 20224
rect 18418 20032 18474 20088
rect 18878 20576 18934 20632
rect 18234 19080 18290 19136
rect 18142 18944 18198 19000
rect 17130 17448 17186 17504
rect 16946 16360 17002 16416
rect 16394 15680 16450 15736
rect 16320 15258 16376 15260
rect 16400 15258 16456 15260
rect 16480 15258 16536 15260
rect 16560 15258 16616 15260
rect 16320 15206 16366 15258
rect 16366 15206 16376 15258
rect 16400 15206 16430 15258
rect 16430 15206 16442 15258
rect 16442 15206 16456 15258
rect 16480 15206 16494 15258
rect 16494 15206 16506 15258
rect 16506 15206 16536 15258
rect 16560 15206 16570 15258
rect 16570 15206 16616 15258
rect 16320 15204 16376 15206
rect 16400 15204 16456 15206
rect 16480 15204 16536 15206
rect 16560 15204 16616 15206
rect 16762 15136 16818 15192
rect 16762 14456 16818 14512
rect 15934 14184 15990 14240
rect 15842 14048 15898 14104
rect 16026 12416 16082 12472
rect 16320 14170 16376 14172
rect 16400 14170 16456 14172
rect 16480 14170 16536 14172
rect 16560 14170 16616 14172
rect 16320 14118 16366 14170
rect 16366 14118 16376 14170
rect 16400 14118 16430 14170
rect 16430 14118 16442 14170
rect 16442 14118 16456 14170
rect 16480 14118 16494 14170
rect 16494 14118 16506 14170
rect 16506 14118 16536 14170
rect 16560 14118 16570 14170
rect 16570 14118 16616 14170
rect 16320 14116 16376 14118
rect 16400 14116 16456 14118
rect 16480 14116 16536 14118
rect 16560 14116 16616 14118
rect 16302 13232 16358 13288
rect 16320 13082 16376 13084
rect 16400 13082 16456 13084
rect 16480 13082 16536 13084
rect 16560 13082 16616 13084
rect 16320 13030 16366 13082
rect 16366 13030 16376 13082
rect 16400 13030 16430 13082
rect 16430 13030 16442 13082
rect 16442 13030 16456 13082
rect 16480 13030 16494 13082
rect 16494 13030 16506 13082
rect 16506 13030 16536 13082
rect 16560 13030 16570 13082
rect 16570 13030 16616 13082
rect 16320 13028 16376 13030
rect 16400 13028 16456 13030
rect 16480 13028 16536 13030
rect 16560 13028 16616 13030
rect 16762 13096 16818 13152
rect 17406 17856 17462 17912
rect 17590 17856 17646 17912
rect 17314 17312 17370 17368
rect 16946 14184 17002 14240
rect 17498 16904 17554 16960
rect 17866 16904 17922 16960
rect 17774 16768 17830 16824
rect 17498 15544 17554 15600
rect 17774 15544 17830 15600
rect 17498 14456 17554 14512
rect 16946 14048 17002 14104
rect 17222 13776 17278 13832
rect 16854 12960 16910 13016
rect 16320 11994 16376 11996
rect 16400 11994 16456 11996
rect 16480 11994 16536 11996
rect 16560 11994 16616 11996
rect 16320 11942 16366 11994
rect 16366 11942 16376 11994
rect 16400 11942 16430 11994
rect 16430 11942 16442 11994
rect 16442 11942 16456 11994
rect 16480 11942 16494 11994
rect 16494 11942 16506 11994
rect 16506 11942 16536 11994
rect 16560 11942 16570 11994
rect 16570 11942 16616 11994
rect 16320 11940 16376 11942
rect 16400 11940 16456 11942
rect 16480 11940 16536 11942
rect 16560 11940 16616 11942
rect 17498 13912 17554 13968
rect 17774 15000 17830 15056
rect 17866 14476 17922 14512
rect 17866 14456 17868 14476
rect 17868 14456 17920 14476
rect 17920 14456 17922 14476
rect 18694 19780 18750 19816
rect 18694 19760 18696 19780
rect 18696 19760 18748 19780
rect 18748 19760 18750 19780
rect 18878 19760 18934 19816
rect 19246 19896 19302 19952
rect 19154 19760 19210 19816
rect 18786 19624 18842 19680
rect 18970 19624 19026 19680
rect 18786 19488 18842 19544
rect 18694 19352 18750 19408
rect 18326 17584 18382 17640
rect 18510 17584 18566 17640
rect 19154 19352 19210 19408
rect 19154 19080 19210 19136
rect 18050 15000 18106 15056
rect 18050 14728 18106 14784
rect 17958 13096 18014 13152
rect 16320 10906 16376 10908
rect 16400 10906 16456 10908
rect 16480 10906 16536 10908
rect 16560 10906 16616 10908
rect 16320 10854 16366 10906
rect 16366 10854 16376 10906
rect 16400 10854 16430 10906
rect 16430 10854 16442 10906
rect 16442 10854 16456 10906
rect 16480 10854 16494 10906
rect 16494 10854 16506 10906
rect 16506 10854 16536 10906
rect 16560 10854 16570 10906
rect 16570 10854 16616 10906
rect 16320 10852 16376 10854
rect 16400 10852 16456 10854
rect 16480 10852 16536 10854
rect 16560 10852 16616 10854
rect 17774 11892 17830 11928
rect 17774 11872 17776 11892
rect 17776 11872 17828 11892
rect 17828 11872 17830 11892
rect 18418 16904 18474 16960
rect 18418 16224 18474 16280
rect 18234 15816 18290 15872
rect 18234 15680 18290 15736
rect 18602 15816 18658 15872
rect 18878 15680 18934 15736
rect 19338 19080 19394 19136
rect 19062 16224 19118 16280
rect 19890 24520 19946 24576
rect 19798 24384 19854 24440
rect 19706 23840 19762 23896
rect 20350 24928 20406 24984
rect 19982 24384 20038 24440
rect 20161 24506 20217 24508
rect 20241 24506 20297 24508
rect 20321 24506 20377 24508
rect 20401 24506 20457 24508
rect 20161 24454 20207 24506
rect 20207 24454 20217 24506
rect 20241 24454 20271 24506
rect 20271 24454 20283 24506
rect 20283 24454 20297 24506
rect 20321 24454 20335 24506
rect 20335 24454 20347 24506
rect 20347 24454 20377 24506
rect 20401 24454 20411 24506
rect 20411 24454 20457 24506
rect 20161 24452 20217 24454
rect 20241 24452 20297 24454
rect 20321 24452 20377 24454
rect 20401 24452 20457 24454
rect 19706 23296 19762 23352
rect 19706 22480 19762 22536
rect 19798 22344 19854 22400
rect 20534 23432 20590 23488
rect 20161 23418 20217 23420
rect 20241 23418 20297 23420
rect 20321 23418 20377 23420
rect 20401 23418 20457 23420
rect 20161 23366 20207 23418
rect 20207 23366 20217 23418
rect 20241 23366 20271 23418
rect 20271 23366 20283 23418
rect 20283 23366 20297 23418
rect 20321 23366 20335 23418
rect 20335 23366 20347 23418
rect 20347 23366 20377 23418
rect 20401 23366 20411 23418
rect 20411 23366 20457 23418
rect 20161 23364 20217 23366
rect 20241 23364 20297 23366
rect 20321 23364 20377 23366
rect 20401 23364 20457 23366
rect 20161 22330 20217 22332
rect 20241 22330 20297 22332
rect 20321 22330 20377 22332
rect 20401 22330 20457 22332
rect 20161 22278 20207 22330
rect 20207 22278 20217 22330
rect 20241 22278 20271 22330
rect 20271 22278 20283 22330
rect 20283 22278 20297 22330
rect 20321 22278 20335 22330
rect 20335 22278 20347 22330
rect 20347 22278 20377 22330
rect 20401 22278 20411 22330
rect 20411 22278 20457 22330
rect 20161 22276 20217 22278
rect 20241 22276 20297 22278
rect 20321 22276 20377 22278
rect 20401 22276 20457 22278
rect 19982 22208 20038 22264
rect 19614 21664 19670 21720
rect 19982 21256 20038 21312
rect 20534 21256 20590 21312
rect 20161 21242 20217 21244
rect 20241 21242 20297 21244
rect 20321 21242 20377 21244
rect 20401 21242 20457 21244
rect 20161 21190 20207 21242
rect 20207 21190 20217 21242
rect 20241 21190 20271 21242
rect 20271 21190 20283 21242
rect 20283 21190 20297 21242
rect 20321 21190 20335 21242
rect 20335 21190 20347 21242
rect 20347 21190 20377 21242
rect 20401 21190 20411 21242
rect 20411 21190 20457 21242
rect 20161 21188 20217 21190
rect 20241 21188 20297 21190
rect 20321 21188 20377 21190
rect 20401 21188 20457 21190
rect 21546 29144 21602 29200
rect 21086 27512 21142 27568
rect 21086 27412 21088 27432
rect 21088 27412 21140 27432
rect 21140 27412 21142 27432
rect 21086 27376 21142 27412
rect 21362 27512 21418 27568
rect 21178 26968 21234 27024
rect 21546 27784 21602 27840
rect 21638 27668 21694 27704
rect 21638 27648 21640 27668
rect 21640 27648 21692 27668
rect 21692 27648 21694 27668
rect 21270 26424 21326 26480
rect 21178 26324 21180 26344
rect 21180 26324 21232 26344
rect 21232 26324 21234 26344
rect 21178 26288 21234 26324
rect 21178 26152 21234 26208
rect 21362 26188 21364 26208
rect 21364 26188 21416 26208
rect 21416 26188 21418 26208
rect 21362 26152 21418 26188
rect 21270 25880 21326 25936
rect 21362 25744 21418 25800
rect 23570 32680 23626 32736
rect 24002 32666 24058 32668
rect 24082 32666 24138 32668
rect 24162 32666 24218 32668
rect 24242 32666 24298 32668
rect 24002 32614 24048 32666
rect 24048 32614 24058 32666
rect 24082 32614 24112 32666
rect 24112 32614 24124 32666
rect 24124 32614 24138 32666
rect 24162 32614 24176 32666
rect 24176 32614 24188 32666
rect 24188 32614 24218 32666
rect 24242 32614 24252 32666
rect 24252 32614 24298 32666
rect 24002 32612 24058 32614
rect 24082 32612 24138 32614
rect 24162 32612 24218 32614
rect 24242 32612 24298 32614
rect 21822 28736 21878 28792
rect 22650 31864 22706 31920
rect 22190 30504 22246 30560
rect 22190 29688 22246 29744
rect 22374 29552 22430 29608
rect 22006 28756 22062 28792
rect 22006 28736 22008 28756
rect 22008 28736 22060 28756
rect 22060 28736 22062 28756
rect 21822 27784 21878 27840
rect 21822 27512 21878 27568
rect 21362 25200 21418 25256
rect 21086 24928 21142 24984
rect 20994 24384 21050 24440
rect 21086 24248 21142 24304
rect 20994 24112 21050 24168
rect 20902 22480 20958 22536
rect 20810 22344 20866 22400
rect 21086 23432 21142 23488
rect 21546 24928 21602 24984
rect 22190 28192 22246 28248
rect 22098 27920 22154 27976
rect 22006 27512 22062 27568
rect 22282 27240 22338 27296
rect 22650 31048 22706 31104
rect 23478 31592 23534 31648
rect 23294 31048 23350 31104
rect 23202 30268 23204 30288
rect 23204 30268 23256 30288
rect 23256 30268 23258 30288
rect 23202 30232 23258 30268
rect 22926 29552 22982 29608
rect 23202 29996 23204 30016
rect 23204 29996 23256 30016
rect 23256 29996 23258 30016
rect 23202 29960 23258 29996
rect 22742 29008 22798 29064
rect 22558 28872 22614 28928
rect 22558 28192 22614 28248
rect 22558 27784 22614 27840
rect 22466 27512 22522 27568
rect 22466 27240 22522 27296
rect 22374 26968 22430 27024
rect 22098 26560 22154 26616
rect 22282 26560 22338 26616
rect 21822 25880 21878 25936
rect 21730 25064 21786 25120
rect 21546 24384 21602 24440
rect 21454 23976 21510 24032
rect 21454 23704 21510 23760
rect 21362 23432 21418 23488
rect 21270 22616 21326 22672
rect 19614 20032 19670 20088
rect 19890 20204 19892 20224
rect 19892 20204 19944 20224
rect 19944 20204 19946 20224
rect 19890 20168 19946 20204
rect 19522 18944 19578 19000
rect 19798 19488 19854 19544
rect 19522 18672 19578 18728
rect 21086 21256 21142 21312
rect 20902 20848 20958 20904
rect 20161 20154 20217 20156
rect 20241 20154 20297 20156
rect 20321 20154 20377 20156
rect 20401 20154 20457 20156
rect 20161 20102 20207 20154
rect 20207 20102 20217 20154
rect 20241 20102 20271 20154
rect 20271 20102 20283 20154
rect 20283 20102 20297 20154
rect 20321 20102 20335 20154
rect 20335 20102 20347 20154
rect 20347 20102 20377 20154
rect 20401 20102 20411 20154
rect 20411 20102 20457 20154
rect 20161 20100 20217 20102
rect 20241 20100 20297 20102
rect 20321 20100 20377 20102
rect 20401 20100 20457 20102
rect 20626 20168 20682 20224
rect 20074 19624 20130 19680
rect 19890 19080 19946 19136
rect 20534 19080 20590 19136
rect 20161 19066 20217 19068
rect 20241 19066 20297 19068
rect 20321 19066 20377 19068
rect 20401 19066 20457 19068
rect 20161 19014 20207 19066
rect 20207 19014 20217 19066
rect 20241 19014 20271 19066
rect 20271 19014 20283 19066
rect 20283 19014 20297 19066
rect 20321 19014 20335 19066
rect 20335 19014 20347 19066
rect 20347 19014 20377 19066
rect 20401 19014 20411 19066
rect 20411 19014 20457 19066
rect 20161 19012 20217 19014
rect 20241 19012 20297 19014
rect 20321 19012 20377 19014
rect 20401 19012 20457 19014
rect 19798 17992 19854 18048
rect 19890 17856 19946 17912
rect 18418 14456 18474 14512
rect 18326 13912 18382 13968
rect 18878 13912 18934 13968
rect 18510 13268 18512 13288
rect 18512 13268 18564 13288
rect 18564 13268 18566 13288
rect 18510 13232 18566 13268
rect 18786 13096 18842 13152
rect 18878 12416 18934 12472
rect 19614 16224 19670 16280
rect 19614 15816 19670 15872
rect 19798 16904 19854 16960
rect 21362 22072 21418 22128
rect 21914 25336 21970 25392
rect 21914 25064 21970 25120
rect 22374 26424 22430 26480
rect 22190 26152 22246 26208
rect 22374 26016 22430 26072
rect 22558 26016 22614 26072
rect 22466 25880 22522 25936
rect 23294 29416 23350 29472
rect 23018 29280 23074 29336
rect 23202 29280 23258 29336
rect 22926 29008 22982 29064
rect 23110 29008 23166 29064
rect 23294 29028 23350 29064
rect 23294 29008 23296 29028
rect 23296 29008 23348 29028
rect 23348 29008 23350 29028
rect 23110 28872 23166 28928
rect 23754 32136 23810 32192
rect 23846 31628 23848 31648
rect 23848 31628 23900 31648
rect 23900 31628 23902 31648
rect 23846 31592 23902 31628
rect 24002 31578 24058 31580
rect 24082 31578 24138 31580
rect 24162 31578 24218 31580
rect 24242 31578 24298 31580
rect 24002 31526 24048 31578
rect 24048 31526 24058 31578
rect 24082 31526 24112 31578
rect 24112 31526 24124 31578
rect 24124 31526 24138 31578
rect 24162 31526 24176 31578
rect 24176 31526 24188 31578
rect 24188 31526 24218 31578
rect 24242 31526 24252 31578
rect 24252 31526 24298 31578
rect 24002 31524 24058 31526
rect 24082 31524 24138 31526
rect 24162 31524 24218 31526
rect 24242 31524 24298 31526
rect 23846 31476 23902 31512
rect 23846 31456 23848 31476
rect 23848 31456 23900 31476
rect 23900 31456 23902 31476
rect 23662 30776 23718 30832
rect 23754 30504 23810 30560
rect 24490 31592 24546 31648
rect 24490 31476 24546 31512
rect 24490 31456 24492 31476
rect 24492 31456 24544 31476
rect 24544 31456 24546 31476
rect 25134 33224 25190 33280
rect 24950 31592 25006 31648
rect 24766 30776 24822 30832
rect 23754 30368 23810 30424
rect 23754 29416 23810 29472
rect 23662 29280 23718 29336
rect 23662 29164 23718 29200
rect 23662 29144 23664 29164
rect 23664 29144 23716 29164
rect 23716 29144 23718 29164
rect 23570 28872 23626 28928
rect 22926 28056 22982 28112
rect 22834 27512 22890 27568
rect 23018 27512 23074 27568
rect 22926 27376 22982 27432
rect 22742 27240 22798 27296
rect 23018 27240 23074 27296
rect 22926 26988 22982 27024
rect 22926 26968 22928 26988
rect 22928 26968 22980 26988
rect 22980 26968 22982 26988
rect 23570 28364 23572 28384
rect 23572 28364 23624 28384
rect 23624 28364 23626 28384
rect 23570 28328 23626 28364
rect 23662 28212 23718 28248
rect 23662 28192 23664 28212
rect 23664 28192 23716 28212
rect 23716 28192 23718 28212
rect 23202 27512 23258 27568
rect 23386 27512 23442 27568
rect 23294 27376 23350 27432
rect 23570 27920 23626 27976
rect 23754 27376 23810 27432
rect 22190 25336 22246 25392
rect 22006 24928 22062 24984
rect 21638 22616 21694 22672
rect 21638 21800 21694 21856
rect 21638 20848 21694 20904
rect 21638 20576 21694 20632
rect 21086 18536 21142 18592
rect 20161 17978 20217 17980
rect 20241 17978 20297 17980
rect 20321 17978 20377 17980
rect 20401 17978 20457 17980
rect 20161 17926 20207 17978
rect 20207 17926 20217 17978
rect 20241 17926 20271 17978
rect 20271 17926 20283 17978
rect 20283 17926 20297 17978
rect 20321 17926 20335 17978
rect 20335 17926 20347 17978
rect 20347 17926 20377 17978
rect 20401 17926 20411 17978
rect 20411 17926 20457 17978
rect 20161 17924 20217 17926
rect 20241 17924 20297 17926
rect 20321 17924 20377 17926
rect 20401 17924 20457 17926
rect 20626 17584 20682 17640
rect 19982 16768 20038 16824
rect 20161 16890 20217 16892
rect 20241 16890 20297 16892
rect 20321 16890 20377 16892
rect 20401 16890 20457 16892
rect 20161 16838 20207 16890
rect 20207 16838 20217 16890
rect 20241 16838 20271 16890
rect 20271 16838 20283 16890
rect 20283 16838 20297 16890
rect 20321 16838 20335 16890
rect 20335 16838 20347 16890
rect 20347 16838 20377 16890
rect 20401 16838 20411 16890
rect 20411 16838 20457 16890
rect 20161 16836 20217 16838
rect 20241 16836 20297 16838
rect 20321 16836 20377 16838
rect 20401 16836 20457 16838
rect 19890 15680 19946 15736
rect 19430 14592 19486 14648
rect 19154 13504 19210 13560
rect 19062 13232 19118 13288
rect 19338 13368 19394 13424
rect 19706 14592 19762 14648
rect 19614 14048 19670 14104
rect 19522 12008 19578 12064
rect 15750 10376 15806 10432
rect 19890 14048 19946 14104
rect 19798 13096 19854 13152
rect 20534 16632 20590 16688
rect 20161 15802 20217 15804
rect 20241 15802 20297 15804
rect 20321 15802 20377 15804
rect 20401 15802 20457 15804
rect 20161 15750 20207 15802
rect 20207 15750 20217 15802
rect 20241 15750 20271 15802
rect 20271 15750 20283 15802
rect 20283 15750 20297 15802
rect 20321 15750 20335 15802
rect 20335 15750 20347 15802
rect 20347 15750 20377 15802
rect 20401 15750 20411 15802
rect 20411 15750 20457 15802
rect 20161 15748 20217 15750
rect 20241 15748 20297 15750
rect 20321 15748 20377 15750
rect 20401 15748 20457 15750
rect 20718 15136 20774 15192
rect 20810 15000 20866 15056
rect 21178 16496 21234 16552
rect 21086 15680 21142 15736
rect 20994 14864 21050 14920
rect 20161 14714 20217 14716
rect 20241 14714 20297 14716
rect 20321 14714 20377 14716
rect 20401 14714 20457 14716
rect 20161 14662 20207 14714
rect 20207 14662 20217 14714
rect 20241 14662 20271 14714
rect 20271 14662 20283 14714
rect 20283 14662 20297 14714
rect 20321 14662 20335 14714
rect 20335 14662 20347 14714
rect 20347 14662 20377 14714
rect 20401 14662 20411 14714
rect 20411 14662 20457 14714
rect 20161 14660 20217 14662
rect 20241 14660 20297 14662
rect 20321 14660 20377 14662
rect 20401 14660 20457 14662
rect 20350 14456 20406 14512
rect 20534 14320 20590 14376
rect 19982 13640 20038 13696
rect 19890 12552 19946 12608
rect 20161 13626 20217 13628
rect 20241 13626 20297 13628
rect 20321 13626 20377 13628
rect 20401 13626 20457 13628
rect 20161 13574 20207 13626
rect 20207 13574 20217 13626
rect 20241 13574 20271 13626
rect 20271 13574 20283 13626
rect 20283 13574 20297 13626
rect 20321 13574 20335 13626
rect 20335 13574 20347 13626
rect 20347 13574 20377 13626
rect 20401 13574 20411 13626
rect 20411 13574 20457 13626
rect 20161 13572 20217 13574
rect 20241 13572 20297 13574
rect 20321 13572 20377 13574
rect 20401 13572 20457 13574
rect 20534 13096 20590 13152
rect 20161 12538 20217 12540
rect 20241 12538 20297 12540
rect 20321 12538 20377 12540
rect 20401 12538 20457 12540
rect 20161 12486 20207 12538
rect 20207 12486 20217 12538
rect 20241 12486 20271 12538
rect 20271 12486 20283 12538
rect 20283 12486 20297 12538
rect 20321 12486 20335 12538
rect 20335 12486 20347 12538
rect 20347 12486 20377 12538
rect 20401 12486 20411 12538
rect 20411 12486 20457 12538
rect 20161 12484 20217 12486
rect 20241 12484 20297 12486
rect 20321 12484 20377 12486
rect 20401 12484 20457 12486
rect 19982 12008 20038 12064
rect 19982 11464 20038 11520
rect 20161 11450 20217 11452
rect 20241 11450 20297 11452
rect 20321 11450 20377 11452
rect 20401 11450 20457 11452
rect 20161 11398 20207 11450
rect 20207 11398 20217 11450
rect 20241 11398 20271 11450
rect 20271 11398 20283 11450
rect 20283 11398 20297 11450
rect 20321 11398 20335 11450
rect 20335 11398 20347 11450
rect 20347 11398 20377 11450
rect 20401 11398 20411 11450
rect 20411 11398 20457 11450
rect 20161 11396 20217 11398
rect 20241 11396 20297 11398
rect 20321 11396 20377 11398
rect 20401 11396 20457 11398
rect 20810 13232 20866 13288
rect 20902 10804 20958 10840
rect 20902 10784 20904 10804
rect 20904 10784 20956 10804
rect 20956 10784 20958 10804
rect 20902 10668 20958 10704
rect 20902 10648 20904 10668
rect 20904 10648 20956 10668
rect 20956 10648 20958 10668
rect 19706 10376 19762 10432
rect 20161 10362 20217 10364
rect 20241 10362 20297 10364
rect 20321 10362 20377 10364
rect 20401 10362 20457 10364
rect 20161 10310 20207 10362
rect 20207 10310 20217 10362
rect 20241 10310 20271 10362
rect 20271 10310 20283 10362
rect 20283 10310 20297 10362
rect 20321 10310 20335 10362
rect 20335 10310 20347 10362
rect 20347 10310 20377 10362
rect 20401 10310 20411 10362
rect 20411 10310 20457 10362
rect 20161 10308 20217 10310
rect 20241 10308 20297 10310
rect 20321 10308 20377 10310
rect 20401 10308 20457 10310
rect 20902 10240 20958 10296
rect 21454 17720 21510 17776
rect 22006 24792 22062 24848
rect 22190 24792 22246 24848
rect 22558 25200 22614 25256
rect 22190 24384 22246 24440
rect 22374 24384 22430 24440
rect 22098 23704 22154 23760
rect 21822 23160 21878 23216
rect 22006 23160 22062 23216
rect 22466 24112 22522 24168
rect 22006 22888 22062 22944
rect 22006 22072 22062 22128
rect 22190 21664 22246 21720
rect 22374 22888 22430 22944
rect 22650 23976 22706 24032
rect 23662 27240 23718 27296
rect 23754 26968 23810 27024
rect 24002 30490 24058 30492
rect 24082 30490 24138 30492
rect 24162 30490 24218 30492
rect 24242 30490 24298 30492
rect 24002 30438 24048 30490
rect 24048 30438 24058 30490
rect 24082 30438 24112 30490
rect 24112 30438 24124 30490
rect 24124 30438 24138 30490
rect 24162 30438 24176 30490
rect 24176 30438 24188 30490
rect 24188 30438 24218 30490
rect 24242 30438 24252 30490
rect 24252 30438 24298 30490
rect 24002 30436 24058 30438
rect 24082 30436 24138 30438
rect 24162 30436 24218 30438
rect 24242 30436 24298 30438
rect 23938 29960 23994 30016
rect 24002 29402 24058 29404
rect 24082 29402 24138 29404
rect 24162 29402 24218 29404
rect 24242 29402 24298 29404
rect 24002 29350 24048 29402
rect 24048 29350 24058 29402
rect 24082 29350 24112 29402
rect 24112 29350 24124 29402
rect 24124 29350 24138 29402
rect 24162 29350 24176 29402
rect 24176 29350 24188 29402
rect 24188 29350 24218 29402
rect 24242 29350 24252 29402
rect 24252 29350 24298 29402
rect 24002 29348 24058 29350
rect 24082 29348 24138 29350
rect 24162 29348 24218 29350
rect 24242 29348 24298 29350
rect 24214 29144 24270 29200
rect 23938 28872 23994 28928
rect 24490 30368 24546 30424
rect 24306 29028 24362 29064
rect 24306 29008 24308 29028
rect 24308 29008 24360 29028
rect 24360 29008 24362 29028
rect 24002 28314 24058 28316
rect 24082 28314 24138 28316
rect 24162 28314 24218 28316
rect 24242 28314 24298 28316
rect 24002 28262 24048 28314
rect 24048 28262 24058 28314
rect 24082 28262 24112 28314
rect 24112 28262 24124 28314
rect 24124 28262 24138 28314
rect 24162 28262 24176 28314
rect 24176 28262 24188 28314
rect 24188 28262 24218 28314
rect 24242 28262 24252 28314
rect 24252 28262 24298 28314
rect 24002 28260 24058 28262
rect 24082 28260 24138 28262
rect 24162 28260 24218 28262
rect 24242 28260 24298 28262
rect 24306 27920 24362 27976
rect 24122 27784 24178 27840
rect 24030 27512 24086 27568
rect 24122 27376 24178 27432
rect 24002 27226 24058 27228
rect 24082 27226 24138 27228
rect 24162 27226 24218 27228
rect 24242 27226 24298 27228
rect 24002 27174 24048 27226
rect 24048 27174 24058 27226
rect 24082 27174 24112 27226
rect 24112 27174 24124 27226
rect 24124 27174 24138 27226
rect 24162 27174 24176 27226
rect 24176 27174 24188 27226
rect 24188 27174 24218 27226
rect 24242 27174 24252 27226
rect 24252 27174 24298 27226
rect 24002 27172 24058 27174
rect 24082 27172 24138 27174
rect 24162 27172 24218 27174
rect 24242 27172 24298 27174
rect 23662 26560 23718 26616
rect 22926 24112 22982 24168
rect 22834 23976 22890 24032
rect 22742 23840 22798 23896
rect 22742 23704 22798 23760
rect 23202 23840 23258 23896
rect 22742 22616 22798 22672
rect 21822 21256 21878 21312
rect 22006 20304 22062 20360
rect 22190 21120 22246 21176
rect 22466 20712 22522 20768
rect 22282 20440 22338 20496
rect 22374 20168 22430 20224
rect 22006 19896 22062 19952
rect 22098 19624 22154 19680
rect 21730 17992 21786 18048
rect 21546 15136 21602 15192
rect 21546 14728 21602 14784
rect 21362 13096 21418 13152
rect 21546 13640 21602 13696
rect 21546 12824 21602 12880
rect 21546 12552 21602 12608
rect 21454 12416 21510 12472
rect 21454 11600 21510 11656
rect 21730 13232 21786 13288
rect 21730 12552 21786 12608
rect 22282 16768 22338 16824
rect 22466 16940 22468 16960
rect 22468 16940 22520 16960
rect 22520 16940 22522 16960
rect 22466 16904 22522 16940
rect 22742 19896 22798 19952
rect 22926 22344 22982 22400
rect 23110 22380 23112 22400
rect 23112 22380 23164 22400
rect 23164 22380 23166 22400
rect 23110 22344 23166 22380
rect 23386 25336 23442 25392
rect 23846 26560 23902 26616
rect 24030 26968 24086 27024
rect 24122 26560 24178 26616
rect 24306 26868 24308 26888
rect 24308 26868 24360 26888
rect 24360 26868 24362 26888
rect 24306 26832 24362 26868
rect 24214 26288 24270 26344
rect 24002 26138 24058 26140
rect 24082 26138 24138 26140
rect 24162 26138 24218 26140
rect 24242 26138 24298 26140
rect 24002 26086 24048 26138
rect 24048 26086 24058 26138
rect 24082 26086 24112 26138
rect 24112 26086 24124 26138
rect 24124 26086 24138 26138
rect 24162 26086 24176 26138
rect 24176 26086 24188 26138
rect 24188 26086 24218 26138
rect 24242 26086 24252 26138
rect 24252 26086 24298 26138
rect 24002 26084 24058 26086
rect 24082 26084 24138 26086
rect 24162 26084 24218 26086
rect 24242 26084 24298 26086
rect 23662 25336 23718 25392
rect 23570 25200 23626 25256
rect 23570 24928 23626 24984
rect 23478 24384 23534 24440
rect 23386 23976 23442 24032
rect 24214 25744 24270 25800
rect 24122 25492 24178 25528
rect 24122 25472 24124 25492
rect 24124 25472 24176 25492
rect 24176 25472 24178 25492
rect 24030 25200 24086 25256
rect 24306 25336 24362 25392
rect 24950 30504 25006 30560
rect 24950 30096 25006 30152
rect 24766 29824 24822 29880
rect 24674 29688 24730 29744
rect 24674 29280 24730 29336
rect 24858 29688 24914 29744
rect 24766 29144 24822 29200
rect 24582 28192 24638 28248
rect 24674 27784 24730 27840
rect 24582 27648 24638 27704
rect 24674 27376 24730 27432
rect 24490 25472 24546 25528
rect 24950 29416 25006 29472
rect 24950 29164 25006 29200
rect 24950 29144 24952 29164
rect 24952 29144 25004 29164
rect 25004 29144 25006 29164
rect 25226 31320 25282 31376
rect 25226 30368 25282 30424
rect 25410 31864 25466 31920
rect 25502 31084 25504 31104
rect 25504 31084 25556 31104
rect 25556 31084 25558 31104
rect 25502 31048 25558 31084
rect 25226 30132 25228 30152
rect 25228 30132 25280 30152
rect 25280 30132 25282 30152
rect 25226 30096 25282 30132
rect 25226 29688 25282 29744
rect 25226 29416 25282 29472
rect 24766 26016 24822 26072
rect 24950 26560 25006 26616
rect 25226 27820 25228 27840
rect 25228 27820 25280 27840
rect 25280 27820 25282 27840
rect 25226 27784 25282 27820
rect 25594 29416 25650 29472
rect 26790 34040 26846 34096
rect 26146 30776 26202 30832
rect 25778 29552 25834 29608
rect 25410 27784 25466 27840
rect 25318 27648 25374 27704
rect 25134 27104 25190 27160
rect 25134 26832 25190 26888
rect 25042 26288 25098 26344
rect 24950 25608 25006 25664
rect 24490 25200 24546 25256
rect 24766 25336 24822 25392
rect 24398 25064 24454 25120
rect 24002 25050 24058 25052
rect 24082 25050 24138 25052
rect 24162 25050 24218 25052
rect 24242 25050 24298 25052
rect 24002 24998 24048 25050
rect 24048 24998 24058 25050
rect 24082 24998 24112 25050
rect 24112 24998 24124 25050
rect 24124 24998 24138 25050
rect 24162 24998 24176 25050
rect 24176 24998 24188 25050
rect 24188 24998 24218 25050
rect 24242 24998 24252 25050
rect 24252 24998 24298 25050
rect 24002 24996 24058 24998
rect 24082 24996 24138 24998
rect 24162 24996 24218 24998
rect 24242 24996 24298 24998
rect 24398 24928 24454 24984
rect 23846 23976 23902 24032
rect 23570 23840 23626 23896
rect 23754 23840 23810 23896
rect 23478 23604 23480 23624
rect 23480 23604 23532 23624
rect 23532 23604 23534 23624
rect 23478 23568 23534 23604
rect 23478 23432 23534 23488
rect 23478 22480 23534 22536
rect 23570 21256 23626 21312
rect 24002 23962 24058 23964
rect 24082 23962 24138 23964
rect 24162 23962 24218 23964
rect 24242 23962 24298 23964
rect 24002 23910 24048 23962
rect 24048 23910 24058 23962
rect 24082 23910 24112 23962
rect 24112 23910 24124 23962
rect 24124 23910 24138 23962
rect 24162 23910 24176 23962
rect 24176 23910 24188 23962
rect 24188 23910 24218 23962
rect 24242 23910 24252 23962
rect 24252 23910 24298 23962
rect 24002 23908 24058 23910
rect 24082 23908 24138 23910
rect 24162 23908 24218 23910
rect 24242 23908 24298 23910
rect 24766 24656 24822 24712
rect 24490 23840 24546 23896
rect 24398 23296 24454 23352
rect 25042 24556 25044 24576
rect 25044 24556 25096 24576
rect 25096 24556 25098 24576
rect 25042 24520 25098 24556
rect 25226 24520 25282 24576
rect 24582 22888 24638 22944
rect 24002 22874 24058 22876
rect 24082 22874 24138 22876
rect 24162 22874 24218 22876
rect 24242 22874 24298 22876
rect 24002 22822 24048 22874
rect 24048 22822 24058 22874
rect 24082 22822 24112 22874
rect 24112 22822 24124 22874
rect 24124 22822 24138 22874
rect 24162 22822 24176 22874
rect 24176 22822 24188 22874
rect 24188 22822 24218 22874
rect 24242 22822 24252 22874
rect 24252 22822 24298 22874
rect 24002 22820 24058 22822
rect 24082 22820 24138 22822
rect 24162 22820 24218 22822
rect 24242 22820 24298 22822
rect 25226 23704 25282 23760
rect 25778 28620 25834 28656
rect 25778 28600 25780 28620
rect 25780 28600 25832 28620
rect 25832 28600 25834 28620
rect 25594 27820 25596 27840
rect 25596 27820 25648 27840
rect 25648 27820 25650 27840
rect 25594 27784 25650 27820
rect 25778 27784 25834 27840
rect 25502 26152 25558 26208
rect 23938 22208 23994 22264
rect 24002 21786 24058 21788
rect 24082 21786 24138 21788
rect 24162 21786 24218 21788
rect 24242 21786 24298 21788
rect 24002 21734 24048 21786
rect 24048 21734 24058 21786
rect 24082 21734 24112 21786
rect 24112 21734 24124 21786
rect 24124 21734 24138 21786
rect 24162 21734 24176 21786
rect 24176 21734 24188 21786
rect 24188 21734 24218 21786
rect 24242 21734 24252 21786
rect 24252 21734 24298 21786
rect 24002 21732 24058 21734
rect 24082 21732 24138 21734
rect 24162 21732 24218 21734
rect 24242 21732 24298 21734
rect 24674 21800 24730 21856
rect 24582 21664 24638 21720
rect 24490 21256 24546 21312
rect 24002 20698 24058 20700
rect 24082 20698 24138 20700
rect 24162 20698 24218 20700
rect 24242 20698 24298 20700
rect 24002 20646 24048 20698
rect 24048 20646 24058 20698
rect 24082 20646 24112 20698
rect 24112 20646 24124 20698
rect 24124 20646 24138 20698
rect 24162 20646 24176 20698
rect 24176 20646 24188 20698
rect 24188 20646 24218 20698
rect 24242 20646 24252 20698
rect 24252 20646 24298 20698
rect 24002 20644 24058 20646
rect 24082 20644 24138 20646
rect 24162 20644 24218 20646
rect 24242 20644 24298 20646
rect 23110 18944 23166 19000
rect 23110 18672 23166 18728
rect 23018 18536 23074 18592
rect 22742 18300 22744 18320
rect 22744 18300 22796 18320
rect 22796 18300 22798 18320
rect 22742 18264 22798 18300
rect 22374 16632 22430 16688
rect 22282 16124 22284 16144
rect 22284 16124 22336 16144
rect 22336 16124 22338 16144
rect 22282 16088 22338 16124
rect 22098 13368 22154 13424
rect 22466 15000 22522 15056
rect 22466 13776 22522 13832
rect 22374 13232 22430 13288
rect 22282 10784 22338 10840
rect 22742 16632 22798 16688
rect 23018 16632 23074 16688
rect 23018 16496 23074 16552
rect 23202 17720 23258 17776
rect 23202 17040 23258 17096
rect 23570 19488 23626 19544
rect 23386 18672 23442 18728
rect 23386 17176 23442 17232
rect 24002 19610 24058 19612
rect 24082 19610 24138 19612
rect 24162 19610 24218 19612
rect 24242 19610 24298 19612
rect 24002 19558 24048 19610
rect 24048 19558 24058 19610
rect 24082 19558 24112 19610
rect 24112 19558 24124 19610
rect 24124 19558 24138 19610
rect 24162 19558 24176 19610
rect 24176 19558 24188 19610
rect 24188 19558 24218 19610
rect 24242 19558 24252 19610
rect 24252 19558 24298 19610
rect 24002 19556 24058 19558
rect 24082 19556 24138 19558
rect 24162 19556 24218 19558
rect 24242 19556 24298 19558
rect 24582 19488 24638 19544
rect 23662 17992 23718 18048
rect 23570 17312 23626 17368
rect 23754 16768 23810 16824
rect 23294 15952 23350 16008
rect 16320 9818 16376 9820
rect 16400 9818 16456 9820
rect 16480 9818 16536 9820
rect 16560 9818 16616 9820
rect 16320 9766 16366 9818
rect 16366 9766 16376 9818
rect 16400 9766 16430 9818
rect 16430 9766 16442 9818
rect 16442 9766 16456 9818
rect 16480 9766 16494 9818
rect 16494 9766 16506 9818
rect 16506 9766 16536 9818
rect 16560 9766 16570 9818
rect 16570 9766 16616 9818
rect 16320 9764 16376 9766
rect 16400 9764 16456 9766
rect 16480 9764 16536 9766
rect 16560 9764 16616 9766
rect 22190 10376 22246 10432
rect 23662 16088 23718 16144
rect 23478 14320 23534 14376
rect 23570 13640 23626 13696
rect 23570 11892 23626 11928
rect 23570 11872 23572 11892
rect 23572 11872 23624 11892
rect 23624 11872 23626 11892
rect 23202 10376 23258 10432
rect 24030 19116 24032 19136
rect 24032 19116 24084 19136
rect 24084 19116 24086 19136
rect 24030 19080 24086 19116
rect 24490 18944 24546 19000
rect 24490 18536 24546 18592
rect 24002 18522 24058 18524
rect 24082 18522 24138 18524
rect 24162 18522 24218 18524
rect 24242 18522 24298 18524
rect 24002 18470 24048 18522
rect 24048 18470 24058 18522
rect 24082 18470 24112 18522
rect 24112 18470 24124 18522
rect 24124 18470 24138 18522
rect 24162 18470 24176 18522
rect 24176 18470 24188 18522
rect 24188 18470 24218 18522
rect 24242 18470 24252 18522
rect 24252 18470 24298 18522
rect 24002 18468 24058 18470
rect 24082 18468 24138 18470
rect 24162 18468 24218 18470
rect 24242 18468 24298 18470
rect 24398 18400 24454 18456
rect 24002 17434 24058 17436
rect 24082 17434 24138 17436
rect 24162 17434 24218 17436
rect 24242 17434 24298 17436
rect 24002 17382 24048 17434
rect 24048 17382 24058 17434
rect 24082 17382 24112 17434
rect 24112 17382 24124 17434
rect 24124 17382 24138 17434
rect 24162 17382 24176 17434
rect 24176 17382 24188 17434
rect 24188 17382 24218 17434
rect 24242 17382 24252 17434
rect 24252 17382 24298 17434
rect 24002 17380 24058 17382
rect 24082 17380 24138 17382
rect 24162 17380 24218 17382
rect 24242 17380 24298 17382
rect 24030 16496 24086 16552
rect 24002 16346 24058 16348
rect 24082 16346 24138 16348
rect 24162 16346 24218 16348
rect 24242 16346 24298 16348
rect 24002 16294 24048 16346
rect 24048 16294 24058 16346
rect 24082 16294 24112 16346
rect 24112 16294 24124 16346
rect 24124 16294 24138 16346
rect 24162 16294 24176 16346
rect 24176 16294 24188 16346
rect 24188 16294 24218 16346
rect 24242 16294 24252 16346
rect 24252 16294 24298 16346
rect 24002 16292 24058 16294
rect 24082 16292 24138 16294
rect 24162 16292 24218 16294
rect 24242 16292 24298 16294
rect 23938 15544 23994 15600
rect 24030 15408 24086 15464
rect 24002 15258 24058 15260
rect 24082 15258 24138 15260
rect 24162 15258 24218 15260
rect 24242 15258 24298 15260
rect 24002 15206 24048 15258
rect 24048 15206 24058 15258
rect 24082 15206 24112 15258
rect 24112 15206 24124 15258
rect 24124 15206 24138 15258
rect 24162 15206 24176 15258
rect 24176 15206 24188 15258
rect 24188 15206 24218 15258
rect 24242 15206 24252 15258
rect 24252 15206 24298 15258
rect 24002 15204 24058 15206
rect 24082 15204 24138 15206
rect 24162 15204 24218 15206
rect 24242 15204 24298 15206
rect 23846 14592 23902 14648
rect 24002 14170 24058 14172
rect 24082 14170 24138 14172
rect 24162 14170 24218 14172
rect 24242 14170 24298 14172
rect 24002 14118 24048 14170
rect 24048 14118 24058 14170
rect 24082 14118 24112 14170
rect 24112 14118 24124 14170
rect 24124 14118 24138 14170
rect 24162 14118 24176 14170
rect 24176 14118 24188 14170
rect 24188 14118 24218 14170
rect 24242 14118 24252 14170
rect 24252 14118 24298 14170
rect 24002 14116 24058 14118
rect 24082 14116 24138 14118
rect 24162 14116 24218 14118
rect 24242 14116 24298 14118
rect 24490 18128 24546 18184
rect 24858 19352 24914 19408
rect 24766 17992 24822 18048
rect 24490 15680 24546 15736
rect 24766 17584 24822 17640
rect 26514 30912 26570 30968
rect 26330 30504 26386 30560
rect 26054 29960 26110 30016
rect 26146 29552 26202 29608
rect 26330 29960 26386 30016
rect 26146 29416 26202 29472
rect 26238 29280 26294 29336
rect 26238 28328 26294 28384
rect 26146 27784 26202 27840
rect 26238 27548 26240 27568
rect 26240 27548 26292 27568
rect 26292 27548 26294 27568
rect 26238 27512 26294 27548
rect 25962 27104 26018 27160
rect 25870 26852 25926 26888
rect 25870 26832 25872 26852
rect 25872 26832 25924 26852
rect 25924 26832 25926 26852
rect 25686 26152 25742 26208
rect 25870 26016 25926 26072
rect 25594 25880 25650 25936
rect 25594 24384 25650 24440
rect 25502 23976 25558 24032
rect 25410 23160 25466 23216
rect 25226 22344 25282 22400
rect 25318 22072 25374 22128
rect 25226 20984 25282 21040
rect 25042 19760 25098 19816
rect 25042 19352 25098 19408
rect 24858 17448 24914 17504
rect 24674 17312 24730 17368
rect 24674 16768 24730 16824
rect 24858 17176 24914 17232
rect 24858 16360 24914 16416
rect 24858 15952 24914 16008
rect 24490 14592 24546 14648
rect 24030 13776 24086 13832
rect 24858 14048 24914 14104
rect 24858 13912 24914 13968
rect 24766 13796 24822 13832
rect 24766 13776 24768 13796
rect 24768 13776 24820 13796
rect 24820 13776 24822 13796
rect 24582 13368 24638 13424
rect 23846 13096 23902 13152
rect 24002 13082 24058 13084
rect 24082 13082 24138 13084
rect 24162 13082 24218 13084
rect 24242 13082 24298 13084
rect 24002 13030 24048 13082
rect 24048 13030 24058 13082
rect 24082 13030 24112 13082
rect 24112 13030 24124 13082
rect 24124 13030 24138 13082
rect 24162 13030 24176 13082
rect 24176 13030 24188 13082
rect 24188 13030 24218 13082
rect 24242 13030 24252 13082
rect 24252 13030 24298 13082
rect 24002 13028 24058 13030
rect 24082 13028 24138 13030
rect 24162 13028 24218 13030
rect 24242 13028 24298 13030
rect 24214 12844 24270 12880
rect 24214 12824 24216 12844
rect 24216 12824 24268 12844
rect 24268 12824 24270 12844
rect 23846 12416 23902 12472
rect 24002 11994 24058 11996
rect 24082 11994 24138 11996
rect 24162 11994 24218 11996
rect 24242 11994 24298 11996
rect 24002 11942 24048 11994
rect 24048 11942 24058 11994
rect 24082 11942 24112 11994
rect 24112 11942 24124 11994
rect 24124 11942 24138 11994
rect 24162 11942 24176 11994
rect 24176 11942 24188 11994
rect 24188 11942 24218 11994
rect 24242 11942 24252 11994
rect 24252 11942 24298 11994
rect 24002 11940 24058 11942
rect 24082 11940 24138 11942
rect 24162 11940 24218 11942
rect 24242 11940 24298 11942
rect 24002 10906 24058 10908
rect 24082 10906 24138 10908
rect 24162 10906 24218 10908
rect 24242 10906 24298 10908
rect 24002 10854 24048 10906
rect 24048 10854 24058 10906
rect 24082 10854 24112 10906
rect 24112 10854 24124 10906
rect 24124 10854 24138 10906
rect 24162 10854 24176 10906
rect 24176 10854 24188 10906
rect 24188 10854 24218 10906
rect 24242 10854 24252 10906
rect 24252 10854 24298 10906
rect 24002 10852 24058 10854
rect 24082 10852 24138 10854
rect 24162 10852 24218 10854
rect 24242 10852 24298 10854
rect 24306 10648 24362 10704
rect 23846 10376 23902 10432
rect 20161 9274 20217 9276
rect 20241 9274 20297 9276
rect 20321 9274 20377 9276
rect 20401 9274 20457 9276
rect 20161 9222 20207 9274
rect 20207 9222 20217 9274
rect 20241 9222 20271 9274
rect 20271 9222 20283 9274
rect 20283 9222 20297 9274
rect 20321 9222 20335 9274
rect 20335 9222 20347 9274
rect 20347 9222 20377 9274
rect 20401 9222 20411 9274
rect 20411 9222 20457 9274
rect 20161 9220 20217 9222
rect 20241 9220 20297 9222
rect 20321 9220 20377 9222
rect 20401 9220 20457 9222
rect 16320 8730 16376 8732
rect 16400 8730 16456 8732
rect 16480 8730 16536 8732
rect 16560 8730 16616 8732
rect 16320 8678 16366 8730
rect 16366 8678 16376 8730
rect 16400 8678 16430 8730
rect 16430 8678 16442 8730
rect 16442 8678 16456 8730
rect 16480 8678 16494 8730
rect 16494 8678 16506 8730
rect 16506 8678 16536 8730
rect 16560 8678 16570 8730
rect 16570 8678 16616 8730
rect 16320 8676 16376 8678
rect 16400 8676 16456 8678
rect 16480 8676 16536 8678
rect 16560 8676 16616 8678
rect 19522 8608 19578 8664
rect 25042 16360 25098 16416
rect 25042 15272 25098 15328
rect 25042 12960 25098 13016
rect 25870 25880 25926 25936
rect 26146 27412 26148 27432
rect 26148 27412 26200 27432
rect 26200 27412 26202 27432
rect 26146 27376 26202 27412
rect 26514 29416 26570 29472
rect 26514 29008 26570 29064
rect 27066 32408 27122 32464
rect 29090 34312 29146 34368
rect 26790 30776 26846 30832
rect 26790 29824 26846 29880
rect 26606 28872 26662 28928
rect 26606 28736 26662 28792
rect 26790 28908 26792 28928
rect 26792 28908 26844 28928
rect 26844 28908 26846 28928
rect 26790 28872 26846 28908
rect 26790 28736 26846 28792
rect 27434 32136 27490 32192
rect 27066 31184 27122 31240
rect 27066 29996 27068 30016
rect 27068 29996 27120 30016
rect 27120 29996 27122 30016
rect 27066 29960 27122 29996
rect 27066 29416 27122 29472
rect 26422 28192 26478 28248
rect 26422 27920 26478 27976
rect 26606 28328 26662 28384
rect 26790 28192 26846 28248
rect 26790 27920 26846 27976
rect 26514 27784 26570 27840
rect 26790 27820 26792 27840
rect 26792 27820 26844 27840
rect 26844 27820 26846 27840
rect 26790 27784 26846 27820
rect 26974 27648 27030 27704
rect 26422 27240 26478 27296
rect 26238 26832 26294 26888
rect 25778 25064 25834 25120
rect 25962 24792 26018 24848
rect 25870 24656 25926 24712
rect 25870 24384 25926 24440
rect 25686 24112 25742 24168
rect 25686 23740 25688 23760
rect 25688 23740 25740 23760
rect 25740 23740 25742 23760
rect 25686 23704 25742 23740
rect 25870 23568 25926 23624
rect 27066 27512 27122 27568
rect 26974 27104 27030 27160
rect 26698 26832 26754 26888
rect 26514 25780 26516 25800
rect 26516 25780 26568 25800
rect 26568 25780 26570 25800
rect 26514 25744 26570 25780
rect 26514 25608 26570 25664
rect 26422 24928 26478 24984
rect 26330 23568 26386 23624
rect 25594 23160 25650 23216
rect 25502 20576 25558 20632
rect 25778 20984 25834 21040
rect 26790 26152 26846 26208
rect 26698 25064 26754 25120
rect 26698 24520 26754 24576
rect 26790 24112 26846 24168
rect 26606 23840 26662 23896
rect 27066 26560 27122 26616
rect 27342 31084 27344 31104
rect 27344 31084 27396 31104
rect 27396 31084 27398 31104
rect 27342 31048 27398 31084
rect 27342 30640 27398 30696
rect 27342 29824 27398 29880
rect 27434 29416 27490 29472
rect 27526 29280 27582 29336
rect 27843 32122 27899 32124
rect 27923 32122 27979 32124
rect 28003 32122 28059 32124
rect 28083 32122 28139 32124
rect 27843 32070 27889 32122
rect 27889 32070 27899 32122
rect 27923 32070 27953 32122
rect 27953 32070 27965 32122
rect 27965 32070 27979 32122
rect 28003 32070 28017 32122
rect 28017 32070 28029 32122
rect 28029 32070 28059 32122
rect 28083 32070 28093 32122
rect 28093 32070 28139 32122
rect 27843 32068 27899 32070
rect 27923 32068 27979 32070
rect 28003 32068 28059 32070
rect 28083 32068 28139 32070
rect 27710 32000 27766 32056
rect 27843 31034 27899 31036
rect 27923 31034 27979 31036
rect 28003 31034 28059 31036
rect 28083 31034 28139 31036
rect 27843 30982 27889 31034
rect 27889 30982 27899 31034
rect 27923 30982 27953 31034
rect 27953 30982 27965 31034
rect 27965 30982 27979 31034
rect 28003 30982 28017 31034
rect 28017 30982 28029 31034
rect 28029 30982 28059 31034
rect 28083 30982 28093 31034
rect 28093 30982 28139 31034
rect 27843 30980 27899 30982
rect 27923 30980 27979 30982
rect 28003 30980 28059 30982
rect 28083 30980 28139 30982
rect 28354 32292 28410 32328
rect 28354 32272 28356 32292
rect 28356 32272 28408 32292
rect 28408 32272 28410 32292
rect 27894 30368 27950 30424
rect 27843 29946 27899 29948
rect 27923 29946 27979 29948
rect 28003 29946 28059 29948
rect 28083 29946 28139 29948
rect 27843 29894 27889 29946
rect 27889 29894 27899 29946
rect 27923 29894 27953 29946
rect 27953 29894 27965 29946
rect 27965 29894 27979 29946
rect 28003 29894 28017 29946
rect 28017 29894 28029 29946
rect 28029 29894 28059 29946
rect 28083 29894 28093 29946
rect 28093 29894 28139 29946
rect 27843 29892 27899 29894
rect 27923 29892 27979 29894
rect 28003 29892 28059 29894
rect 28083 29892 28139 29894
rect 28078 29688 28134 29744
rect 27986 29552 28042 29608
rect 28722 31048 28778 31104
rect 28446 30912 28502 30968
rect 28354 30776 28410 30832
rect 28354 30368 28410 30424
rect 28446 29824 28502 29880
rect 28262 29688 28318 29744
rect 28262 29416 28318 29472
rect 27526 28736 27582 28792
rect 28262 28872 28318 28928
rect 27843 28858 27899 28860
rect 27923 28858 27979 28860
rect 28003 28858 28059 28860
rect 28083 28858 28139 28860
rect 27843 28806 27889 28858
rect 27889 28806 27899 28858
rect 27923 28806 27953 28858
rect 27953 28806 27965 28858
rect 27965 28806 27979 28858
rect 28003 28806 28017 28858
rect 28017 28806 28029 28858
rect 28029 28806 28059 28858
rect 28083 28806 28093 28858
rect 28093 28806 28139 28858
rect 27843 28804 27899 28806
rect 27923 28804 27979 28806
rect 28003 28804 28059 28806
rect 28083 28804 28139 28806
rect 28446 28736 28502 28792
rect 28446 28328 28502 28384
rect 27710 27784 27766 27840
rect 28258 27784 28314 27840
rect 27618 27648 27674 27704
rect 27843 27770 27899 27772
rect 27923 27770 27979 27772
rect 28003 27770 28059 27772
rect 28083 27770 28139 27772
rect 27843 27718 27889 27770
rect 27889 27718 27899 27770
rect 27923 27718 27953 27770
rect 27953 27718 27965 27770
rect 27965 27718 27979 27770
rect 28003 27718 28017 27770
rect 28017 27718 28029 27770
rect 28029 27718 28059 27770
rect 28083 27718 28093 27770
rect 28093 27718 28139 27770
rect 27843 27716 27899 27718
rect 27923 27716 27979 27718
rect 28003 27716 28059 27718
rect 28083 27716 28139 27718
rect 27894 27512 27950 27568
rect 27526 27104 27582 27160
rect 27526 26288 27582 26344
rect 27986 27124 28042 27160
rect 27986 27104 27988 27124
rect 27988 27104 28040 27124
rect 28040 27104 28042 27124
rect 28170 27104 28226 27160
rect 27843 26682 27899 26684
rect 27923 26682 27979 26684
rect 28003 26682 28059 26684
rect 28083 26682 28139 26684
rect 27843 26630 27889 26682
rect 27889 26630 27899 26682
rect 27923 26630 27953 26682
rect 27953 26630 27965 26682
rect 27965 26630 27979 26682
rect 28003 26630 28017 26682
rect 28017 26630 28029 26682
rect 28029 26630 28059 26682
rect 28083 26630 28093 26682
rect 28093 26630 28139 26682
rect 27843 26628 27899 26630
rect 27923 26628 27979 26630
rect 28003 26628 28059 26630
rect 28083 26628 28139 26630
rect 26974 25064 27030 25120
rect 26974 24520 27030 24576
rect 26514 23432 26570 23488
rect 26146 22092 26202 22128
rect 26146 22072 26148 22092
rect 26148 22072 26200 22092
rect 26200 22072 26202 22092
rect 25686 19760 25742 19816
rect 25226 17992 25282 18048
rect 25318 16768 25374 16824
rect 25594 19508 25650 19544
rect 25594 19488 25596 19508
rect 25596 19488 25648 19508
rect 25648 19488 25650 19508
rect 25778 19488 25834 19544
rect 25502 16904 25558 16960
rect 25778 18420 25834 18456
rect 25778 18400 25780 18420
rect 25780 18400 25832 18420
rect 25832 18400 25834 18420
rect 25410 16496 25466 16552
rect 25686 16496 25742 16552
rect 25134 12144 25190 12200
rect 24002 9818 24058 9820
rect 24082 9818 24138 9820
rect 24162 9818 24218 9820
rect 24242 9818 24298 9820
rect 24002 9766 24048 9818
rect 24048 9766 24058 9818
rect 24082 9766 24112 9818
rect 24112 9766 24124 9818
rect 24124 9766 24138 9818
rect 24162 9766 24176 9818
rect 24176 9766 24188 9818
rect 24188 9766 24218 9818
rect 24242 9766 24252 9818
rect 24252 9766 24298 9818
rect 24002 9764 24058 9766
rect 24082 9764 24138 9766
rect 24162 9764 24218 9766
rect 24242 9764 24298 9766
rect 24002 8730 24058 8732
rect 24082 8730 24138 8732
rect 24162 8730 24218 8732
rect 24242 8730 24298 8732
rect 24002 8678 24048 8730
rect 24048 8678 24058 8730
rect 24082 8678 24112 8730
rect 24112 8678 24124 8730
rect 24124 8678 24138 8730
rect 24162 8678 24176 8730
rect 24176 8678 24188 8730
rect 24188 8678 24218 8730
rect 24242 8678 24252 8730
rect 24252 8678 24298 8730
rect 24002 8676 24058 8678
rect 24082 8676 24138 8678
rect 24162 8676 24218 8678
rect 24242 8676 24298 8678
rect 19522 8336 19578 8392
rect 12479 8186 12535 8188
rect 12559 8186 12615 8188
rect 12639 8186 12695 8188
rect 12719 8186 12775 8188
rect 12479 8134 12525 8186
rect 12525 8134 12535 8186
rect 12559 8134 12589 8186
rect 12589 8134 12601 8186
rect 12601 8134 12615 8186
rect 12639 8134 12653 8186
rect 12653 8134 12665 8186
rect 12665 8134 12695 8186
rect 12719 8134 12729 8186
rect 12729 8134 12775 8186
rect 12479 8132 12535 8134
rect 12559 8132 12615 8134
rect 12639 8132 12695 8134
rect 12719 8132 12775 8134
rect 20161 8186 20217 8188
rect 20241 8186 20297 8188
rect 20321 8186 20377 8188
rect 20401 8186 20457 8188
rect 20161 8134 20207 8186
rect 20207 8134 20217 8186
rect 20241 8134 20271 8186
rect 20271 8134 20283 8186
rect 20283 8134 20297 8186
rect 20321 8134 20335 8186
rect 20335 8134 20347 8186
rect 20347 8134 20377 8186
rect 20401 8134 20411 8186
rect 20411 8134 20457 8186
rect 20161 8132 20217 8134
rect 20241 8132 20297 8134
rect 20321 8132 20377 8134
rect 20401 8132 20457 8134
rect 16320 7642 16376 7644
rect 16400 7642 16456 7644
rect 16480 7642 16536 7644
rect 16560 7642 16616 7644
rect 16320 7590 16366 7642
rect 16366 7590 16376 7642
rect 16400 7590 16430 7642
rect 16430 7590 16442 7642
rect 16442 7590 16456 7642
rect 16480 7590 16494 7642
rect 16494 7590 16506 7642
rect 16506 7590 16536 7642
rect 16560 7590 16570 7642
rect 16570 7590 16616 7642
rect 16320 7588 16376 7590
rect 16400 7588 16456 7590
rect 16480 7588 16536 7590
rect 16560 7588 16616 7590
rect 24002 7642 24058 7644
rect 24082 7642 24138 7644
rect 24162 7642 24218 7644
rect 24242 7642 24298 7644
rect 24002 7590 24048 7642
rect 24048 7590 24058 7642
rect 24082 7590 24112 7642
rect 24112 7590 24124 7642
rect 24124 7590 24138 7642
rect 24162 7590 24176 7642
rect 24176 7590 24188 7642
rect 24188 7590 24218 7642
rect 24242 7590 24252 7642
rect 24252 7590 24298 7642
rect 24002 7588 24058 7590
rect 24082 7588 24138 7590
rect 24162 7588 24218 7590
rect 24242 7588 24298 7590
rect 12479 7098 12535 7100
rect 12559 7098 12615 7100
rect 12639 7098 12695 7100
rect 12719 7098 12775 7100
rect 12479 7046 12525 7098
rect 12525 7046 12535 7098
rect 12559 7046 12589 7098
rect 12589 7046 12601 7098
rect 12601 7046 12615 7098
rect 12639 7046 12653 7098
rect 12653 7046 12665 7098
rect 12665 7046 12695 7098
rect 12719 7046 12729 7098
rect 12729 7046 12775 7098
rect 12479 7044 12535 7046
rect 12559 7044 12615 7046
rect 12639 7044 12695 7046
rect 12719 7044 12775 7046
rect 20161 7098 20217 7100
rect 20241 7098 20297 7100
rect 20321 7098 20377 7100
rect 20401 7098 20457 7100
rect 20161 7046 20207 7098
rect 20207 7046 20217 7098
rect 20241 7046 20271 7098
rect 20271 7046 20283 7098
rect 20283 7046 20297 7098
rect 20321 7046 20335 7098
rect 20335 7046 20347 7098
rect 20347 7046 20377 7098
rect 20401 7046 20411 7098
rect 20411 7046 20457 7098
rect 20161 7044 20217 7046
rect 20241 7044 20297 7046
rect 20321 7044 20377 7046
rect 20401 7044 20457 7046
rect 8638 6554 8694 6556
rect 8718 6554 8774 6556
rect 8798 6554 8854 6556
rect 8878 6554 8934 6556
rect 8638 6502 8684 6554
rect 8684 6502 8694 6554
rect 8718 6502 8748 6554
rect 8748 6502 8760 6554
rect 8760 6502 8774 6554
rect 8798 6502 8812 6554
rect 8812 6502 8824 6554
rect 8824 6502 8854 6554
rect 8878 6502 8888 6554
rect 8888 6502 8934 6554
rect 8638 6500 8694 6502
rect 8718 6500 8774 6502
rect 8798 6500 8854 6502
rect 8878 6500 8934 6502
rect 8638 5466 8694 5468
rect 8718 5466 8774 5468
rect 8798 5466 8854 5468
rect 8878 5466 8934 5468
rect 8638 5414 8684 5466
rect 8684 5414 8694 5466
rect 8718 5414 8748 5466
rect 8748 5414 8760 5466
rect 8760 5414 8774 5466
rect 8798 5414 8812 5466
rect 8812 5414 8824 5466
rect 8824 5414 8854 5466
rect 8878 5414 8888 5466
rect 8888 5414 8934 5466
rect 8638 5412 8694 5414
rect 8718 5412 8774 5414
rect 8798 5412 8854 5414
rect 8878 5412 8934 5414
rect 16320 6554 16376 6556
rect 16400 6554 16456 6556
rect 16480 6554 16536 6556
rect 16560 6554 16616 6556
rect 16320 6502 16366 6554
rect 16366 6502 16376 6554
rect 16400 6502 16430 6554
rect 16430 6502 16442 6554
rect 16442 6502 16456 6554
rect 16480 6502 16494 6554
rect 16494 6502 16506 6554
rect 16506 6502 16536 6554
rect 16560 6502 16570 6554
rect 16570 6502 16616 6554
rect 16320 6500 16376 6502
rect 16400 6500 16456 6502
rect 16480 6500 16536 6502
rect 16560 6500 16616 6502
rect 24002 6554 24058 6556
rect 24082 6554 24138 6556
rect 24162 6554 24218 6556
rect 24242 6554 24298 6556
rect 24002 6502 24048 6554
rect 24048 6502 24058 6554
rect 24082 6502 24112 6554
rect 24112 6502 24124 6554
rect 24124 6502 24138 6554
rect 24162 6502 24176 6554
rect 24176 6502 24188 6554
rect 24188 6502 24218 6554
rect 24242 6502 24252 6554
rect 24252 6502 24298 6554
rect 24002 6500 24058 6502
rect 24082 6500 24138 6502
rect 24162 6500 24218 6502
rect 24242 6500 24298 6502
rect 12479 6010 12535 6012
rect 12559 6010 12615 6012
rect 12639 6010 12695 6012
rect 12719 6010 12775 6012
rect 12479 5958 12525 6010
rect 12525 5958 12535 6010
rect 12559 5958 12589 6010
rect 12589 5958 12601 6010
rect 12601 5958 12615 6010
rect 12639 5958 12653 6010
rect 12653 5958 12665 6010
rect 12665 5958 12695 6010
rect 12719 5958 12729 6010
rect 12729 5958 12775 6010
rect 12479 5956 12535 5958
rect 12559 5956 12615 5958
rect 12639 5956 12695 5958
rect 12719 5956 12775 5958
rect 20161 6010 20217 6012
rect 20241 6010 20297 6012
rect 20321 6010 20377 6012
rect 20401 6010 20457 6012
rect 20161 5958 20207 6010
rect 20207 5958 20217 6010
rect 20241 5958 20271 6010
rect 20271 5958 20283 6010
rect 20283 5958 20297 6010
rect 20321 5958 20335 6010
rect 20335 5958 20347 6010
rect 20347 5958 20377 6010
rect 20401 5958 20411 6010
rect 20411 5958 20457 6010
rect 20161 5956 20217 5958
rect 20241 5956 20297 5958
rect 20321 5956 20377 5958
rect 20401 5956 20457 5958
rect 16320 5466 16376 5468
rect 16400 5466 16456 5468
rect 16480 5466 16536 5468
rect 16560 5466 16616 5468
rect 16320 5414 16366 5466
rect 16366 5414 16376 5466
rect 16400 5414 16430 5466
rect 16430 5414 16442 5466
rect 16442 5414 16456 5466
rect 16480 5414 16494 5466
rect 16494 5414 16506 5466
rect 16506 5414 16536 5466
rect 16560 5414 16570 5466
rect 16570 5414 16616 5466
rect 16320 5412 16376 5414
rect 16400 5412 16456 5414
rect 16480 5412 16536 5414
rect 16560 5412 16616 5414
rect 24002 5466 24058 5468
rect 24082 5466 24138 5468
rect 24162 5466 24218 5468
rect 24242 5466 24298 5468
rect 24002 5414 24048 5466
rect 24048 5414 24058 5466
rect 24082 5414 24112 5466
rect 24112 5414 24124 5466
rect 24124 5414 24138 5466
rect 24162 5414 24176 5466
rect 24176 5414 24188 5466
rect 24188 5414 24218 5466
rect 24242 5414 24252 5466
rect 24252 5414 24298 5466
rect 24002 5412 24058 5414
rect 24082 5412 24138 5414
rect 24162 5412 24218 5414
rect 24242 5412 24298 5414
rect 5170 5208 5226 5264
rect 25134 10240 25190 10296
rect 25410 16360 25466 16416
rect 25594 15952 25650 16008
rect 25502 14592 25558 14648
rect 25410 13504 25466 13560
rect 25502 13096 25558 13152
rect 25410 12688 25466 12744
rect 25042 9424 25098 9480
rect 25410 9596 25412 9616
rect 25412 9596 25464 9616
rect 25464 9596 25466 9616
rect 25410 9560 25466 9596
rect 25410 9016 25466 9072
rect 25226 8880 25282 8936
rect 25686 13912 25742 13968
rect 25686 13232 25742 13288
rect 26238 20712 26294 20768
rect 26422 21256 26478 21312
rect 26422 20712 26478 20768
rect 26422 20304 26478 20360
rect 26146 20032 26202 20088
rect 26698 23704 26754 23760
rect 26882 23704 26938 23760
rect 26606 22480 26662 22536
rect 26698 20984 26754 21040
rect 27250 23976 27306 24032
rect 27526 25744 27582 25800
rect 27434 25608 27490 25664
rect 28354 26560 28410 26616
rect 27894 26324 27896 26344
rect 27896 26324 27948 26344
rect 27948 26324 27950 26344
rect 27894 26288 27950 26324
rect 28170 25880 28226 25936
rect 27843 25594 27899 25596
rect 27923 25594 27979 25596
rect 28003 25594 28059 25596
rect 28083 25594 28139 25596
rect 27843 25542 27889 25594
rect 27889 25542 27899 25594
rect 27923 25542 27953 25594
rect 27953 25542 27965 25594
rect 27965 25542 27979 25594
rect 28003 25542 28017 25594
rect 28017 25542 28029 25594
rect 28029 25542 28059 25594
rect 28083 25542 28093 25594
rect 28093 25542 28139 25594
rect 27843 25540 27899 25542
rect 27923 25540 27979 25542
rect 28003 25540 28059 25542
rect 28083 25540 28139 25542
rect 27434 25472 27490 25528
rect 27618 25472 27674 25528
rect 27434 24792 27490 24848
rect 28262 25472 28318 25528
rect 27843 24506 27899 24508
rect 27923 24506 27979 24508
rect 28003 24506 28059 24508
rect 28083 24506 28139 24508
rect 27843 24454 27889 24506
rect 27889 24454 27899 24506
rect 27923 24454 27953 24506
rect 27953 24454 27965 24506
rect 27965 24454 27979 24506
rect 28003 24454 28017 24506
rect 28017 24454 28029 24506
rect 28029 24454 28059 24506
rect 28083 24454 28093 24506
rect 28093 24454 28139 24506
rect 27843 24452 27899 24454
rect 27923 24452 27979 24454
rect 28003 24452 28059 24454
rect 28083 24452 28139 24454
rect 28630 27784 28686 27840
rect 28538 26424 28594 26480
rect 27158 23568 27214 23624
rect 27434 23432 27490 23488
rect 27158 22888 27214 22944
rect 26974 22072 27030 22128
rect 26974 21664 27030 21720
rect 26698 20304 26754 20360
rect 26882 20304 26938 20360
rect 26514 18944 26570 19000
rect 26882 19760 26938 19816
rect 25962 18164 25964 18184
rect 25964 18164 26016 18184
rect 26016 18164 26018 18184
rect 25962 18128 26018 18164
rect 26330 18128 26386 18184
rect 26238 17720 26294 17776
rect 26238 17176 26294 17232
rect 26054 15408 26110 15464
rect 25962 15272 26018 15328
rect 26698 18672 26754 18728
rect 26974 19080 27030 19136
rect 26514 18264 26570 18320
rect 26882 18264 26938 18320
rect 26054 14864 26110 14920
rect 26054 14456 26110 14512
rect 25962 13776 26018 13832
rect 25870 12316 25872 12336
rect 25872 12316 25924 12336
rect 25924 12316 25926 12336
rect 25870 12280 25926 12316
rect 26330 14592 26386 14648
rect 26238 13912 26294 13968
rect 26514 16632 26570 16688
rect 26974 18128 27030 18184
rect 26698 17856 26754 17912
rect 26974 17856 27030 17912
rect 26790 17448 26846 17504
rect 26698 16904 26754 16960
rect 26698 16088 26754 16144
rect 26330 13368 26386 13424
rect 26606 13912 26662 13968
rect 26974 17604 27030 17640
rect 26974 17584 26976 17604
rect 26976 17584 27028 17604
rect 27028 17584 27030 17604
rect 26882 17176 26938 17232
rect 26974 16768 27030 16824
rect 26882 16396 26884 16416
rect 26884 16396 26936 16416
rect 26936 16396 26938 16416
rect 26882 16360 26938 16396
rect 26790 15952 26846 16008
rect 26882 15444 26884 15464
rect 26884 15444 26936 15464
rect 26936 15444 26938 15464
rect 26882 15408 26938 15444
rect 27250 22480 27306 22536
rect 27843 23418 27899 23420
rect 27923 23418 27979 23420
rect 28003 23418 28059 23420
rect 28083 23418 28139 23420
rect 27843 23366 27889 23418
rect 27889 23366 27899 23418
rect 27923 23366 27953 23418
rect 27953 23366 27965 23418
rect 27965 23366 27979 23418
rect 28003 23366 28017 23418
rect 28017 23366 28029 23418
rect 28029 23366 28059 23418
rect 28083 23366 28093 23418
rect 28093 23366 28139 23418
rect 27843 23364 27899 23366
rect 27923 23364 27979 23366
rect 28003 23364 28059 23366
rect 28083 23364 28139 23366
rect 27710 23316 27766 23352
rect 27710 23296 27712 23316
rect 27712 23296 27764 23316
rect 27764 23296 27766 23316
rect 27526 22480 27582 22536
rect 28078 22752 28134 22808
rect 27618 22344 27674 22400
rect 28538 23432 28594 23488
rect 28446 23296 28502 23352
rect 28998 29280 29054 29336
rect 28814 29008 28870 29064
rect 28906 28872 28962 28928
rect 28906 28600 28962 28656
rect 30378 33904 30434 33960
rect 29090 27668 29146 27704
rect 29090 27648 29092 27668
rect 29092 27648 29144 27668
rect 29144 27648 29146 27668
rect 28906 27104 28962 27160
rect 28814 26696 28870 26752
rect 28906 26424 28962 26480
rect 29090 26424 29146 26480
rect 28722 26324 28724 26344
rect 28724 26324 28776 26344
rect 28776 26324 28778 26344
rect 28722 26288 28778 26324
rect 29090 26324 29092 26344
rect 29092 26324 29144 26344
rect 29144 26324 29146 26344
rect 29090 26288 29146 26324
rect 29642 31864 29698 31920
rect 29274 28328 29330 28384
rect 29274 27784 29330 27840
rect 29274 27648 29330 27704
rect 29458 28600 29514 28656
rect 29458 27920 29514 27976
rect 29274 26016 29330 26072
rect 29182 25880 29238 25936
rect 29366 25744 29422 25800
rect 29090 24792 29146 24848
rect 28998 24384 29054 24440
rect 28998 24112 29054 24168
rect 28722 23432 28778 23488
rect 28262 22752 28318 22808
rect 28446 22480 28502 22536
rect 27843 22330 27899 22332
rect 27923 22330 27979 22332
rect 28003 22330 28059 22332
rect 28083 22330 28139 22332
rect 27843 22278 27889 22330
rect 27889 22278 27899 22330
rect 27923 22278 27953 22330
rect 27953 22278 27965 22330
rect 27965 22278 27979 22330
rect 28003 22278 28017 22330
rect 28017 22278 28029 22330
rect 28029 22278 28059 22330
rect 28083 22278 28093 22330
rect 28093 22278 28139 22330
rect 27843 22276 27899 22278
rect 27923 22276 27979 22278
rect 28003 22276 28059 22278
rect 28083 22276 28139 22278
rect 27250 20984 27306 21040
rect 27618 21256 27674 21312
rect 27434 20984 27490 21040
rect 28354 22344 28410 22400
rect 28354 22208 28410 22264
rect 27843 21242 27899 21244
rect 27923 21242 27979 21244
rect 28003 21242 28059 21244
rect 28083 21242 28139 21244
rect 27843 21190 27889 21242
rect 27889 21190 27899 21242
rect 27923 21190 27953 21242
rect 27953 21190 27965 21242
rect 27965 21190 27979 21242
rect 28003 21190 28017 21242
rect 28017 21190 28029 21242
rect 28029 21190 28059 21242
rect 28083 21190 28093 21242
rect 28093 21190 28139 21242
rect 27843 21188 27899 21190
rect 27923 21188 27979 21190
rect 28003 21188 28059 21190
rect 28083 21188 28139 21190
rect 27526 20576 27582 20632
rect 26790 14184 26846 14240
rect 24950 7384 25006 7440
rect 26146 11892 26202 11928
rect 26146 11872 26148 11892
rect 26148 11872 26200 11892
rect 26200 11872 26202 11892
rect 4797 4922 4853 4924
rect 4877 4922 4933 4924
rect 4957 4922 5013 4924
rect 5037 4922 5093 4924
rect 4797 4870 4843 4922
rect 4843 4870 4853 4922
rect 4877 4870 4907 4922
rect 4907 4870 4919 4922
rect 4919 4870 4933 4922
rect 4957 4870 4971 4922
rect 4971 4870 4983 4922
rect 4983 4870 5013 4922
rect 5037 4870 5047 4922
rect 5047 4870 5093 4922
rect 4797 4868 4853 4870
rect 4877 4868 4933 4870
rect 4957 4868 5013 4870
rect 5037 4868 5093 4870
rect 12479 4922 12535 4924
rect 12559 4922 12615 4924
rect 12639 4922 12695 4924
rect 12719 4922 12775 4924
rect 12479 4870 12525 4922
rect 12525 4870 12535 4922
rect 12559 4870 12589 4922
rect 12589 4870 12601 4922
rect 12601 4870 12615 4922
rect 12639 4870 12653 4922
rect 12653 4870 12665 4922
rect 12665 4870 12695 4922
rect 12719 4870 12729 4922
rect 12729 4870 12775 4922
rect 12479 4868 12535 4870
rect 12559 4868 12615 4870
rect 12639 4868 12695 4870
rect 12719 4868 12775 4870
rect 20161 4922 20217 4924
rect 20241 4922 20297 4924
rect 20321 4922 20377 4924
rect 20401 4922 20457 4924
rect 20161 4870 20207 4922
rect 20207 4870 20217 4922
rect 20241 4870 20271 4922
rect 20271 4870 20283 4922
rect 20283 4870 20297 4922
rect 20321 4870 20335 4922
rect 20335 4870 20347 4922
rect 20347 4870 20377 4922
rect 20401 4870 20411 4922
rect 20411 4870 20457 4922
rect 20161 4868 20217 4870
rect 20241 4868 20297 4870
rect 20321 4868 20377 4870
rect 20401 4868 20457 4870
rect 26882 13776 26938 13832
rect 26606 11348 26662 11384
rect 26606 11328 26608 11348
rect 26608 11328 26660 11348
rect 26660 11328 26662 11348
rect 26606 10412 26608 10432
rect 26608 10412 26660 10432
rect 26660 10412 26662 10432
rect 26606 10376 26662 10412
rect 26422 9696 26478 9752
rect 26422 9324 26424 9344
rect 26424 9324 26476 9344
rect 26476 9324 26478 9344
rect 26422 9288 26478 9324
rect 27250 20032 27306 20088
rect 27250 19372 27306 19408
rect 27250 19352 27252 19372
rect 27252 19352 27304 19372
rect 27304 19352 27306 19372
rect 27250 18672 27306 18728
rect 26974 11872 27030 11928
rect 27434 20032 27490 20088
rect 27802 20304 27858 20360
rect 27843 20154 27899 20156
rect 27923 20154 27979 20156
rect 28003 20154 28059 20156
rect 28083 20154 28139 20156
rect 27843 20102 27889 20154
rect 27889 20102 27899 20154
rect 27923 20102 27953 20154
rect 27953 20102 27965 20154
rect 27965 20102 27979 20154
rect 28003 20102 28017 20154
rect 28017 20102 28029 20154
rect 28029 20102 28059 20154
rect 28083 20102 28093 20154
rect 28093 20102 28139 20154
rect 27843 20100 27899 20102
rect 27923 20100 27979 20102
rect 28003 20100 28059 20102
rect 28083 20100 28139 20102
rect 27434 18944 27490 19000
rect 27434 18708 27436 18728
rect 27436 18708 27488 18728
rect 27488 18708 27490 18728
rect 27434 18672 27490 18708
rect 27710 19624 27766 19680
rect 27710 19352 27766 19408
rect 28262 21120 28318 21176
rect 28262 20032 28318 20088
rect 28814 23316 28870 23352
rect 28814 23296 28816 23316
rect 28816 23296 28868 23316
rect 28868 23296 28870 23316
rect 28630 23024 28686 23080
rect 28814 23060 28816 23080
rect 28816 23060 28868 23080
rect 28868 23060 28870 23080
rect 28814 23024 28870 23060
rect 29274 24112 29330 24168
rect 29090 23432 29146 23488
rect 29734 31456 29790 31512
rect 30010 30640 30066 30696
rect 29918 29588 29920 29608
rect 29920 29588 29972 29608
rect 29972 29588 29974 29608
rect 29918 29552 29974 29588
rect 29826 29008 29882 29064
rect 29550 27240 29606 27296
rect 29826 28056 29882 28112
rect 29826 27648 29882 27704
rect 29826 27240 29882 27296
rect 29826 26016 29882 26072
rect 29642 25608 29698 25664
rect 29642 25492 29698 25528
rect 29826 25608 29882 25664
rect 29642 25472 29644 25492
rect 29644 25472 29696 25492
rect 29696 25472 29698 25492
rect 29734 25200 29790 25256
rect 30010 28328 30066 28384
rect 29826 24812 29882 24848
rect 29826 24792 29828 24812
rect 29828 24792 29880 24812
rect 29880 24792 29882 24812
rect 30562 32408 30618 32464
rect 31684 32666 31740 32668
rect 31764 32666 31820 32668
rect 31844 32666 31900 32668
rect 31924 32666 31980 32668
rect 31684 32614 31730 32666
rect 31730 32614 31740 32666
rect 31764 32614 31794 32666
rect 31794 32614 31806 32666
rect 31806 32614 31820 32666
rect 31844 32614 31858 32666
rect 31858 32614 31870 32666
rect 31870 32614 31900 32666
rect 31924 32614 31934 32666
rect 31934 32614 31980 32666
rect 31684 32612 31740 32614
rect 31764 32612 31820 32614
rect 31844 32612 31900 32614
rect 31924 32612 31980 32614
rect 30378 28464 30434 28520
rect 30102 27104 30158 27160
rect 30102 26460 30104 26480
rect 30104 26460 30156 26480
rect 30156 26460 30158 26480
rect 30102 26424 30158 26460
rect 29826 24248 29882 24304
rect 28630 21120 28686 21176
rect 28998 21800 29054 21856
rect 28814 21392 28870 21448
rect 28998 21392 29054 21448
rect 28814 20304 28870 20360
rect 28630 20168 28686 20224
rect 28630 19352 28686 19408
rect 27843 19066 27899 19068
rect 27923 19066 27979 19068
rect 28003 19066 28059 19068
rect 28083 19066 28139 19068
rect 27843 19014 27889 19066
rect 27889 19014 27899 19066
rect 27923 19014 27953 19066
rect 27953 19014 27965 19066
rect 27965 19014 27979 19066
rect 28003 19014 28017 19066
rect 28017 19014 28029 19066
rect 28029 19014 28059 19066
rect 28083 19014 28093 19066
rect 28093 19014 28139 19066
rect 27843 19012 27899 19014
rect 27923 19012 27979 19014
rect 28003 19012 28059 19014
rect 28083 19012 28139 19014
rect 27526 18128 27582 18184
rect 27434 17992 27490 18048
rect 27802 18672 27858 18728
rect 28262 19080 28318 19136
rect 28446 18964 28502 19000
rect 28446 18944 28448 18964
rect 28448 18944 28500 18964
rect 28500 18944 28502 18964
rect 28078 18164 28080 18184
rect 28080 18164 28132 18184
rect 28132 18164 28134 18184
rect 28078 18128 28134 18164
rect 27843 17978 27899 17980
rect 27923 17978 27979 17980
rect 28003 17978 28059 17980
rect 28083 17978 28139 17980
rect 27843 17926 27889 17978
rect 27889 17926 27899 17978
rect 27923 17926 27953 17978
rect 27953 17926 27965 17978
rect 27965 17926 27979 17978
rect 28003 17926 28017 17978
rect 28017 17926 28029 17978
rect 28029 17926 28059 17978
rect 28083 17926 28093 17978
rect 28093 17926 28139 17978
rect 27843 17924 27899 17926
rect 27923 17924 27979 17926
rect 28003 17924 28059 17926
rect 28083 17924 28139 17926
rect 27710 17856 27766 17912
rect 28262 17856 28318 17912
rect 27710 17740 27766 17776
rect 27710 17720 27712 17740
rect 27712 17720 27764 17740
rect 27764 17720 27766 17740
rect 27434 17448 27490 17504
rect 28078 17448 28134 17504
rect 28538 18264 28594 18320
rect 28262 17484 28264 17504
rect 28264 17484 28316 17504
rect 28316 17484 28318 17504
rect 28262 17448 28318 17484
rect 27434 16768 27490 16824
rect 27434 16652 27490 16688
rect 27434 16632 27436 16652
rect 27436 16632 27488 16652
rect 27488 16632 27490 16652
rect 27843 16890 27899 16892
rect 27923 16890 27979 16892
rect 28003 16890 28059 16892
rect 28083 16890 28139 16892
rect 27843 16838 27889 16890
rect 27889 16838 27899 16890
rect 27923 16838 27953 16890
rect 27953 16838 27965 16890
rect 27965 16838 27979 16890
rect 28003 16838 28017 16890
rect 28017 16838 28029 16890
rect 28029 16838 28059 16890
rect 28083 16838 28093 16890
rect 28093 16838 28139 16890
rect 27843 16836 27899 16838
rect 27923 16836 27979 16838
rect 28003 16836 28059 16838
rect 28083 16836 28139 16838
rect 28170 16632 28226 16688
rect 28630 18128 28686 18184
rect 28630 17720 28686 17776
rect 28538 17176 28594 17232
rect 28538 16768 28594 16824
rect 28078 16224 28134 16280
rect 27843 15802 27899 15804
rect 27923 15802 27979 15804
rect 28003 15802 28059 15804
rect 28083 15802 28139 15804
rect 27843 15750 27889 15802
rect 27889 15750 27899 15802
rect 27923 15750 27953 15802
rect 27953 15750 27965 15802
rect 27965 15750 27979 15802
rect 28003 15750 28017 15802
rect 28017 15750 28029 15802
rect 28029 15750 28059 15802
rect 28083 15750 28093 15802
rect 28093 15750 28139 15802
rect 27843 15748 27899 15750
rect 27923 15748 27979 15750
rect 28003 15748 28059 15750
rect 28083 15748 28139 15750
rect 28446 16224 28502 16280
rect 27894 15272 27950 15328
rect 27342 12980 27398 13016
rect 27342 12960 27344 12980
rect 27344 12960 27396 12980
rect 27396 12960 27398 12980
rect 27843 14714 27899 14716
rect 27923 14714 27979 14716
rect 28003 14714 28059 14716
rect 28083 14714 28139 14716
rect 27843 14662 27889 14714
rect 27889 14662 27899 14714
rect 27923 14662 27953 14714
rect 27953 14662 27965 14714
rect 27965 14662 27979 14714
rect 28003 14662 28017 14714
rect 28017 14662 28029 14714
rect 28029 14662 28059 14714
rect 28083 14662 28093 14714
rect 28093 14662 28139 14714
rect 27843 14660 27899 14662
rect 27923 14660 27979 14662
rect 28003 14660 28059 14662
rect 28083 14660 28139 14662
rect 28078 14456 28134 14512
rect 28170 13776 28226 13832
rect 27843 13626 27899 13628
rect 27923 13626 27979 13628
rect 28003 13626 28059 13628
rect 28083 13626 28139 13628
rect 27843 13574 27889 13626
rect 27889 13574 27899 13626
rect 27923 13574 27953 13626
rect 27953 13574 27965 13626
rect 27965 13574 27979 13626
rect 28003 13574 28017 13626
rect 28017 13574 28029 13626
rect 28029 13574 28059 13626
rect 28083 13574 28093 13626
rect 28093 13574 28139 13626
rect 27843 13572 27899 13574
rect 27923 13572 27979 13574
rect 28003 13572 28059 13574
rect 28083 13572 28139 13574
rect 27710 12824 27766 12880
rect 27618 12416 27674 12472
rect 27843 12538 27899 12540
rect 27923 12538 27979 12540
rect 28003 12538 28059 12540
rect 28083 12538 28139 12540
rect 27843 12486 27889 12538
rect 27889 12486 27899 12538
rect 27923 12486 27953 12538
rect 27953 12486 27965 12538
rect 27965 12486 27979 12538
rect 28003 12486 28017 12538
rect 28017 12486 28029 12538
rect 28029 12486 28059 12538
rect 28083 12486 28093 12538
rect 28093 12486 28139 12538
rect 27843 12484 27899 12486
rect 27923 12484 27979 12486
rect 28003 12484 28059 12486
rect 28083 12484 28139 12486
rect 27843 11450 27899 11452
rect 27923 11450 27979 11452
rect 28003 11450 28059 11452
rect 28083 11450 28139 11452
rect 27843 11398 27889 11450
rect 27889 11398 27899 11450
rect 27923 11398 27953 11450
rect 27953 11398 27965 11450
rect 27965 11398 27979 11450
rect 28003 11398 28017 11450
rect 28017 11398 28029 11450
rect 28029 11398 28059 11450
rect 28083 11398 28093 11450
rect 28093 11398 28139 11450
rect 27843 11396 27899 11398
rect 27923 11396 27979 11398
rect 28003 11396 28059 11398
rect 28083 11396 28139 11398
rect 28446 14340 28502 14376
rect 28446 14320 28448 14340
rect 28448 14320 28500 14340
rect 28500 14320 28502 14340
rect 28630 15564 28686 15600
rect 28630 15544 28632 15564
rect 28632 15544 28684 15564
rect 28684 15544 28686 15564
rect 28630 15020 28686 15056
rect 28630 15000 28632 15020
rect 28632 15000 28684 15020
rect 28684 15000 28686 15020
rect 28630 14728 28686 14784
rect 28630 14592 28686 14648
rect 28814 19080 28870 19136
rect 28998 21256 29054 21312
rect 29090 20848 29146 20904
rect 28998 20304 29054 20360
rect 28998 19372 29054 19408
rect 28998 19352 29000 19372
rect 29000 19352 29052 19372
rect 29052 19352 29054 19372
rect 29182 19116 29184 19136
rect 29184 19116 29236 19136
rect 29236 19116 29238 19136
rect 29182 19080 29238 19116
rect 29182 18944 29238 19000
rect 29090 18536 29146 18592
rect 28906 17176 28962 17232
rect 28722 13232 28778 13288
rect 28538 12824 28594 12880
rect 27618 10920 27674 10976
rect 27843 10362 27899 10364
rect 27923 10362 27979 10364
rect 28003 10362 28059 10364
rect 28083 10362 28139 10364
rect 27843 10310 27889 10362
rect 27889 10310 27899 10362
rect 27923 10310 27953 10362
rect 27953 10310 27965 10362
rect 27965 10310 27979 10362
rect 28003 10310 28017 10362
rect 28017 10310 28029 10362
rect 28029 10310 28059 10362
rect 28083 10310 28093 10362
rect 28093 10310 28139 10362
rect 27843 10308 27899 10310
rect 27923 10308 27979 10310
rect 28003 10308 28059 10310
rect 28083 10308 28139 10310
rect 27843 9274 27899 9276
rect 27923 9274 27979 9276
rect 28003 9274 28059 9276
rect 28083 9274 28139 9276
rect 27843 9222 27889 9274
rect 27889 9222 27899 9274
rect 27923 9222 27953 9274
rect 27953 9222 27965 9274
rect 27965 9222 27979 9274
rect 28003 9222 28017 9274
rect 28017 9222 28029 9274
rect 28029 9222 28059 9274
rect 28083 9222 28093 9274
rect 28093 9222 28139 9274
rect 27843 9220 27899 9222
rect 27923 9220 27979 9222
rect 28003 9220 28059 9222
rect 28083 9220 28139 9222
rect 27843 8186 27899 8188
rect 27923 8186 27979 8188
rect 28003 8186 28059 8188
rect 28083 8186 28139 8188
rect 27843 8134 27889 8186
rect 27889 8134 27899 8186
rect 27923 8134 27953 8186
rect 27953 8134 27965 8186
rect 27965 8134 27979 8186
rect 28003 8134 28017 8186
rect 28017 8134 28029 8186
rect 28029 8134 28059 8186
rect 28083 8134 28093 8186
rect 28093 8134 28139 8186
rect 27843 8132 27899 8134
rect 27923 8132 27979 8134
rect 28003 8132 28059 8134
rect 28083 8132 28139 8134
rect 27618 7792 27674 7848
rect 27843 7098 27899 7100
rect 27923 7098 27979 7100
rect 28003 7098 28059 7100
rect 28083 7098 28139 7100
rect 27843 7046 27889 7098
rect 27889 7046 27899 7098
rect 27923 7046 27953 7098
rect 27953 7046 27965 7098
rect 27965 7046 27979 7098
rect 28003 7046 28017 7098
rect 28017 7046 28029 7098
rect 28029 7046 28059 7098
rect 28083 7046 28093 7098
rect 28093 7046 28139 7098
rect 27843 7044 27899 7046
rect 27923 7044 27979 7046
rect 28003 7044 28059 7046
rect 28083 7044 28139 7046
rect 27843 6010 27899 6012
rect 27923 6010 27979 6012
rect 28003 6010 28059 6012
rect 28083 6010 28139 6012
rect 27843 5958 27889 6010
rect 27889 5958 27899 6010
rect 27923 5958 27953 6010
rect 27953 5958 27965 6010
rect 27965 5958 27979 6010
rect 28003 5958 28017 6010
rect 28017 5958 28029 6010
rect 28029 5958 28059 6010
rect 28083 5958 28093 6010
rect 28093 5958 28139 6010
rect 27843 5956 27899 5958
rect 27923 5956 27979 5958
rect 28003 5956 28059 5958
rect 28083 5956 28139 5958
rect 28538 11056 28594 11112
rect 28998 16632 29054 16688
rect 29826 23568 29882 23624
rect 29642 22888 29698 22944
rect 29826 23024 29882 23080
rect 29734 22752 29790 22808
rect 29550 21800 29606 21856
rect 29458 20712 29514 20768
rect 29734 21664 29790 21720
rect 30010 23724 30066 23760
rect 30010 23704 30012 23724
rect 30012 23704 30064 23724
rect 30064 23704 30066 23724
rect 30194 23704 30250 23760
rect 30102 23316 30158 23352
rect 30562 30368 30618 30424
rect 30654 28464 30710 28520
rect 30654 27648 30710 27704
rect 30470 27240 30526 27296
rect 30378 25900 30434 25936
rect 30378 25880 30380 25900
rect 30380 25880 30432 25900
rect 30432 25880 30434 25900
rect 30286 23568 30342 23624
rect 30102 23296 30104 23316
rect 30104 23296 30156 23316
rect 30156 23296 30158 23316
rect 30010 22072 30066 22128
rect 29918 21800 29974 21856
rect 29918 21664 29974 21720
rect 29642 20984 29698 21040
rect 29826 21004 29882 21040
rect 29826 20984 29828 21004
rect 29828 20984 29880 21004
rect 29880 20984 29882 21004
rect 30010 20848 30066 20904
rect 29642 20712 29698 20768
rect 29734 20440 29790 20496
rect 29366 18264 29422 18320
rect 29366 17720 29422 17776
rect 29182 17060 29238 17096
rect 29182 17040 29184 17060
rect 29184 17040 29236 17060
rect 29236 17040 29238 17060
rect 29274 16904 29330 16960
rect 28998 16224 29054 16280
rect 29366 16496 29422 16552
rect 29274 16360 29330 16416
rect 29090 15952 29146 16008
rect 29182 15816 29238 15872
rect 29274 15408 29330 15464
rect 29182 15136 29238 15192
rect 28998 14456 29054 14512
rect 29090 14048 29146 14104
rect 29550 16768 29606 16824
rect 29734 18128 29790 18184
rect 29918 20712 29974 20768
rect 29918 20476 29920 20496
rect 29920 20476 29972 20496
rect 29972 20476 29974 20496
rect 29918 20440 29974 20476
rect 30286 21936 30342 21992
rect 30194 20848 30250 20904
rect 30378 20712 30434 20768
rect 30286 20576 30342 20632
rect 31206 31728 31262 31784
rect 31684 31578 31740 31580
rect 31764 31578 31820 31580
rect 31844 31578 31900 31580
rect 31924 31578 31980 31580
rect 31684 31526 31730 31578
rect 31730 31526 31740 31578
rect 31764 31526 31794 31578
rect 31794 31526 31806 31578
rect 31806 31526 31820 31578
rect 31844 31526 31858 31578
rect 31858 31526 31870 31578
rect 31870 31526 31900 31578
rect 31924 31526 31934 31578
rect 31934 31526 31980 31578
rect 31684 31524 31740 31526
rect 31764 31524 31820 31526
rect 31844 31524 31900 31526
rect 31924 31524 31980 31526
rect 30930 30504 30986 30560
rect 31482 30096 31538 30152
rect 31206 29688 31262 29744
rect 30838 26460 30840 26480
rect 30840 26460 30892 26480
rect 30892 26460 30894 26480
rect 30838 26424 30894 26460
rect 30838 26324 30840 26344
rect 30840 26324 30892 26344
rect 30892 26324 30894 26344
rect 30838 26288 30894 26324
rect 31022 26152 31078 26208
rect 30930 25336 30986 25392
rect 30930 25064 30986 25120
rect 30930 24656 30986 24712
rect 30838 24520 30894 24576
rect 30838 23976 30894 24032
rect 31206 27648 31262 27704
rect 31114 24928 31170 24984
rect 31298 25608 31354 25664
rect 31298 25336 31354 25392
rect 31022 23180 31078 23216
rect 31022 23160 31024 23180
rect 31024 23160 31076 23180
rect 31076 23160 31078 23180
rect 30930 22344 30986 22400
rect 30654 21936 30710 21992
rect 29918 19488 29974 19544
rect 30010 19352 30066 19408
rect 29826 17856 29882 17912
rect 29550 16360 29606 16416
rect 29366 14184 29422 14240
rect 28906 13132 28908 13152
rect 28908 13132 28960 13152
rect 28960 13132 28962 13152
rect 28906 13096 28962 13132
rect 28814 11192 28870 11248
rect 29182 13368 29238 13424
rect 29642 15272 29698 15328
rect 29642 13912 29698 13968
rect 30102 18536 30158 18592
rect 30286 19388 30288 19408
rect 30288 19388 30340 19408
rect 30340 19388 30342 19408
rect 30286 19352 30342 19388
rect 30194 18128 30250 18184
rect 30102 17720 30158 17776
rect 29918 15952 29974 16008
rect 30286 17856 30342 17912
rect 30470 20304 30526 20360
rect 30470 19896 30526 19952
rect 30470 19796 30472 19816
rect 30472 19796 30524 19816
rect 30524 19796 30526 19816
rect 30470 19760 30526 19796
rect 30470 18944 30526 19000
rect 30470 18808 30526 18864
rect 30470 17332 30526 17368
rect 30470 17312 30472 17332
rect 30472 17312 30524 17332
rect 30524 17312 30526 17332
rect 30470 17040 30526 17096
rect 30378 16496 30434 16552
rect 30010 15000 30066 15056
rect 29734 13776 29790 13832
rect 28722 6196 28724 6216
rect 28724 6196 28776 6216
rect 28776 6196 28778 6216
rect 28722 6160 28778 6196
rect 29090 8780 29092 8800
rect 29092 8780 29144 8800
rect 29144 8780 29146 8800
rect 29090 8744 29146 8780
rect 29366 6840 29422 6896
rect 30010 13912 30066 13968
rect 30286 14592 30342 14648
rect 29642 10784 29698 10840
rect 29918 10548 29920 10568
rect 29920 10548 29972 10568
rect 29972 10548 29974 10568
rect 29918 10512 29974 10548
rect 29734 9968 29790 10024
rect 30470 15272 30526 15328
rect 30838 21392 30894 21448
rect 30838 21256 30894 21312
rect 30746 20032 30802 20088
rect 31114 21528 31170 21584
rect 31114 21120 31170 21176
rect 31482 24656 31538 24712
rect 31298 22752 31354 22808
rect 31298 22616 31354 22672
rect 31206 20848 31262 20904
rect 31114 19624 31170 19680
rect 31022 19216 31078 19272
rect 31022 18808 31078 18864
rect 30838 18536 30894 18592
rect 30838 18420 30894 18456
rect 30838 18400 30840 18420
rect 30840 18400 30892 18420
rect 30892 18400 30894 18420
rect 30838 18128 30894 18184
rect 30746 17992 30802 18048
rect 30654 17312 30710 17368
rect 30746 17040 30802 17096
rect 30654 16088 30710 16144
rect 30746 15972 30802 16008
rect 30746 15952 30748 15972
rect 30748 15952 30800 15972
rect 30800 15952 30802 15972
rect 30746 15408 30802 15464
rect 30470 14864 30526 14920
rect 30378 14320 30434 14376
rect 29734 8628 29790 8664
rect 29734 8608 29736 8628
rect 29736 8608 29788 8628
rect 29788 8608 29790 8628
rect 30102 8472 30158 8528
rect 30378 8356 30434 8392
rect 30378 8336 30380 8356
rect 30380 8336 30432 8356
rect 30432 8336 30434 8356
rect 29918 7284 29920 7304
rect 29920 7284 29972 7304
rect 29972 7284 29974 7304
rect 29918 7248 29974 7284
rect 30470 6724 30526 6760
rect 30470 6704 30472 6724
rect 30472 6704 30524 6724
rect 30524 6704 30526 6724
rect 28630 5072 28686 5128
rect 27843 4922 27899 4924
rect 27923 4922 27979 4924
rect 28003 4922 28059 4924
rect 28083 4922 28139 4924
rect 27843 4870 27889 4922
rect 27889 4870 27899 4922
rect 27923 4870 27953 4922
rect 27953 4870 27965 4922
rect 27965 4870 27979 4922
rect 28003 4870 28017 4922
rect 28017 4870 28029 4922
rect 28029 4870 28059 4922
rect 28083 4870 28093 4922
rect 28093 4870 28139 4922
rect 27843 4868 27899 4870
rect 27923 4868 27979 4870
rect 28003 4868 28059 4870
rect 28083 4868 28139 4870
rect 8638 4378 8694 4380
rect 8718 4378 8774 4380
rect 8798 4378 8854 4380
rect 8878 4378 8934 4380
rect 8638 4326 8684 4378
rect 8684 4326 8694 4378
rect 8718 4326 8748 4378
rect 8748 4326 8760 4378
rect 8760 4326 8774 4378
rect 8798 4326 8812 4378
rect 8812 4326 8824 4378
rect 8824 4326 8854 4378
rect 8878 4326 8888 4378
rect 8888 4326 8934 4378
rect 8638 4324 8694 4326
rect 8718 4324 8774 4326
rect 8798 4324 8854 4326
rect 8878 4324 8934 4326
rect 16320 4378 16376 4380
rect 16400 4378 16456 4380
rect 16480 4378 16536 4380
rect 16560 4378 16616 4380
rect 16320 4326 16366 4378
rect 16366 4326 16376 4378
rect 16400 4326 16430 4378
rect 16430 4326 16442 4378
rect 16442 4326 16456 4378
rect 16480 4326 16494 4378
rect 16494 4326 16506 4378
rect 16506 4326 16536 4378
rect 16560 4326 16570 4378
rect 16570 4326 16616 4378
rect 16320 4324 16376 4326
rect 16400 4324 16456 4326
rect 16480 4324 16536 4326
rect 16560 4324 16616 4326
rect 24002 4378 24058 4380
rect 24082 4378 24138 4380
rect 24162 4378 24218 4380
rect 24242 4378 24298 4380
rect 24002 4326 24048 4378
rect 24048 4326 24058 4378
rect 24082 4326 24112 4378
rect 24112 4326 24124 4378
rect 24124 4326 24138 4378
rect 24162 4326 24176 4378
rect 24176 4326 24188 4378
rect 24188 4326 24218 4378
rect 24242 4326 24252 4378
rect 24252 4326 24298 4378
rect 24002 4324 24058 4326
rect 24082 4324 24138 4326
rect 24162 4324 24218 4326
rect 24242 4324 24298 4326
rect 1582 4020 1584 4040
rect 1584 4020 1636 4040
rect 1636 4020 1638 4040
rect 1582 3984 1638 4020
rect 31114 13504 31170 13560
rect 31022 10804 31078 10840
rect 31022 10784 31024 10804
rect 31024 10784 31076 10804
rect 31076 10784 31078 10804
rect 30930 10104 30986 10160
rect 31298 20712 31354 20768
rect 31684 30490 31740 30492
rect 31764 30490 31820 30492
rect 31844 30490 31900 30492
rect 31924 30490 31980 30492
rect 31684 30438 31730 30490
rect 31730 30438 31740 30490
rect 31764 30438 31794 30490
rect 31794 30438 31806 30490
rect 31806 30438 31820 30490
rect 31844 30438 31858 30490
rect 31858 30438 31870 30490
rect 31870 30438 31900 30490
rect 31924 30438 31934 30490
rect 31934 30438 31980 30490
rect 31684 30436 31740 30438
rect 31764 30436 31820 30438
rect 31844 30436 31900 30438
rect 31924 30436 31980 30438
rect 31684 29402 31740 29404
rect 31764 29402 31820 29404
rect 31844 29402 31900 29404
rect 31924 29402 31980 29404
rect 31684 29350 31730 29402
rect 31730 29350 31740 29402
rect 31764 29350 31794 29402
rect 31794 29350 31806 29402
rect 31806 29350 31820 29402
rect 31844 29350 31858 29402
rect 31858 29350 31870 29402
rect 31870 29350 31900 29402
rect 31924 29350 31934 29402
rect 31934 29350 31980 29402
rect 31684 29348 31740 29350
rect 31764 29348 31820 29350
rect 31844 29348 31900 29350
rect 31924 29348 31980 29350
rect 31684 28314 31740 28316
rect 31764 28314 31820 28316
rect 31844 28314 31900 28316
rect 31924 28314 31980 28316
rect 31684 28262 31730 28314
rect 31730 28262 31740 28314
rect 31764 28262 31794 28314
rect 31794 28262 31806 28314
rect 31806 28262 31820 28314
rect 31844 28262 31858 28314
rect 31858 28262 31870 28314
rect 31870 28262 31900 28314
rect 31924 28262 31934 28314
rect 31934 28262 31980 28314
rect 31684 28260 31740 28262
rect 31764 28260 31820 28262
rect 31844 28260 31900 28262
rect 31924 28260 31980 28262
rect 31684 27226 31740 27228
rect 31764 27226 31820 27228
rect 31844 27226 31900 27228
rect 31924 27226 31980 27228
rect 31684 27174 31730 27226
rect 31730 27174 31740 27226
rect 31764 27174 31794 27226
rect 31794 27174 31806 27226
rect 31806 27174 31820 27226
rect 31844 27174 31858 27226
rect 31858 27174 31870 27226
rect 31870 27174 31900 27226
rect 31924 27174 31934 27226
rect 31934 27174 31980 27226
rect 31684 27172 31740 27174
rect 31764 27172 31820 27174
rect 31844 27172 31900 27174
rect 31924 27172 31980 27174
rect 31850 26968 31906 27024
rect 32126 26560 32182 26616
rect 32034 26288 32090 26344
rect 31684 26138 31740 26140
rect 31764 26138 31820 26140
rect 31844 26138 31900 26140
rect 31924 26138 31980 26140
rect 31684 26086 31730 26138
rect 31730 26086 31740 26138
rect 31764 26086 31794 26138
rect 31794 26086 31806 26138
rect 31806 26086 31820 26138
rect 31844 26086 31858 26138
rect 31858 26086 31870 26138
rect 31870 26086 31900 26138
rect 31924 26086 31934 26138
rect 31934 26086 31980 26138
rect 31684 26084 31740 26086
rect 31764 26084 31820 26086
rect 31844 26084 31900 26086
rect 31924 26084 31980 26086
rect 31684 25050 31740 25052
rect 31764 25050 31820 25052
rect 31844 25050 31900 25052
rect 31924 25050 31980 25052
rect 31684 24998 31730 25050
rect 31730 24998 31740 25050
rect 31764 24998 31794 25050
rect 31794 24998 31806 25050
rect 31806 24998 31820 25050
rect 31844 24998 31858 25050
rect 31858 24998 31870 25050
rect 31870 24998 31900 25050
rect 31924 24998 31934 25050
rect 31934 24998 31980 25050
rect 31684 24996 31740 24998
rect 31764 24996 31820 24998
rect 31844 24996 31900 24998
rect 31924 24996 31980 24998
rect 32034 24384 32090 24440
rect 31574 24248 31630 24304
rect 31684 23962 31740 23964
rect 31764 23962 31820 23964
rect 31844 23962 31900 23964
rect 31924 23962 31980 23964
rect 31684 23910 31730 23962
rect 31730 23910 31740 23962
rect 31764 23910 31794 23962
rect 31794 23910 31806 23962
rect 31806 23910 31820 23962
rect 31844 23910 31858 23962
rect 31858 23910 31870 23962
rect 31870 23910 31900 23962
rect 31924 23910 31934 23962
rect 31934 23910 31980 23962
rect 31684 23908 31740 23910
rect 31764 23908 31820 23910
rect 31844 23908 31900 23910
rect 31924 23908 31980 23910
rect 31684 22874 31740 22876
rect 31764 22874 31820 22876
rect 31844 22874 31900 22876
rect 31924 22874 31980 22876
rect 31684 22822 31730 22874
rect 31730 22822 31740 22874
rect 31764 22822 31794 22874
rect 31794 22822 31806 22874
rect 31806 22822 31820 22874
rect 31844 22822 31858 22874
rect 31858 22822 31870 22874
rect 31870 22822 31900 22874
rect 31924 22822 31934 22874
rect 31934 22822 31980 22874
rect 31684 22820 31740 22822
rect 31764 22820 31820 22822
rect 31844 22820 31900 22822
rect 31924 22820 31980 22822
rect 31684 21786 31740 21788
rect 31764 21786 31820 21788
rect 31844 21786 31900 21788
rect 31924 21786 31980 21788
rect 31684 21734 31730 21786
rect 31730 21734 31740 21786
rect 31764 21734 31794 21786
rect 31794 21734 31806 21786
rect 31806 21734 31820 21786
rect 31844 21734 31858 21786
rect 31858 21734 31870 21786
rect 31870 21734 31900 21786
rect 31924 21734 31934 21786
rect 31934 21734 31980 21786
rect 31684 21732 31740 21734
rect 31764 21732 31820 21734
rect 31844 21732 31900 21734
rect 31924 21732 31980 21734
rect 31684 20698 31740 20700
rect 31764 20698 31820 20700
rect 31844 20698 31900 20700
rect 31924 20698 31980 20700
rect 31684 20646 31730 20698
rect 31730 20646 31740 20698
rect 31764 20646 31794 20698
rect 31794 20646 31806 20698
rect 31806 20646 31820 20698
rect 31844 20646 31858 20698
rect 31858 20646 31870 20698
rect 31870 20646 31900 20698
rect 31924 20646 31934 20698
rect 31934 20646 31980 20698
rect 31684 20644 31740 20646
rect 31764 20644 31820 20646
rect 31844 20644 31900 20646
rect 31924 20644 31980 20646
rect 31482 20168 31538 20224
rect 31390 19760 31446 19816
rect 31390 19352 31446 19408
rect 31298 16632 31354 16688
rect 31298 16088 31354 16144
rect 31684 19610 31740 19612
rect 31764 19610 31820 19612
rect 31844 19610 31900 19612
rect 31924 19610 31980 19612
rect 31684 19558 31730 19610
rect 31730 19558 31740 19610
rect 31764 19558 31794 19610
rect 31794 19558 31806 19610
rect 31806 19558 31820 19610
rect 31844 19558 31858 19610
rect 31858 19558 31870 19610
rect 31870 19558 31900 19610
rect 31924 19558 31934 19610
rect 31934 19558 31980 19610
rect 31684 19556 31740 19558
rect 31764 19556 31820 19558
rect 31844 19556 31900 19558
rect 31924 19556 31980 19558
rect 31666 18708 31668 18728
rect 31668 18708 31720 18728
rect 31720 18708 31722 18728
rect 31666 18672 31722 18708
rect 31684 18522 31740 18524
rect 31764 18522 31820 18524
rect 31844 18522 31900 18524
rect 31924 18522 31980 18524
rect 31684 18470 31730 18522
rect 31730 18470 31740 18522
rect 31764 18470 31794 18522
rect 31794 18470 31806 18522
rect 31806 18470 31820 18522
rect 31844 18470 31858 18522
rect 31858 18470 31870 18522
rect 31870 18470 31900 18522
rect 31924 18470 31934 18522
rect 31934 18470 31980 18522
rect 31684 18468 31740 18470
rect 31764 18468 31820 18470
rect 31844 18468 31900 18470
rect 31924 18468 31980 18470
rect 32034 17584 32090 17640
rect 31684 17434 31740 17436
rect 31764 17434 31820 17436
rect 31844 17434 31900 17436
rect 31924 17434 31980 17436
rect 31684 17382 31730 17434
rect 31730 17382 31740 17434
rect 31764 17382 31794 17434
rect 31794 17382 31806 17434
rect 31806 17382 31820 17434
rect 31844 17382 31858 17434
rect 31858 17382 31870 17434
rect 31870 17382 31900 17434
rect 31924 17382 31934 17434
rect 31934 17382 31980 17434
rect 31684 17380 31740 17382
rect 31764 17380 31820 17382
rect 31844 17380 31900 17382
rect 31924 17380 31980 17382
rect 32586 30096 32642 30152
rect 32494 25880 32550 25936
rect 32494 25336 32550 25392
rect 32678 29280 32734 29336
rect 32770 26696 32826 26752
rect 32402 23296 32458 23352
rect 31390 13368 31446 13424
rect 31666 17040 31722 17096
rect 32034 16904 32090 16960
rect 31684 16346 31740 16348
rect 31764 16346 31820 16348
rect 31844 16346 31900 16348
rect 31924 16346 31980 16348
rect 31684 16294 31730 16346
rect 31730 16294 31740 16346
rect 31764 16294 31794 16346
rect 31794 16294 31806 16346
rect 31806 16294 31820 16346
rect 31844 16294 31858 16346
rect 31858 16294 31870 16346
rect 31870 16294 31900 16346
rect 31924 16294 31934 16346
rect 31934 16294 31980 16346
rect 31684 16292 31740 16294
rect 31764 16292 31820 16294
rect 31844 16292 31900 16294
rect 31924 16292 31980 16294
rect 31684 15258 31740 15260
rect 31764 15258 31820 15260
rect 31844 15258 31900 15260
rect 31924 15258 31980 15260
rect 31684 15206 31730 15258
rect 31730 15206 31740 15258
rect 31764 15206 31794 15258
rect 31794 15206 31806 15258
rect 31806 15206 31820 15258
rect 31844 15206 31858 15258
rect 31858 15206 31870 15258
rect 31870 15206 31900 15258
rect 31924 15206 31934 15258
rect 31934 15206 31980 15258
rect 31684 15204 31740 15206
rect 31764 15204 31820 15206
rect 31844 15204 31900 15206
rect 31924 15204 31980 15206
rect 31684 14170 31740 14172
rect 31764 14170 31820 14172
rect 31844 14170 31900 14172
rect 31924 14170 31980 14172
rect 31684 14118 31730 14170
rect 31730 14118 31740 14170
rect 31764 14118 31794 14170
rect 31794 14118 31806 14170
rect 31806 14118 31820 14170
rect 31844 14118 31858 14170
rect 31858 14118 31870 14170
rect 31870 14118 31900 14170
rect 31924 14118 31934 14170
rect 31934 14118 31980 14170
rect 31684 14116 31740 14118
rect 31764 14116 31820 14118
rect 31844 14116 31900 14118
rect 31924 14116 31980 14118
rect 31684 13082 31740 13084
rect 31764 13082 31820 13084
rect 31844 13082 31900 13084
rect 31924 13082 31980 13084
rect 31684 13030 31730 13082
rect 31730 13030 31740 13082
rect 31764 13030 31794 13082
rect 31794 13030 31806 13082
rect 31806 13030 31820 13082
rect 31844 13030 31858 13082
rect 31858 13030 31870 13082
rect 31870 13030 31900 13082
rect 31924 13030 31934 13082
rect 31934 13030 31980 13082
rect 31684 13028 31740 13030
rect 31764 13028 31820 13030
rect 31844 13028 31900 13030
rect 31924 13028 31980 13030
rect 31574 12144 31630 12200
rect 31684 11994 31740 11996
rect 31764 11994 31820 11996
rect 31844 11994 31900 11996
rect 31924 11994 31980 11996
rect 31684 11942 31730 11994
rect 31730 11942 31740 11994
rect 31764 11942 31794 11994
rect 31794 11942 31806 11994
rect 31806 11942 31820 11994
rect 31844 11942 31858 11994
rect 31858 11942 31870 11994
rect 31870 11942 31900 11994
rect 31924 11942 31934 11994
rect 31934 11942 31980 11994
rect 31684 11940 31740 11942
rect 31764 11940 31820 11942
rect 31844 11940 31900 11942
rect 31924 11940 31980 11942
rect 31298 11756 31354 11792
rect 31298 11736 31300 11756
rect 31300 11736 31352 11756
rect 31352 11736 31354 11756
rect 31298 11348 31354 11384
rect 31298 11328 31300 11348
rect 31300 11328 31352 11348
rect 31352 11328 31354 11348
rect 31390 10920 31446 10976
rect 31684 10906 31740 10908
rect 31764 10906 31820 10908
rect 31844 10906 31900 10908
rect 31924 10906 31980 10908
rect 31684 10854 31730 10906
rect 31730 10854 31740 10906
rect 31764 10854 31794 10906
rect 31794 10854 31806 10906
rect 31806 10854 31820 10906
rect 31844 10854 31858 10906
rect 31858 10854 31870 10906
rect 31870 10854 31900 10906
rect 31924 10854 31934 10906
rect 31934 10854 31980 10906
rect 31684 10852 31740 10854
rect 31764 10852 31820 10854
rect 31844 10852 31900 10854
rect 31924 10852 31980 10854
rect 31298 10004 31300 10024
rect 31300 10004 31352 10024
rect 31352 10004 31354 10024
rect 31298 9968 31354 10004
rect 31298 9324 31300 9344
rect 31300 9324 31352 9344
rect 31352 9324 31354 9344
rect 31298 9288 31354 9324
rect 31684 9818 31740 9820
rect 31764 9818 31820 9820
rect 31844 9818 31900 9820
rect 31924 9818 31980 9820
rect 31684 9766 31730 9818
rect 31730 9766 31740 9818
rect 31764 9766 31794 9818
rect 31794 9766 31806 9818
rect 31806 9766 31820 9818
rect 31844 9766 31858 9818
rect 31858 9766 31870 9818
rect 31870 9766 31900 9818
rect 31924 9766 31934 9818
rect 31934 9766 31980 9818
rect 31684 9764 31740 9766
rect 31764 9764 31820 9766
rect 31844 9764 31900 9766
rect 31924 9764 31980 9766
rect 31684 8730 31740 8732
rect 31764 8730 31820 8732
rect 31844 8730 31900 8732
rect 31924 8730 31980 8732
rect 31684 8678 31730 8730
rect 31730 8678 31740 8730
rect 31764 8678 31794 8730
rect 31794 8678 31806 8730
rect 31806 8678 31820 8730
rect 31844 8678 31858 8730
rect 31858 8678 31870 8730
rect 31870 8678 31900 8730
rect 31924 8678 31934 8730
rect 31934 8678 31980 8730
rect 31684 8676 31740 8678
rect 31764 8676 31820 8678
rect 31844 8676 31900 8678
rect 31924 8676 31980 8678
rect 32126 15680 32182 15736
rect 31298 7928 31354 7984
rect 31684 7642 31740 7644
rect 31764 7642 31820 7644
rect 31844 7642 31900 7644
rect 31924 7642 31980 7644
rect 31684 7590 31730 7642
rect 31730 7590 31740 7642
rect 31764 7590 31794 7642
rect 31794 7590 31806 7642
rect 31806 7590 31820 7642
rect 31844 7590 31858 7642
rect 31858 7590 31870 7642
rect 31870 7590 31900 7642
rect 31924 7590 31934 7642
rect 31934 7590 31980 7642
rect 31684 7588 31740 7590
rect 31764 7588 31820 7590
rect 31844 7588 31900 7590
rect 31924 7588 31980 7590
rect 32218 14320 32274 14376
rect 32678 15816 32734 15872
rect 31298 7268 31354 7304
rect 31298 7248 31300 7268
rect 31300 7248 31352 7268
rect 31352 7248 31354 7268
rect 31684 6554 31740 6556
rect 31764 6554 31820 6556
rect 31844 6554 31900 6556
rect 31924 6554 31980 6556
rect 31684 6502 31730 6554
rect 31730 6502 31740 6554
rect 31764 6502 31794 6554
rect 31794 6502 31806 6554
rect 31806 6502 31820 6554
rect 31844 6502 31858 6554
rect 31858 6502 31870 6554
rect 31870 6502 31900 6554
rect 31924 6502 31934 6554
rect 31934 6502 31980 6554
rect 31684 6500 31740 6502
rect 31764 6500 31820 6502
rect 31844 6500 31900 6502
rect 31924 6500 31980 6502
rect 31298 5888 31354 5944
rect 31684 5466 31740 5468
rect 31764 5466 31820 5468
rect 31844 5466 31900 5468
rect 31924 5466 31980 5468
rect 31684 5414 31730 5466
rect 31730 5414 31740 5466
rect 31764 5414 31794 5466
rect 31794 5414 31806 5466
rect 31806 5414 31820 5466
rect 31844 5414 31858 5466
rect 31858 5414 31870 5466
rect 31870 5414 31900 5466
rect 31924 5414 31934 5466
rect 31934 5414 31980 5466
rect 31684 5412 31740 5414
rect 31764 5412 31820 5414
rect 31844 5412 31900 5414
rect 31924 5412 31980 5414
rect 31298 5208 31354 5264
rect 31684 4378 31740 4380
rect 31764 4378 31820 4380
rect 31844 4378 31900 4380
rect 31924 4378 31980 4380
rect 31684 4326 31730 4378
rect 31730 4326 31740 4378
rect 31764 4326 31794 4378
rect 31794 4326 31806 4378
rect 31806 4326 31820 4378
rect 31844 4326 31858 4378
rect 31858 4326 31870 4378
rect 31870 4326 31900 4378
rect 31924 4326 31934 4378
rect 31934 4326 31980 4378
rect 31684 4324 31740 4326
rect 31764 4324 31820 4326
rect 31844 4324 31900 4326
rect 31924 4324 31980 4326
rect 31298 3884 31300 3904
rect 31300 3884 31352 3904
rect 31352 3884 31354 3904
rect 4797 3834 4853 3836
rect 4877 3834 4933 3836
rect 4957 3834 5013 3836
rect 5037 3834 5093 3836
rect 4797 3782 4843 3834
rect 4843 3782 4853 3834
rect 4877 3782 4907 3834
rect 4907 3782 4919 3834
rect 4919 3782 4933 3834
rect 4957 3782 4971 3834
rect 4971 3782 4983 3834
rect 4983 3782 5013 3834
rect 5037 3782 5047 3834
rect 5047 3782 5093 3834
rect 4797 3780 4853 3782
rect 4877 3780 4933 3782
rect 4957 3780 5013 3782
rect 5037 3780 5093 3782
rect 12479 3834 12535 3836
rect 12559 3834 12615 3836
rect 12639 3834 12695 3836
rect 12719 3834 12775 3836
rect 12479 3782 12525 3834
rect 12525 3782 12535 3834
rect 12559 3782 12589 3834
rect 12589 3782 12601 3834
rect 12601 3782 12615 3834
rect 12639 3782 12653 3834
rect 12653 3782 12665 3834
rect 12665 3782 12695 3834
rect 12719 3782 12729 3834
rect 12729 3782 12775 3834
rect 12479 3780 12535 3782
rect 12559 3780 12615 3782
rect 12639 3780 12695 3782
rect 12719 3780 12775 3782
rect 20161 3834 20217 3836
rect 20241 3834 20297 3836
rect 20321 3834 20377 3836
rect 20401 3834 20457 3836
rect 20161 3782 20207 3834
rect 20207 3782 20217 3834
rect 20241 3782 20271 3834
rect 20271 3782 20283 3834
rect 20283 3782 20297 3834
rect 20321 3782 20335 3834
rect 20335 3782 20347 3834
rect 20347 3782 20377 3834
rect 20401 3782 20411 3834
rect 20411 3782 20457 3834
rect 20161 3780 20217 3782
rect 20241 3780 20297 3782
rect 20321 3780 20377 3782
rect 20401 3780 20457 3782
rect 27843 3834 27899 3836
rect 27923 3834 27979 3836
rect 28003 3834 28059 3836
rect 28083 3834 28139 3836
rect 27843 3782 27889 3834
rect 27889 3782 27899 3834
rect 27923 3782 27953 3834
rect 27953 3782 27965 3834
rect 27965 3782 27979 3834
rect 28003 3782 28017 3834
rect 28017 3782 28029 3834
rect 28029 3782 28059 3834
rect 28083 3782 28093 3834
rect 28093 3782 28139 3834
rect 27843 3780 27899 3782
rect 27923 3780 27979 3782
rect 28003 3780 28059 3782
rect 28083 3780 28139 3782
rect 31298 3848 31354 3884
rect 31298 3476 31300 3496
rect 31300 3476 31352 3496
rect 31352 3476 31354 3496
rect 31298 3440 31354 3476
rect 8638 3290 8694 3292
rect 8718 3290 8774 3292
rect 8798 3290 8854 3292
rect 8878 3290 8934 3292
rect 8638 3238 8684 3290
rect 8684 3238 8694 3290
rect 8718 3238 8748 3290
rect 8748 3238 8760 3290
rect 8760 3238 8774 3290
rect 8798 3238 8812 3290
rect 8812 3238 8824 3290
rect 8824 3238 8854 3290
rect 8878 3238 8888 3290
rect 8888 3238 8934 3290
rect 8638 3236 8694 3238
rect 8718 3236 8774 3238
rect 8798 3236 8854 3238
rect 8878 3236 8934 3238
rect 16320 3290 16376 3292
rect 16400 3290 16456 3292
rect 16480 3290 16536 3292
rect 16560 3290 16616 3292
rect 16320 3238 16366 3290
rect 16366 3238 16376 3290
rect 16400 3238 16430 3290
rect 16430 3238 16442 3290
rect 16442 3238 16456 3290
rect 16480 3238 16494 3290
rect 16494 3238 16506 3290
rect 16506 3238 16536 3290
rect 16560 3238 16570 3290
rect 16570 3238 16616 3290
rect 16320 3236 16376 3238
rect 16400 3236 16456 3238
rect 16480 3236 16536 3238
rect 16560 3236 16616 3238
rect 24002 3290 24058 3292
rect 24082 3290 24138 3292
rect 24162 3290 24218 3292
rect 24242 3290 24298 3292
rect 24002 3238 24048 3290
rect 24048 3238 24058 3290
rect 24082 3238 24112 3290
rect 24112 3238 24124 3290
rect 24124 3238 24138 3290
rect 24162 3238 24176 3290
rect 24176 3238 24188 3290
rect 24188 3238 24218 3290
rect 24242 3238 24252 3290
rect 24252 3238 24298 3290
rect 24002 3236 24058 3238
rect 24082 3236 24138 3238
rect 24162 3236 24218 3238
rect 24242 3236 24298 3238
rect 31684 3290 31740 3292
rect 31764 3290 31820 3292
rect 31844 3290 31900 3292
rect 31924 3290 31980 3292
rect 31684 3238 31730 3290
rect 31730 3238 31740 3290
rect 31764 3238 31794 3290
rect 31794 3238 31806 3290
rect 31806 3238 31820 3290
rect 31844 3238 31858 3290
rect 31858 3238 31870 3290
rect 31870 3238 31900 3290
rect 31924 3238 31934 3290
rect 31934 3238 31980 3290
rect 31684 3236 31740 3238
rect 31764 3236 31820 3238
rect 31844 3236 31900 3238
rect 31924 3236 31980 3238
rect 1582 3168 1638 3224
rect 4797 2746 4853 2748
rect 4877 2746 4933 2748
rect 4957 2746 5013 2748
rect 5037 2746 5093 2748
rect 4797 2694 4843 2746
rect 4843 2694 4853 2746
rect 4877 2694 4907 2746
rect 4907 2694 4919 2746
rect 4919 2694 4933 2746
rect 4957 2694 4971 2746
rect 4971 2694 4983 2746
rect 4983 2694 5013 2746
rect 5037 2694 5047 2746
rect 5047 2694 5093 2746
rect 4797 2692 4853 2694
rect 4877 2692 4933 2694
rect 4957 2692 5013 2694
rect 5037 2692 5093 2694
rect 12479 2746 12535 2748
rect 12559 2746 12615 2748
rect 12639 2746 12695 2748
rect 12719 2746 12775 2748
rect 12479 2694 12525 2746
rect 12525 2694 12535 2746
rect 12559 2694 12589 2746
rect 12589 2694 12601 2746
rect 12601 2694 12615 2746
rect 12639 2694 12653 2746
rect 12653 2694 12665 2746
rect 12665 2694 12695 2746
rect 12719 2694 12729 2746
rect 12729 2694 12775 2746
rect 12479 2692 12535 2694
rect 12559 2692 12615 2694
rect 12639 2692 12695 2694
rect 12719 2692 12775 2694
rect 20161 2746 20217 2748
rect 20241 2746 20297 2748
rect 20321 2746 20377 2748
rect 20401 2746 20457 2748
rect 20161 2694 20207 2746
rect 20207 2694 20217 2746
rect 20241 2694 20271 2746
rect 20271 2694 20283 2746
rect 20283 2694 20297 2746
rect 20321 2694 20335 2746
rect 20335 2694 20347 2746
rect 20347 2694 20377 2746
rect 20401 2694 20411 2746
rect 20411 2694 20457 2746
rect 20161 2692 20217 2694
rect 20241 2692 20297 2694
rect 20321 2692 20377 2694
rect 20401 2692 20457 2694
rect 27843 2746 27899 2748
rect 27923 2746 27979 2748
rect 28003 2746 28059 2748
rect 28083 2746 28139 2748
rect 27843 2694 27889 2746
rect 27889 2694 27899 2746
rect 27923 2694 27953 2746
rect 27953 2694 27965 2746
rect 27965 2694 27979 2746
rect 28003 2694 28017 2746
rect 28017 2694 28029 2746
rect 28029 2694 28059 2746
rect 28083 2694 28093 2746
rect 28093 2694 28139 2746
rect 27843 2692 27899 2694
rect 27923 2692 27979 2694
rect 28003 2692 28059 2694
rect 28083 2692 28139 2694
rect 8638 2202 8694 2204
rect 8718 2202 8774 2204
rect 8798 2202 8854 2204
rect 8878 2202 8934 2204
rect 8638 2150 8684 2202
rect 8684 2150 8694 2202
rect 8718 2150 8748 2202
rect 8748 2150 8760 2202
rect 8760 2150 8774 2202
rect 8798 2150 8812 2202
rect 8812 2150 8824 2202
rect 8824 2150 8854 2202
rect 8878 2150 8888 2202
rect 8888 2150 8934 2202
rect 8638 2148 8694 2150
rect 8718 2148 8774 2150
rect 8798 2148 8854 2150
rect 8878 2148 8934 2150
rect 16320 2202 16376 2204
rect 16400 2202 16456 2204
rect 16480 2202 16536 2204
rect 16560 2202 16616 2204
rect 16320 2150 16366 2202
rect 16366 2150 16376 2202
rect 16400 2150 16430 2202
rect 16430 2150 16442 2202
rect 16442 2150 16456 2202
rect 16480 2150 16494 2202
rect 16494 2150 16506 2202
rect 16506 2150 16536 2202
rect 16560 2150 16570 2202
rect 16570 2150 16616 2202
rect 16320 2148 16376 2150
rect 16400 2148 16456 2150
rect 16480 2148 16536 2150
rect 16560 2148 16616 2150
rect 24002 2202 24058 2204
rect 24082 2202 24138 2204
rect 24162 2202 24218 2204
rect 24242 2202 24298 2204
rect 24002 2150 24048 2202
rect 24048 2150 24058 2202
rect 24082 2150 24112 2202
rect 24112 2150 24124 2202
rect 24124 2150 24138 2202
rect 24162 2150 24176 2202
rect 24176 2150 24188 2202
rect 24188 2150 24218 2202
rect 24242 2150 24252 2202
rect 24252 2150 24298 2202
rect 24002 2148 24058 2150
rect 24082 2148 24138 2150
rect 24162 2148 24218 2150
rect 24242 2148 24298 2150
rect 31684 2202 31740 2204
rect 31764 2202 31820 2204
rect 31844 2202 31900 2204
rect 31924 2202 31980 2204
rect 31684 2150 31730 2202
rect 31730 2150 31740 2202
rect 31764 2150 31794 2202
rect 31794 2150 31806 2202
rect 31806 2150 31820 2202
rect 31844 2150 31858 2202
rect 31858 2150 31870 2202
rect 31870 2150 31900 2202
rect 31924 2150 31934 2202
rect 31934 2150 31980 2202
rect 31684 2148 31740 2150
rect 31764 2148 31820 2150
rect 31844 2148 31900 2150
rect 31924 2148 31980 2150
rect 1582 1536 1638 1592
rect 1398 720 1454 776
<< metal3 >>
rect 6637 34914 6703 34917
rect 22134 34914 22140 34916
rect 6637 34912 22140 34914
rect 6637 34856 6642 34912
rect 6698 34856 22140 34912
rect 6637 34854 22140 34856
rect 6637 34851 6703 34854
rect 22134 34852 22140 34854
rect 22204 34852 22210 34916
rect 3969 34778 4035 34781
rect 20846 34778 20852 34780
rect 3969 34776 20852 34778
rect 3969 34720 3974 34776
rect 4030 34720 20852 34776
rect 3969 34718 20852 34720
rect 3969 34715 4035 34718
rect 20846 34716 20852 34718
rect 20916 34716 20922 34780
rect 10174 34580 10180 34644
rect 10244 34642 10250 34644
rect 25313 34642 25379 34645
rect 10244 34640 25379 34642
rect 10244 34584 25318 34640
rect 25374 34584 25379 34640
rect 10244 34582 25379 34584
rect 10244 34580 10250 34582
rect 25313 34579 25379 34582
rect 14825 34506 14891 34509
rect 24945 34506 25011 34509
rect 14825 34504 25011 34506
rect 14825 34448 14830 34504
rect 14886 34448 24950 34504
rect 25006 34448 25011 34504
rect 14825 34446 25011 34448
rect 14825 34443 14891 34446
rect 24945 34443 25011 34446
rect 17309 34370 17375 34373
rect 29085 34370 29151 34373
rect 17309 34368 29151 34370
rect 17309 34312 17314 34368
rect 17370 34312 29090 34368
rect 29146 34312 29151 34368
rect 17309 34310 29151 34312
rect 17309 34307 17375 34310
rect 29085 34307 29151 34310
rect 0 34144 800 34264
rect 13261 34234 13327 34237
rect 26550 34234 26556 34236
rect 13261 34232 26556 34234
rect 13261 34176 13266 34232
rect 13322 34176 26556 34232
rect 13261 34174 26556 34176
rect 13261 34171 13327 34174
rect 26550 34172 26556 34174
rect 26620 34172 26626 34236
rect 9254 34036 9260 34100
rect 9324 34098 9330 34100
rect 26785 34098 26851 34101
rect 9324 34096 26851 34098
rect 9324 34040 26790 34096
rect 26846 34040 26851 34096
rect 9324 34038 26851 34040
rect 9324 34036 9330 34038
rect 26785 34035 26851 34038
rect 12065 33962 12131 33965
rect 30373 33962 30439 33965
rect 12065 33960 30439 33962
rect 12065 33904 12070 33960
rect 12126 33904 30378 33960
rect 30434 33904 30439 33960
rect 12065 33902 30439 33904
rect 12065 33899 12131 33902
rect 30373 33899 30439 33902
rect 12198 33764 12204 33828
rect 12268 33826 12274 33828
rect 23790 33826 23796 33828
rect 12268 33766 23796 33826
rect 12268 33764 12274 33766
rect 23790 33764 23796 33766
rect 23860 33764 23866 33828
rect 0 33418 800 33448
rect 2865 33418 2931 33421
rect 0 33416 2931 33418
rect 0 33360 2870 33416
rect 2926 33360 2931 33416
rect 0 33358 2931 33360
rect 0 33328 800 33358
rect 2865 33355 2931 33358
rect 15142 33356 15148 33420
rect 15212 33418 15218 33420
rect 30230 33418 30236 33420
rect 15212 33358 30236 33418
rect 15212 33356 15218 33358
rect 30230 33356 30236 33358
rect 30300 33356 30306 33420
rect 16062 33220 16068 33284
rect 16132 33282 16138 33284
rect 25129 33282 25195 33285
rect 16132 33280 25195 33282
rect 16132 33224 25134 33280
rect 25190 33224 25195 33280
rect 16132 33222 25195 33224
rect 16132 33220 16138 33222
rect 25129 33219 25195 33222
rect 6310 33084 6316 33148
rect 6380 33146 6386 33148
rect 19517 33146 19583 33149
rect 6380 33144 19583 33146
rect 6380 33088 19522 33144
rect 19578 33088 19583 33144
rect 6380 33086 19583 33088
rect 6380 33084 6386 33086
rect 19517 33083 19583 33086
rect 19241 32874 19307 32877
rect 30046 32874 30052 32876
rect 19241 32872 30052 32874
rect 19241 32816 19246 32872
rect 19302 32816 30052 32872
rect 19241 32814 30052 32816
rect 19241 32811 19307 32814
rect 30046 32812 30052 32814
rect 30116 32812 30122 32876
rect 19926 32676 19932 32740
rect 19996 32738 20002 32740
rect 23565 32738 23631 32741
rect 19996 32736 23631 32738
rect 19996 32680 23570 32736
rect 23626 32680 23631 32736
rect 19996 32678 23631 32680
rect 19996 32676 20002 32678
rect 23565 32675 23631 32678
rect 8628 32672 8944 32673
rect 0 32602 800 32632
rect 8628 32608 8634 32672
rect 8698 32608 8714 32672
rect 8778 32608 8794 32672
rect 8858 32608 8874 32672
rect 8938 32608 8944 32672
rect 8628 32607 8944 32608
rect 16310 32672 16626 32673
rect 16310 32608 16316 32672
rect 16380 32608 16396 32672
rect 16460 32608 16476 32672
rect 16540 32608 16556 32672
rect 16620 32608 16626 32672
rect 16310 32607 16626 32608
rect 23992 32672 24308 32673
rect 23992 32608 23998 32672
rect 24062 32608 24078 32672
rect 24142 32608 24158 32672
rect 24222 32608 24238 32672
rect 24302 32608 24308 32672
rect 23992 32607 24308 32608
rect 31674 32672 31990 32673
rect 31674 32608 31680 32672
rect 31744 32608 31760 32672
rect 31824 32608 31840 32672
rect 31904 32608 31920 32672
rect 31984 32608 31990 32672
rect 31674 32607 31990 32608
rect 1577 32602 1643 32605
rect 22318 32602 22324 32604
rect 0 32600 1643 32602
rect 0 32544 1582 32600
rect 1638 32544 1643 32600
rect 0 32542 1643 32544
rect 0 32512 800 32542
rect 1577 32539 1643 32542
rect 17910 32542 22324 32602
rect 4337 32466 4403 32469
rect 17910 32466 17970 32542
rect 22318 32540 22324 32542
rect 22388 32540 22394 32604
rect 4337 32464 17970 32466
rect 4337 32408 4342 32464
rect 4398 32408 17970 32464
rect 4337 32406 17970 32408
rect 18045 32466 18111 32469
rect 20662 32466 20668 32468
rect 18045 32464 20668 32466
rect 18045 32408 18050 32464
rect 18106 32408 20668 32464
rect 18045 32406 20668 32408
rect 4337 32403 4403 32406
rect 18045 32403 18111 32406
rect 20662 32404 20668 32406
rect 20732 32404 20738 32468
rect 21357 32466 21423 32469
rect 27061 32466 27127 32469
rect 21357 32464 27127 32466
rect 21357 32408 21362 32464
rect 21418 32408 27066 32464
rect 27122 32408 27127 32464
rect 21357 32406 27127 32408
rect 21357 32403 21423 32406
rect 27061 32403 27127 32406
rect 30557 32466 30623 32469
rect 32206 32466 33006 32496
rect 30557 32464 33006 32466
rect 30557 32408 30562 32464
rect 30618 32408 33006 32464
rect 30557 32406 33006 32408
rect 30557 32403 30623 32406
rect 32206 32376 33006 32406
rect 14365 32330 14431 32333
rect 28349 32330 28415 32333
rect 14365 32328 28415 32330
rect 14365 32272 14370 32328
rect 14426 32272 28354 32328
rect 28410 32272 28415 32328
rect 14365 32270 28415 32272
rect 14365 32267 14431 32270
rect 28349 32267 28415 32270
rect 23749 32194 23815 32197
rect 27429 32194 27495 32197
rect 23749 32192 27495 32194
rect 23749 32136 23754 32192
rect 23810 32136 27434 32192
rect 27490 32136 27495 32192
rect 23749 32134 27495 32136
rect 23749 32131 23815 32134
rect 27429 32131 27495 32134
rect 4787 32128 5103 32129
rect 4787 32064 4793 32128
rect 4857 32064 4873 32128
rect 4937 32064 4953 32128
rect 5017 32064 5033 32128
rect 5097 32064 5103 32128
rect 4787 32063 5103 32064
rect 12469 32128 12785 32129
rect 12469 32064 12475 32128
rect 12539 32064 12555 32128
rect 12619 32064 12635 32128
rect 12699 32064 12715 32128
rect 12779 32064 12785 32128
rect 12469 32063 12785 32064
rect 20151 32128 20467 32129
rect 20151 32064 20157 32128
rect 20221 32064 20237 32128
rect 20301 32064 20317 32128
rect 20381 32064 20397 32128
rect 20461 32064 20467 32128
rect 20151 32063 20467 32064
rect 27833 32128 28149 32129
rect 27833 32064 27839 32128
rect 27903 32064 27919 32128
rect 27983 32064 27999 32128
rect 28063 32064 28079 32128
rect 28143 32064 28149 32128
rect 27833 32063 28149 32064
rect 20529 32058 20595 32061
rect 26182 32058 26188 32060
rect 20529 32056 26188 32058
rect 20529 32000 20534 32056
rect 20590 32000 26188 32056
rect 20529 31998 26188 32000
rect 20529 31995 20595 31998
rect 26182 31996 26188 31998
rect 26252 32058 26258 32060
rect 27705 32058 27771 32061
rect 26252 32056 27771 32058
rect 26252 32000 27710 32056
rect 27766 32000 27771 32056
rect 26252 31998 27771 32000
rect 26252 31996 26258 31998
rect 27705 31995 27771 31998
rect 8150 31860 8156 31924
rect 8220 31922 8226 31924
rect 21950 31922 21956 31924
rect 8220 31862 21956 31922
rect 8220 31860 8226 31862
rect 21950 31860 21956 31862
rect 22020 31860 22026 31924
rect 22645 31922 22711 31925
rect 25405 31922 25471 31925
rect 29637 31922 29703 31925
rect 22645 31920 29703 31922
rect 22645 31864 22650 31920
rect 22706 31864 25410 31920
rect 25466 31864 29642 31920
rect 29698 31864 29703 31920
rect 22645 31862 29703 31864
rect 22645 31859 22711 31862
rect 25405 31859 25471 31862
rect 29637 31859 29703 31862
rect 0 31696 800 31816
rect 10041 31786 10107 31789
rect 25446 31786 25452 31788
rect 10041 31784 25452 31786
rect 10041 31728 10046 31784
rect 10102 31728 25452 31784
rect 10041 31726 25452 31728
rect 10041 31723 10107 31726
rect 25446 31724 25452 31726
rect 25516 31724 25522 31788
rect 31201 31786 31267 31789
rect 32206 31786 33006 31816
rect 31201 31784 33006 31786
rect 31201 31728 31206 31784
rect 31262 31728 33006 31784
rect 31201 31726 33006 31728
rect 31201 31723 31267 31726
rect 32206 31696 33006 31726
rect 19609 31650 19675 31653
rect 23473 31650 23539 31653
rect 23841 31650 23907 31653
rect 19609 31648 23907 31650
rect 19609 31592 19614 31648
rect 19670 31592 23478 31648
rect 23534 31592 23846 31648
rect 23902 31592 23907 31648
rect 19609 31590 23907 31592
rect 19609 31587 19675 31590
rect 23473 31587 23539 31590
rect 23841 31587 23907 31590
rect 24485 31652 24551 31653
rect 24485 31648 24532 31652
rect 24596 31650 24602 31652
rect 24945 31650 25011 31653
rect 25998 31650 26004 31652
rect 24485 31592 24490 31648
rect 24485 31588 24532 31592
rect 24596 31590 24642 31650
rect 24945 31648 26004 31650
rect 24945 31592 24950 31648
rect 25006 31592 26004 31648
rect 24945 31590 26004 31592
rect 24596 31588 24602 31590
rect 24485 31587 24551 31588
rect 24945 31587 25011 31590
rect 25998 31588 26004 31590
rect 26068 31588 26074 31652
rect 27286 31588 27292 31652
rect 27356 31650 27362 31652
rect 28758 31650 28764 31652
rect 27356 31590 28764 31650
rect 27356 31588 27362 31590
rect 28758 31588 28764 31590
rect 28828 31588 28834 31652
rect 8628 31584 8944 31585
rect 8628 31520 8634 31584
rect 8698 31520 8714 31584
rect 8778 31520 8794 31584
rect 8858 31520 8874 31584
rect 8938 31520 8944 31584
rect 8628 31519 8944 31520
rect 16310 31584 16626 31585
rect 16310 31520 16316 31584
rect 16380 31520 16396 31584
rect 16460 31520 16476 31584
rect 16540 31520 16556 31584
rect 16620 31520 16626 31584
rect 16310 31519 16626 31520
rect 23992 31584 24308 31585
rect 23992 31520 23998 31584
rect 24062 31520 24078 31584
rect 24142 31520 24158 31584
rect 24222 31520 24238 31584
rect 24302 31520 24308 31584
rect 23992 31519 24308 31520
rect 31674 31584 31990 31585
rect 31674 31520 31680 31584
rect 31744 31520 31760 31584
rect 31824 31520 31840 31584
rect 31904 31520 31920 31584
rect 31984 31520 31990 31584
rect 31674 31519 31990 31520
rect 17769 31514 17835 31517
rect 22502 31514 22508 31516
rect 17588 31512 22508 31514
rect 17588 31456 17774 31512
rect 17830 31456 22508 31512
rect 17588 31454 22508 31456
rect 8201 31378 8267 31381
rect 13537 31378 13603 31381
rect 17588 31378 17648 31454
rect 17769 31451 17835 31454
rect 22502 31452 22508 31454
rect 22572 31514 22578 31516
rect 23841 31514 23907 31517
rect 22572 31512 23907 31514
rect 22572 31456 23846 31512
rect 23902 31456 23907 31512
rect 22572 31454 23907 31456
rect 22572 31452 22578 31454
rect 23841 31451 23907 31454
rect 24485 31514 24551 31517
rect 29729 31514 29795 31517
rect 24485 31512 29795 31514
rect 24485 31456 24490 31512
rect 24546 31456 29734 31512
rect 29790 31456 29795 31512
rect 24485 31454 29795 31456
rect 24485 31451 24551 31454
rect 29729 31451 29795 31454
rect 8201 31376 17648 31378
rect 8201 31320 8206 31376
rect 8262 31320 13542 31376
rect 13598 31320 17648 31376
rect 8201 31318 17648 31320
rect 8201 31315 8267 31318
rect 13537 31315 13603 31318
rect 17718 31316 17724 31380
rect 17788 31378 17794 31380
rect 25221 31378 25287 31381
rect 32254 31378 32260 31380
rect 17788 31376 25287 31378
rect 17788 31320 25226 31376
rect 25282 31320 25287 31376
rect 17788 31318 25287 31320
rect 17788 31316 17794 31318
rect 25221 31315 25287 31318
rect 25408 31318 32260 31378
rect 10726 31180 10732 31244
rect 10796 31242 10802 31244
rect 13169 31242 13235 31245
rect 10796 31240 13235 31242
rect 10796 31184 13174 31240
rect 13230 31184 13235 31240
rect 10796 31182 13235 31184
rect 10796 31180 10802 31182
rect 13169 31179 13235 31182
rect 16113 31242 16179 31245
rect 22686 31242 22692 31244
rect 16113 31240 22692 31242
rect 16113 31184 16118 31240
rect 16174 31184 22692 31240
rect 16113 31182 22692 31184
rect 16113 31179 16179 31182
rect 22686 31180 22692 31182
rect 22756 31242 22762 31244
rect 25408 31242 25468 31318
rect 32254 31316 32260 31318
rect 32324 31316 32330 31380
rect 22756 31182 25468 31242
rect 27061 31242 27127 31245
rect 30782 31242 30788 31244
rect 27061 31240 30788 31242
rect 27061 31184 27066 31240
rect 27122 31184 30788 31240
rect 27061 31182 30788 31184
rect 22756 31180 22762 31182
rect 27061 31179 27127 31182
rect 30782 31180 30788 31182
rect 30852 31180 30858 31244
rect 14733 31106 14799 31109
rect 18086 31106 18092 31108
rect 14733 31104 18092 31106
rect 14733 31048 14738 31104
rect 14794 31048 18092 31104
rect 14733 31046 18092 31048
rect 14733 31043 14799 31046
rect 18086 31044 18092 31046
rect 18156 31106 18162 31108
rect 19977 31106 20043 31109
rect 18156 31104 20043 31106
rect 18156 31048 19982 31104
rect 20038 31048 20043 31104
rect 18156 31046 20043 31048
rect 18156 31044 18162 31046
rect 19977 31043 20043 31046
rect 20713 31106 20779 31109
rect 22645 31106 22711 31109
rect 20713 31104 22711 31106
rect 20713 31048 20718 31104
rect 20774 31048 22650 31104
rect 22706 31048 22711 31104
rect 20713 31046 22711 31048
rect 20713 31043 20779 31046
rect 22645 31043 22711 31046
rect 23289 31106 23355 31109
rect 25262 31106 25268 31108
rect 23289 31104 25268 31106
rect 23289 31048 23294 31104
rect 23350 31048 25268 31104
rect 23289 31046 25268 31048
rect 23289 31043 23355 31046
rect 25262 31044 25268 31046
rect 25332 31044 25338 31108
rect 25497 31106 25563 31109
rect 27337 31106 27403 31109
rect 25497 31104 27403 31106
rect 25497 31048 25502 31104
rect 25558 31048 27342 31104
rect 27398 31048 27403 31104
rect 25497 31046 27403 31048
rect 25497 31043 25563 31046
rect 27337 31043 27403 31046
rect 28717 31106 28783 31109
rect 29310 31106 29316 31108
rect 28717 31104 29316 31106
rect 28717 31048 28722 31104
rect 28778 31048 29316 31104
rect 28717 31046 29316 31048
rect 28717 31043 28783 31046
rect 29310 31044 29316 31046
rect 29380 31044 29386 31108
rect 4787 31040 5103 31041
rect 0 30970 800 31000
rect 4787 30976 4793 31040
rect 4857 30976 4873 31040
rect 4937 30976 4953 31040
rect 5017 30976 5033 31040
rect 5097 30976 5103 31040
rect 4787 30975 5103 30976
rect 12469 31040 12785 31041
rect 12469 30976 12475 31040
rect 12539 30976 12555 31040
rect 12619 30976 12635 31040
rect 12699 30976 12715 31040
rect 12779 30976 12785 31040
rect 12469 30975 12785 30976
rect 20151 31040 20467 31041
rect 20151 30976 20157 31040
rect 20221 30976 20237 31040
rect 20301 30976 20317 31040
rect 20381 30976 20397 31040
rect 20461 30976 20467 31040
rect 20151 30975 20467 30976
rect 27833 31040 28149 31041
rect 27833 30976 27839 31040
rect 27903 30976 27919 31040
rect 27983 30976 27999 31040
rect 28063 30976 28079 31040
rect 28143 30976 28149 31040
rect 32206 31016 33006 31136
rect 27833 30975 28149 30976
rect 1577 30970 1643 30973
rect 0 30968 1643 30970
rect 0 30912 1582 30968
rect 1638 30912 1643 30968
rect 0 30910 1643 30912
rect 0 30880 800 30910
rect 1577 30907 1643 30910
rect 14222 30908 14228 30972
rect 14292 30970 14298 30972
rect 14917 30970 14983 30973
rect 14292 30968 14983 30970
rect 14292 30912 14922 30968
rect 14978 30912 14983 30968
rect 14292 30910 14983 30912
rect 14292 30908 14298 30910
rect 14917 30907 14983 30910
rect 15510 30908 15516 30972
rect 15580 30970 15586 30972
rect 16205 30970 16271 30973
rect 15580 30968 16271 30970
rect 15580 30912 16210 30968
rect 16266 30912 16271 30968
rect 15580 30910 16271 30912
rect 15580 30908 15586 30910
rect 16205 30907 16271 30910
rect 20529 30970 20595 30973
rect 26509 30970 26575 30973
rect 28441 30972 28507 30973
rect 20529 30968 26575 30970
rect 20529 30912 20534 30968
rect 20590 30912 26514 30968
rect 26570 30912 26575 30968
rect 20529 30910 26575 30912
rect 20529 30907 20595 30910
rect 26509 30907 26575 30910
rect 28390 30908 28396 30972
rect 28460 30970 28507 30972
rect 28460 30968 28552 30970
rect 28502 30912 28552 30968
rect 28460 30910 28552 30912
rect 28460 30908 28507 30910
rect 28441 30907 28507 30908
rect 6678 30772 6684 30836
rect 6748 30834 6754 30836
rect 11421 30834 11487 30837
rect 17217 30834 17283 30837
rect 19241 30834 19307 30837
rect 19742 30834 19748 30836
rect 6748 30832 17283 30834
rect 6748 30776 11426 30832
rect 11482 30776 17222 30832
rect 17278 30776 17283 30832
rect 6748 30774 17283 30776
rect 6748 30772 6754 30774
rect 11421 30771 11487 30774
rect 17217 30771 17283 30774
rect 17542 30832 19748 30834
rect 17542 30776 19246 30832
rect 19302 30776 19748 30832
rect 17542 30774 19748 30776
rect 6862 30636 6868 30700
rect 6932 30698 6938 30700
rect 6932 30638 10242 30698
rect 6932 30636 6938 30638
rect 10182 30562 10242 30638
rect 11462 30636 11468 30700
rect 11532 30698 11538 30700
rect 17125 30698 17191 30701
rect 17542 30698 17602 30774
rect 19241 30771 19307 30774
rect 19742 30772 19748 30774
rect 19812 30772 19818 30836
rect 20345 30834 20411 30837
rect 23657 30834 23723 30837
rect 24761 30834 24827 30837
rect 25814 30834 25820 30836
rect 20345 30832 24594 30834
rect 20345 30776 20350 30832
rect 20406 30776 23662 30832
rect 23718 30776 24594 30832
rect 20345 30774 24594 30776
rect 20345 30771 20411 30774
rect 23657 30771 23723 30774
rect 11532 30696 17602 30698
rect 11532 30640 17130 30696
rect 17186 30640 17602 30696
rect 11532 30638 17602 30640
rect 18965 30698 19031 30701
rect 19190 30698 19196 30700
rect 18965 30696 19196 30698
rect 18965 30640 18970 30696
rect 19026 30640 19196 30696
rect 18965 30638 19196 30640
rect 11532 30636 11538 30638
rect 17125 30635 17191 30638
rect 18965 30635 19031 30638
rect 19190 30636 19196 30638
rect 19260 30636 19266 30700
rect 20069 30698 20135 30701
rect 24534 30698 24594 30774
rect 24761 30832 25820 30834
rect 24761 30776 24766 30832
rect 24822 30776 25820 30832
rect 24761 30774 25820 30776
rect 24761 30771 24827 30774
rect 25814 30772 25820 30774
rect 25884 30834 25890 30836
rect 26141 30834 26207 30837
rect 25884 30832 26207 30834
rect 25884 30776 26146 30832
rect 26202 30776 26207 30832
rect 25884 30774 26207 30776
rect 25884 30772 25890 30774
rect 26141 30771 26207 30774
rect 26785 30834 26851 30837
rect 27470 30834 27476 30836
rect 26785 30832 27476 30834
rect 26785 30776 26790 30832
rect 26846 30776 27476 30832
rect 26785 30774 27476 30776
rect 26785 30771 26851 30774
rect 27470 30772 27476 30774
rect 27540 30834 27546 30836
rect 28349 30834 28415 30837
rect 30414 30834 30420 30836
rect 27540 30832 28415 30834
rect 27540 30776 28354 30832
rect 28410 30776 28415 30832
rect 27540 30774 28415 30776
rect 27540 30772 27546 30774
rect 28349 30771 28415 30774
rect 28536 30774 30420 30834
rect 27102 30698 27108 30700
rect 20069 30696 24456 30698
rect 20069 30640 20074 30696
rect 20130 30640 24456 30696
rect 20069 30638 24456 30640
rect 24534 30638 27108 30698
rect 20069 30635 20135 30638
rect 16113 30562 16179 30565
rect 10182 30560 16179 30562
rect 10182 30504 16118 30560
rect 16174 30504 16179 30560
rect 10182 30502 16179 30504
rect 16113 30499 16179 30502
rect 16849 30562 16915 30565
rect 20345 30562 20411 30565
rect 16849 30560 20411 30562
rect 16849 30504 16854 30560
rect 16910 30504 20350 30560
rect 20406 30504 20411 30560
rect 16849 30502 20411 30504
rect 16849 30499 16915 30502
rect 20345 30499 20411 30502
rect 20989 30562 21055 30565
rect 22185 30562 22251 30565
rect 20989 30560 22251 30562
rect 20989 30504 20994 30560
rect 21050 30504 22190 30560
rect 22246 30504 22251 30560
rect 20989 30502 22251 30504
rect 20989 30499 21055 30502
rect 22185 30499 22251 30502
rect 23422 30500 23428 30564
rect 23492 30562 23498 30564
rect 23749 30562 23815 30565
rect 23492 30560 23815 30562
rect 23492 30504 23754 30560
rect 23810 30504 23815 30560
rect 23492 30502 23815 30504
rect 24396 30562 24456 30638
rect 27102 30636 27108 30638
rect 27172 30636 27178 30700
rect 27337 30698 27403 30701
rect 28536 30698 28596 30774
rect 30414 30772 30420 30774
rect 30484 30772 30490 30836
rect 27337 30696 28596 30698
rect 27337 30640 27342 30696
rect 27398 30640 28596 30696
rect 27337 30638 28596 30640
rect 30005 30698 30071 30701
rect 30005 30696 32138 30698
rect 30005 30640 30010 30696
rect 30066 30640 32138 30696
rect 30005 30638 32138 30640
rect 27337 30635 27403 30638
rect 30005 30635 30071 30638
rect 24945 30562 25011 30565
rect 26325 30562 26391 30565
rect 26734 30562 26740 30564
rect 24396 30560 25468 30562
rect 24396 30504 24950 30560
rect 25006 30504 25468 30560
rect 24396 30502 25468 30504
rect 23492 30500 23498 30502
rect 23749 30499 23815 30502
rect 24945 30499 25011 30502
rect 8628 30496 8944 30497
rect 8628 30432 8634 30496
rect 8698 30432 8714 30496
rect 8778 30432 8794 30496
rect 8858 30432 8874 30496
rect 8938 30432 8944 30496
rect 8628 30431 8944 30432
rect 16310 30496 16626 30497
rect 16310 30432 16316 30496
rect 16380 30432 16396 30496
rect 16460 30432 16476 30496
rect 16540 30432 16556 30496
rect 16620 30432 16626 30496
rect 16310 30431 16626 30432
rect 23992 30496 24308 30497
rect 23992 30432 23998 30496
rect 24062 30432 24078 30496
rect 24142 30432 24158 30496
rect 24222 30432 24238 30496
rect 24302 30432 24308 30496
rect 23992 30431 24308 30432
rect 11830 30364 11836 30428
rect 11900 30426 11906 30428
rect 12801 30426 12867 30429
rect 11900 30424 12867 30426
rect 11900 30368 12806 30424
rect 12862 30368 12867 30424
rect 11900 30366 12867 30368
rect 11900 30364 11906 30366
rect 12801 30363 12867 30366
rect 13353 30426 13419 30429
rect 14406 30426 14412 30428
rect 13353 30424 14412 30426
rect 13353 30368 13358 30424
rect 13414 30368 14412 30424
rect 13353 30366 14412 30368
rect 13353 30363 13419 30366
rect 14406 30364 14412 30366
rect 14476 30364 14482 30428
rect 19006 30364 19012 30428
rect 19076 30426 19082 30428
rect 19333 30426 19399 30429
rect 19076 30424 19399 30426
rect 19076 30368 19338 30424
rect 19394 30368 19399 30424
rect 19076 30366 19399 30368
rect 19076 30364 19082 30366
rect 19333 30363 19399 30366
rect 19926 30364 19932 30428
rect 19996 30426 20002 30428
rect 20253 30426 20319 30429
rect 19996 30424 20319 30426
rect 19996 30368 20258 30424
rect 20314 30368 20319 30424
rect 19996 30366 20319 30368
rect 19996 30364 20002 30366
rect 20253 30363 20319 30366
rect 20437 30426 20503 30429
rect 21030 30426 21036 30428
rect 20437 30424 21036 30426
rect 20437 30368 20442 30424
rect 20498 30368 21036 30424
rect 20437 30366 21036 30368
rect 20437 30363 20503 30366
rect 21030 30364 21036 30366
rect 21100 30364 21106 30428
rect 21541 30426 21607 30429
rect 23749 30426 23815 30429
rect 21541 30424 23815 30426
rect 21541 30368 21546 30424
rect 21602 30368 23754 30424
rect 23810 30368 23815 30424
rect 21541 30366 23815 30368
rect 21541 30363 21607 30366
rect 23749 30363 23815 30366
rect 24485 30426 24551 30429
rect 25221 30426 25287 30429
rect 24485 30424 25287 30426
rect 24485 30368 24490 30424
rect 24546 30368 25226 30424
rect 25282 30368 25287 30424
rect 24485 30366 25287 30368
rect 25408 30426 25468 30502
rect 26325 30560 26740 30562
rect 26325 30504 26330 30560
rect 26386 30504 26740 30560
rect 26325 30502 26740 30504
rect 26325 30499 26391 30502
rect 26734 30500 26740 30502
rect 26804 30500 26810 30564
rect 26918 30500 26924 30564
rect 26988 30562 26994 30564
rect 30925 30562 30991 30565
rect 26988 30560 30991 30562
rect 26988 30504 30930 30560
rect 30986 30504 30991 30560
rect 26988 30502 30991 30504
rect 26988 30500 26994 30502
rect 30925 30499 30991 30502
rect 31674 30496 31990 30497
rect 31674 30432 31680 30496
rect 31744 30432 31760 30496
rect 31824 30432 31840 30496
rect 31904 30432 31920 30496
rect 31984 30432 31990 30496
rect 31674 30431 31990 30432
rect 27654 30426 27660 30428
rect 25408 30366 27660 30426
rect 24485 30363 24551 30366
rect 25221 30363 25287 30366
rect 27654 30364 27660 30366
rect 27724 30364 27730 30428
rect 27889 30426 27955 30429
rect 28349 30426 28415 30429
rect 30557 30428 30623 30429
rect 30557 30426 30604 30428
rect 27889 30424 28415 30426
rect 27889 30368 27894 30424
rect 27950 30368 28354 30424
rect 28410 30368 28415 30424
rect 27889 30366 28415 30368
rect 30512 30424 30604 30426
rect 30512 30368 30562 30424
rect 30512 30366 30604 30368
rect 27889 30363 27955 30366
rect 28349 30363 28415 30366
rect 30557 30364 30604 30366
rect 30668 30364 30674 30428
rect 32078 30426 32138 30638
rect 32206 30426 33006 30456
rect 32078 30366 33006 30426
rect 30557 30363 30623 30364
rect 32206 30336 33006 30366
rect 13353 30290 13419 30293
rect 18137 30290 18203 30293
rect 13353 30288 18203 30290
rect 13353 30232 13358 30288
rect 13414 30232 18142 30288
rect 18198 30232 18203 30288
rect 13353 30230 18203 30232
rect 13353 30227 13419 30230
rect 18137 30227 18203 30230
rect 19374 30228 19380 30292
rect 19444 30290 19450 30292
rect 19517 30290 19583 30293
rect 19444 30288 19583 30290
rect 19444 30232 19522 30288
rect 19578 30232 19583 30288
rect 19444 30230 19583 30232
rect 19444 30228 19450 30230
rect 19517 30227 19583 30230
rect 19885 30290 19951 30293
rect 20713 30290 20779 30293
rect 19885 30288 20779 30290
rect 19885 30232 19890 30288
rect 19946 30232 20718 30288
rect 20774 30232 20779 30288
rect 19885 30230 20779 30232
rect 19885 30227 19951 30230
rect 20713 30227 20779 30230
rect 20897 30290 20963 30293
rect 22870 30290 22876 30292
rect 20897 30288 22876 30290
rect 20897 30232 20902 30288
rect 20958 30232 22876 30288
rect 20897 30230 22876 30232
rect 20897 30227 20963 30230
rect 22870 30228 22876 30230
rect 22940 30228 22946 30292
rect 23197 30290 23263 30293
rect 23197 30288 32138 30290
rect 23197 30232 23202 30288
rect 23258 30232 32138 30288
rect 23197 30230 32138 30232
rect 23197 30227 23263 30230
rect 0 30154 800 30184
rect 1577 30154 1643 30157
rect 0 30152 1643 30154
rect 0 30096 1582 30152
rect 1638 30096 1643 30152
rect 0 30094 1643 30096
rect 0 30064 800 30094
rect 1577 30091 1643 30094
rect 7046 30092 7052 30156
rect 7116 30154 7122 30156
rect 9949 30154 10015 30157
rect 15142 30154 15148 30156
rect 7116 30152 15148 30154
rect 7116 30096 9954 30152
rect 10010 30096 15148 30152
rect 7116 30094 15148 30096
rect 7116 30092 7122 30094
rect 9949 30091 10015 30094
rect 15142 30092 15148 30094
rect 15212 30092 15218 30156
rect 15377 30154 15443 30157
rect 15837 30154 15903 30157
rect 24945 30154 25011 30157
rect 15377 30152 25011 30154
rect 15377 30096 15382 30152
rect 15438 30096 15842 30152
rect 15898 30096 24950 30152
rect 25006 30096 25011 30152
rect 15377 30094 25011 30096
rect 15377 30091 15443 30094
rect 15837 30091 15903 30094
rect 24945 30091 25011 30094
rect 25078 30092 25084 30156
rect 25148 30154 25154 30156
rect 25221 30154 25287 30157
rect 25148 30152 25287 30154
rect 25148 30096 25226 30152
rect 25282 30096 25287 30152
rect 25148 30094 25287 30096
rect 25148 30092 25154 30094
rect 25221 30091 25287 30094
rect 25630 30092 25636 30156
rect 25700 30154 25706 30156
rect 31477 30154 31543 30157
rect 25700 30152 31543 30154
rect 25700 30096 31482 30152
rect 31538 30096 31543 30152
rect 25700 30094 31543 30096
rect 32078 30154 32138 30230
rect 32581 30154 32647 30157
rect 32078 30152 32647 30154
rect 32078 30096 32586 30152
rect 32642 30096 32647 30152
rect 32078 30094 32647 30096
rect 25700 30092 25706 30094
rect 31477 30091 31543 30094
rect 32581 30091 32647 30094
rect 17902 29956 17908 30020
rect 17972 30018 17978 30020
rect 19425 30018 19491 30021
rect 17972 30016 19491 30018
rect 17972 29960 19430 30016
rect 19486 29960 19491 30016
rect 17972 29958 19491 29960
rect 17972 29956 17978 29958
rect 19425 29955 19491 29958
rect 20621 30018 20687 30021
rect 23197 30018 23263 30021
rect 20621 30016 23263 30018
rect 20621 29960 20626 30016
rect 20682 29960 23202 30016
rect 23258 29960 23263 30016
rect 20621 29958 23263 29960
rect 20621 29955 20687 29958
rect 23197 29955 23263 29958
rect 23933 30018 23999 30021
rect 26049 30018 26115 30021
rect 23933 30016 26115 30018
rect 23933 29960 23938 30016
rect 23994 29960 26054 30016
rect 26110 29960 26115 30016
rect 23933 29958 26115 29960
rect 23933 29955 23999 29958
rect 26049 29955 26115 29958
rect 26325 30020 26391 30021
rect 26325 30016 26372 30020
rect 26436 30018 26442 30020
rect 27061 30018 27127 30021
rect 27286 30018 27292 30020
rect 26325 29960 26330 30016
rect 26325 29956 26372 29960
rect 26436 29958 26482 30018
rect 27061 30016 27292 30018
rect 27061 29960 27066 30016
rect 27122 29960 27292 30016
rect 27061 29958 27292 29960
rect 26436 29956 26442 29958
rect 26325 29955 26391 29956
rect 27061 29955 27127 29958
rect 27286 29956 27292 29958
rect 27356 29956 27362 30020
rect 28252 29956 28258 30020
rect 28322 30018 28328 30020
rect 32622 30018 32628 30020
rect 28322 29958 32628 30018
rect 28322 29956 28328 29958
rect 32622 29956 32628 29958
rect 32692 29956 32698 30020
rect 4787 29952 5103 29953
rect 4787 29888 4793 29952
rect 4857 29888 4873 29952
rect 4937 29888 4953 29952
rect 5017 29888 5033 29952
rect 5097 29888 5103 29952
rect 4787 29887 5103 29888
rect 12469 29952 12785 29953
rect 12469 29888 12475 29952
rect 12539 29888 12555 29952
rect 12619 29888 12635 29952
rect 12699 29888 12715 29952
rect 12779 29888 12785 29952
rect 12469 29887 12785 29888
rect 20151 29952 20467 29953
rect 20151 29888 20157 29952
rect 20221 29888 20237 29952
rect 20301 29888 20317 29952
rect 20381 29888 20397 29952
rect 20461 29888 20467 29952
rect 20151 29887 20467 29888
rect 27833 29952 28149 29953
rect 27833 29888 27839 29952
rect 27903 29888 27919 29952
rect 27983 29888 27999 29952
rect 28063 29888 28079 29952
rect 28143 29888 28149 29952
rect 27833 29887 28149 29888
rect 17166 29820 17172 29884
rect 17236 29882 17242 29884
rect 19885 29882 19951 29885
rect 24761 29882 24827 29885
rect 26785 29882 26851 29885
rect 27337 29884 27403 29885
rect 27286 29882 27292 29884
rect 17236 29880 19951 29882
rect 17236 29824 19890 29880
rect 19946 29824 19951 29880
rect 17236 29822 19951 29824
rect 17236 29820 17242 29822
rect 19885 29819 19951 29822
rect 20532 29880 26851 29882
rect 20532 29824 24766 29880
rect 24822 29824 26790 29880
rect 26846 29824 26851 29880
rect 20532 29822 26851 29824
rect 27246 29822 27292 29882
rect 27356 29880 27403 29884
rect 27398 29824 27403 29880
rect 4521 29746 4587 29749
rect 12801 29746 12867 29749
rect 12934 29746 12940 29748
rect 4521 29744 9690 29746
rect 4521 29688 4526 29744
rect 4582 29688 9690 29744
rect 4521 29686 9690 29688
rect 4521 29683 4587 29686
rect 9630 29610 9690 29686
rect 12801 29744 12940 29746
rect 12801 29688 12806 29744
rect 12862 29688 12940 29744
rect 12801 29686 12940 29688
rect 12801 29683 12867 29686
rect 12934 29684 12940 29686
rect 13004 29684 13010 29748
rect 18270 29684 18276 29748
rect 18340 29746 18346 29748
rect 18781 29746 18847 29749
rect 20532 29746 20592 29822
rect 24761 29819 24827 29822
rect 26785 29819 26851 29822
rect 27286 29820 27292 29822
rect 27356 29820 27403 29824
rect 27337 29819 27403 29820
rect 28441 29882 28507 29885
rect 29494 29882 29500 29884
rect 28441 29880 29500 29882
rect 28441 29824 28446 29880
rect 28502 29824 29500 29880
rect 28441 29822 29500 29824
rect 28441 29819 28507 29822
rect 29494 29820 29500 29822
rect 29564 29820 29570 29884
rect 18340 29744 20592 29746
rect 18340 29688 18786 29744
rect 18842 29688 20592 29744
rect 18340 29686 20592 29688
rect 20805 29746 20871 29749
rect 21449 29746 21515 29749
rect 21766 29746 21772 29748
rect 20805 29744 21772 29746
rect 20805 29688 20810 29744
rect 20866 29688 21454 29744
rect 21510 29688 21772 29744
rect 20805 29686 21772 29688
rect 18340 29684 18346 29686
rect 18781 29683 18847 29686
rect 20805 29683 20871 29686
rect 21449 29683 21515 29686
rect 21766 29684 21772 29686
rect 21836 29684 21842 29748
rect 22185 29746 22251 29749
rect 24669 29746 24735 29749
rect 22185 29744 24735 29746
rect 22185 29688 22190 29744
rect 22246 29688 24674 29744
rect 24730 29688 24735 29744
rect 22185 29686 24735 29688
rect 22185 29683 22251 29686
rect 24669 29683 24735 29686
rect 24853 29746 24919 29749
rect 25078 29746 25084 29748
rect 24853 29744 25084 29746
rect 24853 29688 24858 29744
rect 24914 29688 25084 29744
rect 24853 29686 25084 29688
rect 24853 29683 24919 29686
rect 25078 29684 25084 29686
rect 25148 29684 25154 29748
rect 25221 29746 25287 29749
rect 25446 29746 25452 29748
rect 25221 29744 25452 29746
rect 25221 29688 25226 29744
rect 25282 29688 25452 29744
rect 25221 29686 25452 29688
rect 25221 29683 25287 29686
rect 25446 29684 25452 29686
rect 25516 29746 25522 29748
rect 28073 29746 28139 29749
rect 25516 29744 28139 29746
rect 25516 29688 28078 29744
rect 28134 29688 28139 29744
rect 25516 29686 28139 29688
rect 25516 29684 25522 29686
rect 28073 29683 28139 29686
rect 28257 29746 28323 29749
rect 28574 29746 28580 29748
rect 28257 29744 28580 29746
rect 28257 29688 28262 29744
rect 28318 29688 28580 29744
rect 28257 29686 28580 29688
rect 28257 29683 28323 29686
rect 28574 29684 28580 29686
rect 28644 29684 28650 29748
rect 31201 29746 31267 29749
rect 32206 29746 33006 29776
rect 28812 29686 31080 29746
rect 18505 29610 18571 29613
rect 18689 29610 18755 29613
rect 9630 29608 18755 29610
rect 9630 29552 18510 29608
rect 18566 29552 18694 29608
rect 18750 29552 18755 29608
rect 9630 29550 18755 29552
rect 18505 29547 18571 29550
rect 18689 29547 18755 29550
rect 19333 29610 19399 29613
rect 20621 29610 20687 29613
rect 22369 29610 22435 29613
rect 22502 29610 22508 29612
rect 19333 29608 20132 29610
rect 19333 29552 19338 29608
rect 19394 29552 20132 29608
rect 19333 29550 20132 29552
rect 19333 29547 19399 29550
rect 17217 29474 17283 29477
rect 17534 29474 17540 29476
rect 17217 29472 17540 29474
rect 17217 29416 17222 29472
rect 17278 29416 17540 29472
rect 17217 29414 17540 29416
rect 17217 29411 17283 29414
rect 17534 29412 17540 29414
rect 17604 29412 17610 29476
rect 17769 29474 17835 29477
rect 19885 29474 19951 29477
rect 17769 29472 19951 29474
rect 17769 29416 17774 29472
rect 17830 29416 19890 29472
rect 19946 29416 19951 29472
rect 17769 29414 19951 29416
rect 20072 29474 20132 29550
rect 20621 29608 22110 29610
rect 20621 29552 20626 29608
rect 20682 29552 22110 29608
rect 20621 29550 22110 29552
rect 20621 29547 20687 29550
rect 20989 29474 21055 29477
rect 21449 29476 21515 29477
rect 20072 29472 21055 29474
rect 20072 29416 20994 29472
rect 21050 29416 21055 29472
rect 20072 29414 21055 29416
rect 17769 29411 17835 29414
rect 19885 29411 19951 29414
rect 20989 29411 21055 29414
rect 21398 29412 21404 29476
rect 21468 29474 21515 29476
rect 22050 29474 22110 29550
rect 22369 29608 22508 29610
rect 22369 29552 22374 29608
rect 22430 29552 22508 29608
rect 22369 29550 22508 29552
rect 22369 29547 22435 29550
rect 22502 29548 22508 29550
rect 22572 29548 22578 29612
rect 22921 29610 22987 29613
rect 25773 29610 25839 29613
rect 22921 29608 25839 29610
rect 22921 29552 22926 29608
rect 22982 29552 25778 29608
rect 25834 29552 25839 29608
rect 22921 29550 25839 29552
rect 22921 29547 22987 29550
rect 25773 29547 25839 29550
rect 26141 29610 26207 29613
rect 27981 29610 28047 29613
rect 28812 29610 28872 29686
rect 26141 29608 27906 29610
rect 26141 29552 26146 29608
rect 26202 29552 27906 29608
rect 26141 29550 27906 29552
rect 26141 29547 26207 29550
rect 23054 29474 23060 29476
rect 21468 29472 21560 29474
rect 21510 29416 21560 29472
rect 21468 29414 21560 29416
rect 22050 29414 23060 29474
rect 21468 29412 21515 29414
rect 23054 29412 23060 29414
rect 23124 29412 23130 29476
rect 23289 29474 23355 29477
rect 23749 29474 23815 29477
rect 23289 29472 23815 29474
rect 23289 29416 23294 29472
rect 23350 29416 23754 29472
rect 23810 29416 23815 29472
rect 23289 29414 23815 29416
rect 21449 29411 21515 29412
rect 23289 29411 23355 29414
rect 23749 29411 23815 29414
rect 24945 29474 25011 29477
rect 25221 29474 25287 29477
rect 25589 29476 25655 29477
rect 25446 29474 25452 29476
rect 24945 29472 25452 29474
rect 24945 29416 24950 29472
rect 25006 29416 25226 29472
rect 25282 29416 25452 29472
rect 24945 29414 25452 29416
rect 24945 29411 25011 29414
rect 25221 29411 25287 29414
rect 25446 29412 25452 29414
rect 25516 29412 25522 29476
rect 25589 29472 25636 29476
rect 25700 29474 25706 29476
rect 25589 29416 25594 29472
rect 25589 29412 25636 29416
rect 25700 29414 25746 29474
rect 25700 29412 25706 29414
rect 25998 29412 26004 29476
rect 26068 29474 26074 29476
rect 26141 29474 26207 29477
rect 26068 29472 26207 29474
rect 26068 29416 26146 29472
rect 26202 29416 26207 29472
rect 26068 29414 26207 29416
rect 26068 29412 26074 29414
rect 25589 29411 25655 29412
rect 26141 29411 26207 29414
rect 26509 29474 26575 29477
rect 26918 29474 26924 29476
rect 26509 29472 26924 29474
rect 26509 29416 26514 29472
rect 26570 29416 26924 29472
rect 26509 29414 26924 29416
rect 26509 29411 26575 29414
rect 26918 29412 26924 29414
rect 26988 29412 26994 29476
rect 27061 29474 27127 29477
rect 27429 29474 27495 29477
rect 27061 29472 27495 29474
rect 27061 29416 27066 29472
rect 27122 29416 27434 29472
rect 27490 29416 27495 29472
rect 27061 29414 27495 29416
rect 27846 29474 27906 29550
rect 27981 29608 28872 29610
rect 27981 29552 27986 29608
rect 28042 29552 28872 29608
rect 27981 29550 28872 29552
rect 27981 29547 28047 29550
rect 28942 29548 28948 29612
rect 29012 29610 29018 29612
rect 29913 29610 29979 29613
rect 29012 29608 29979 29610
rect 29012 29552 29918 29608
rect 29974 29552 29979 29608
rect 29012 29550 29979 29552
rect 31020 29610 31080 29686
rect 31201 29744 33006 29746
rect 31201 29688 31206 29744
rect 31262 29688 33006 29744
rect 31201 29686 33006 29688
rect 31201 29683 31267 29686
rect 32206 29656 33006 29686
rect 31150 29610 31156 29612
rect 31020 29550 31156 29610
rect 29012 29548 29018 29550
rect 29913 29547 29979 29550
rect 31150 29548 31156 29550
rect 31220 29548 31226 29612
rect 28257 29474 28323 29477
rect 29126 29474 29132 29476
rect 27846 29472 29132 29474
rect 27846 29416 28262 29472
rect 28318 29416 29132 29472
rect 27846 29414 29132 29416
rect 27061 29411 27127 29414
rect 27429 29411 27495 29414
rect 28257 29411 28323 29414
rect 29126 29412 29132 29414
rect 29196 29412 29202 29476
rect 8628 29408 8944 29409
rect 0 29248 800 29368
rect 8628 29344 8634 29408
rect 8698 29344 8714 29408
rect 8778 29344 8794 29408
rect 8858 29344 8874 29408
rect 8938 29344 8944 29408
rect 8628 29343 8944 29344
rect 16310 29408 16626 29409
rect 16310 29344 16316 29408
rect 16380 29344 16396 29408
rect 16460 29344 16476 29408
rect 16540 29344 16556 29408
rect 16620 29344 16626 29408
rect 16310 29343 16626 29344
rect 23992 29408 24308 29409
rect 23992 29344 23998 29408
rect 24062 29344 24078 29408
rect 24142 29344 24158 29408
rect 24222 29344 24238 29408
rect 24302 29344 24308 29408
rect 23992 29343 24308 29344
rect 31674 29408 31990 29409
rect 31674 29344 31680 29408
rect 31744 29344 31760 29408
rect 31824 29344 31840 29408
rect 31904 29344 31920 29408
rect 31984 29344 31990 29408
rect 31674 29343 31990 29344
rect 13486 29276 13492 29340
rect 13556 29338 13562 29340
rect 14365 29338 14431 29341
rect 13556 29336 14431 29338
rect 13556 29280 14370 29336
rect 14426 29280 14431 29336
rect 13556 29278 14431 29280
rect 13556 29276 13562 29278
rect 14365 29275 14431 29278
rect 16757 29338 16823 29341
rect 18597 29338 18663 29341
rect 20805 29338 20871 29341
rect 16757 29336 20871 29338
rect 16757 29280 16762 29336
rect 16818 29280 18602 29336
rect 18658 29280 20810 29336
rect 20866 29280 20871 29336
rect 16757 29278 20871 29280
rect 16757 29275 16823 29278
rect 18597 29275 18663 29278
rect 20805 29275 20871 29278
rect 21214 29276 21220 29340
rect 21284 29338 21290 29340
rect 21582 29338 21588 29340
rect 21284 29278 21588 29338
rect 21284 29276 21290 29278
rect 21582 29276 21588 29278
rect 21652 29276 21658 29340
rect 21950 29276 21956 29340
rect 22020 29338 22026 29340
rect 23013 29338 23079 29341
rect 22020 29336 23079 29338
rect 22020 29280 23018 29336
rect 23074 29280 23079 29336
rect 22020 29278 23079 29280
rect 22020 29276 22026 29278
rect 23013 29275 23079 29278
rect 23197 29340 23263 29341
rect 23657 29340 23723 29341
rect 23197 29336 23244 29340
rect 23308 29338 23314 29340
rect 23606 29338 23612 29340
rect 23197 29280 23202 29336
rect 23197 29276 23244 29280
rect 23308 29278 23354 29338
rect 23566 29278 23612 29338
rect 23676 29336 23723 29340
rect 23718 29280 23723 29336
rect 23308 29276 23314 29278
rect 23606 29276 23612 29278
rect 23676 29276 23723 29280
rect 23197 29275 23263 29276
rect 23657 29275 23723 29276
rect 24669 29338 24735 29341
rect 26233 29338 26299 29341
rect 27521 29338 27587 29341
rect 28206 29338 28212 29340
rect 24669 29336 28212 29338
rect 24669 29280 24674 29336
rect 24730 29280 26238 29336
rect 26294 29280 27526 29336
rect 27582 29280 28212 29336
rect 24669 29278 28212 29280
rect 24669 29275 24735 29278
rect 26233 29275 26299 29278
rect 27521 29275 27587 29278
rect 28206 29276 28212 29278
rect 28276 29276 28282 29340
rect 28993 29338 29059 29341
rect 29678 29338 29684 29340
rect 28993 29336 29684 29338
rect 28993 29280 28998 29336
rect 29054 29280 29684 29336
rect 28993 29278 29684 29280
rect 28993 29275 29059 29278
rect 29678 29276 29684 29278
rect 29748 29276 29754 29340
rect 32673 29338 32739 29341
rect 32078 29336 32739 29338
rect 32078 29280 32678 29336
rect 32734 29280 32739 29336
rect 32078 29278 32739 29280
rect 7373 29202 7439 29205
rect 12893 29202 12959 29205
rect 15745 29202 15811 29205
rect 19241 29202 19307 29205
rect 19926 29202 19932 29204
rect 7373 29200 12450 29202
rect 7373 29144 7378 29200
rect 7434 29144 12450 29200
rect 7373 29142 12450 29144
rect 7373 29139 7439 29142
rect 9438 29004 9444 29068
rect 9508 29066 9514 29068
rect 9949 29066 10015 29069
rect 9508 29064 10015 29066
rect 9508 29008 9954 29064
rect 10010 29008 10015 29064
rect 9508 29006 10015 29008
rect 12390 29066 12450 29142
rect 12893 29200 17280 29202
rect 12893 29144 12898 29200
rect 12954 29144 15750 29200
rect 15806 29144 17280 29200
rect 12893 29142 17280 29144
rect 12893 29139 12959 29142
rect 15745 29139 15811 29142
rect 13353 29066 13419 29069
rect 14457 29066 14523 29069
rect 12390 29006 13232 29066
rect 9508 29004 9514 29006
rect 9949 29003 10015 29006
rect 13172 28930 13232 29006
rect 13353 29064 14523 29066
rect 13353 29008 13358 29064
rect 13414 29008 14462 29064
rect 14518 29008 14523 29064
rect 13353 29006 14523 29008
rect 13353 29003 13419 29006
rect 14457 29003 14523 29006
rect 15694 29004 15700 29068
rect 15764 29066 15770 29068
rect 16205 29066 16271 29069
rect 15764 29064 16271 29066
rect 15764 29008 16210 29064
rect 16266 29008 16271 29064
rect 15764 29006 16271 29008
rect 17220 29066 17280 29142
rect 19241 29200 19932 29202
rect 19241 29144 19246 29200
rect 19302 29144 19932 29200
rect 19241 29142 19932 29144
rect 19241 29139 19307 29142
rect 19926 29140 19932 29142
rect 19996 29202 20002 29204
rect 21541 29202 21607 29205
rect 19996 29200 21607 29202
rect 19996 29144 21546 29200
rect 21602 29144 21607 29200
rect 19996 29142 21607 29144
rect 19996 29140 20002 29142
rect 21541 29139 21607 29142
rect 21950 29140 21956 29204
rect 22020 29202 22026 29204
rect 23657 29202 23723 29205
rect 22020 29200 23723 29202
rect 22020 29144 23662 29200
rect 23718 29144 23723 29200
rect 22020 29142 23723 29144
rect 22020 29140 22026 29142
rect 23657 29139 23723 29142
rect 24209 29202 24275 29205
rect 24761 29202 24827 29205
rect 24209 29200 24827 29202
rect 24209 29144 24214 29200
rect 24270 29144 24766 29200
rect 24822 29144 24827 29200
rect 24209 29142 24827 29144
rect 24209 29139 24275 29142
rect 24761 29139 24827 29142
rect 24945 29202 25011 29205
rect 26550 29202 26556 29204
rect 24945 29200 26556 29202
rect 24945 29144 24950 29200
rect 25006 29144 26556 29200
rect 24945 29142 26556 29144
rect 24945 29139 25011 29142
rect 26550 29140 26556 29142
rect 26620 29140 26626 29204
rect 26918 29140 26924 29204
rect 26988 29202 26994 29204
rect 32078 29202 32138 29278
rect 32673 29275 32739 29278
rect 26988 29142 32138 29202
rect 26988 29140 26994 29142
rect 22737 29066 22803 29069
rect 22921 29066 22987 29069
rect 17220 29064 22987 29066
rect 17220 29008 22742 29064
rect 22798 29008 22926 29064
rect 22982 29008 22987 29064
rect 17220 29006 22987 29008
rect 15764 29004 15770 29006
rect 16205 29003 16271 29006
rect 22737 29003 22803 29006
rect 22921 29003 22987 29006
rect 23105 29066 23171 29069
rect 23289 29066 23355 29069
rect 24301 29066 24367 29069
rect 23105 29064 23355 29066
rect 23105 29008 23110 29064
rect 23166 29008 23294 29064
rect 23350 29008 23355 29064
rect 23105 29006 23355 29008
rect 23105 29003 23171 29006
rect 23289 29003 23355 29006
rect 23568 29064 24367 29066
rect 23568 29008 24306 29064
rect 24362 29008 24367 29064
rect 23568 29006 24367 29008
rect 23568 28933 23628 29006
rect 24301 29003 24367 29006
rect 24894 29004 24900 29068
rect 24964 29066 24970 29068
rect 26509 29066 26575 29069
rect 24964 29064 26575 29066
rect 24964 29008 26514 29064
rect 26570 29008 26575 29064
rect 24964 29006 26575 29008
rect 24964 29004 24970 29006
rect 26509 29003 26575 29006
rect 26918 29004 26924 29068
rect 26988 29066 26994 29068
rect 27286 29066 27292 29068
rect 26988 29006 27292 29066
rect 26988 29004 26994 29006
rect 27286 29004 27292 29006
rect 27356 29004 27362 29068
rect 28809 29066 28875 29069
rect 27432 29064 28875 29066
rect 27432 29008 28814 29064
rect 28870 29008 28875 29064
rect 27432 29006 28875 29008
rect 18229 28930 18295 28933
rect 13172 28928 18295 28930
rect 13172 28872 18234 28928
rect 18290 28872 18295 28928
rect 13172 28870 18295 28872
rect 18229 28867 18295 28870
rect 18505 28930 18571 28933
rect 19241 28930 19307 28933
rect 18505 28928 19307 28930
rect 18505 28872 18510 28928
rect 18566 28872 19246 28928
rect 19302 28872 19307 28928
rect 18505 28870 19307 28872
rect 18505 28867 18571 28870
rect 19241 28867 19307 28870
rect 19425 28930 19491 28933
rect 19558 28930 19564 28932
rect 19425 28928 19564 28930
rect 19425 28872 19430 28928
rect 19486 28872 19564 28928
rect 19425 28870 19564 28872
rect 19425 28867 19491 28870
rect 19558 28868 19564 28870
rect 19628 28868 19634 28932
rect 20621 28930 20687 28933
rect 22553 28930 22619 28933
rect 20621 28928 22619 28930
rect 20621 28872 20626 28928
rect 20682 28872 22558 28928
rect 22614 28872 22619 28928
rect 20621 28870 22619 28872
rect 20621 28867 20687 28870
rect 22553 28867 22619 28870
rect 22686 28868 22692 28932
rect 22756 28930 22762 28932
rect 23105 28930 23171 28933
rect 22756 28928 23171 28930
rect 22756 28872 23110 28928
rect 23166 28872 23171 28928
rect 22756 28870 23171 28872
rect 22756 28868 22762 28870
rect 23105 28867 23171 28870
rect 23565 28928 23631 28933
rect 23565 28872 23570 28928
rect 23626 28872 23631 28928
rect 23565 28867 23631 28872
rect 23933 28930 23999 28933
rect 26601 28930 26667 28933
rect 23933 28928 26667 28930
rect 23933 28872 23938 28928
rect 23994 28872 26606 28928
rect 26662 28872 26667 28928
rect 23933 28870 26667 28872
rect 23933 28867 23999 28870
rect 26601 28867 26667 28870
rect 26785 28930 26851 28933
rect 27432 28930 27492 29006
rect 28809 29003 28875 29006
rect 29821 29066 29887 29069
rect 31518 29066 31524 29068
rect 29821 29064 31524 29066
rect 29821 29008 29826 29064
rect 29882 29008 31524 29064
rect 29821 29006 31524 29008
rect 29821 29003 29887 29006
rect 31518 29004 31524 29006
rect 31588 29004 31594 29068
rect 32206 28976 33006 29096
rect 26785 28928 27492 28930
rect 26785 28872 26790 28928
rect 26846 28872 27492 28928
rect 26785 28870 27492 28872
rect 28257 28930 28323 28933
rect 28257 28928 28642 28930
rect 28257 28872 28262 28928
rect 28318 28872 28642 28928
rect 28257 28870 28642 28872
rect 26785 28867 26851 28870
rect 28257 28867 28323 28870
rect 4787 28864 5103 28865
rect 4787 28800 4793 28864
rect 4857 28800 4873 28864
rect 4937 28800 4953 28864
rect 5017 28800 5033 28864
rect 5097 28800 5103 28864
rect 4787 28799 5103 28800
rect 12469 28864 12785 28865
rect 12469 28800 12475 28864
rect 12539 28800 12555 28864
rect 12619 28800 12635 28864
rect 12699 28800 12715 28864
rect 12779 28800 12785 28864
rect 12469 28799 12785 28800
rect 20151 28864 20467 28865
rect 20151 28800 20157 28864
rect 20221 28800 20237 28864
rect 20301 28800 20317 28864
rect 20381 28800 20397 28864
rect 20461 28800 20467 28864
rect 20151 28799 20467 28800
rect 27833 28864 28149 28865
rect 27833 28800 27839 28864
rect 27903 28800 27919 28864
rect 27983 28800 27999 28864
rect 28063 28800 28079 28864
rect 28143 28800 28149 28864
rect 27833 28799 28149 28800
rect 13813 28794 13879 28797
rect 19977 28794 20043 28797
rect 13813 28792 20043 28794
rect 13813 28736 13818 28792
rect 13874 28736 19982 28792
rect 20038 28736 20043 28792
rect 13813 28734 20043 28736
rect 13813 28731 13879 28734
rect 19977 28731 20043 28734
rect 20713 28794 20779 28797
rect 20846 28794 20852 28796
rect 20713 28792 20852 28794
rect 20713 28736 20718 28792
rect 20774 28736 20852 28792
rect 20713 28734 20852 28736
rect 20713 28731 20779 28734
rect 20846 28732 20852 28734
rect 20916 28794 20922 28796
rect 21817 28794 21883 28797
rect 20916 28792 21883 28794
rect 20916 28736 21822 28792
rect 21878 28736 21883 28792
rect 20916 28734 21883 28736
rect 20916 28732 20922 28734
rect 21817 28731 21883 28734
rect 22001 28794 22067 28797
rect 26601 28794 26667 28797
rect 22001 28792 26667 28794
rect 22001 28736 22006 28792
rect 22062 28736 26606 28792
rect 26662 28736 26667 28792
rect 22001 28734 26667 28736
rect 22001 28731 22067 28734
rect 26601 28731 26667 28734
rect 26785 28794 26851 28797
rect 27521 28794 27587 28797
rect 26785 28792 27587 28794
rect 26785 28736 26790 28792
rect 26846 28736 27526 28792
rect 27582 28736 27587 28792
rect 28441 28792 28507 28797
rect 28441 28760 28446 28792
rect 26785 28734 27587 28736
rect 26785 28731 26851 28734
rect 27521 28731 27587 28734
rect 28352 28736 28446 28760
rect 28502 28736 28507 28792
rect 28352 28731 28507 28736
rect 28582 28794 28642 28870
rect 28758 28868 28764 28932
rect 28828 28930 28834 28932
rect 28901 28930 28967 28933
rect 28828 28928 28967 28930
rect 28828 28872 28906 28928
rect 28962 28872 28967 28928
rect 28828 28870 28967 28872
rect 28828 28868 28834 28870
rect 28901 28867 28967 28870
rect 32438 28794 32444 28796
rect 28582 28734 32444 28794
rect 32438 28732 32444 28734
rect 32508 28732 32514 28796
rect 28352 28700 28504 28731
rect 15469 28658 15535 28661
rect 18781 28658 18847 28661
rect 15469 28656 18847 28658
rect 15469 28600 15474 28656
rect 15530 28600 18786 28656
rect 18842 28600 18847 28656
rect 15469 28598 18847 28600
rect 15469 28595 15535 28598
rect 18781 28595 18847 28598
rect 19006 28596 19012 28660
rect 19076 28658 19082 28660
rect 19333 28658 19399 28661
rect 19076 28656 19399 28658
rect 19076 28600 19338 28656
rect 19394 28600 19399 28656
rect 19076 28598 19399 28600
rect 19076 28596 19082 28598
rect 19333 28595 19399 28598
rect 19742 28596 19748 28660
rect 19812 28658 19818 28660
rect 20345 28658 20411 28661
rect 25773 28658 25839 28661
rect 19812 28656 20411 28658
rect 19812 28600 20350 28656
rect 20406 28600 20411 28656
rect 19812 28598 20411 28600
rect 19812 28596 19818 28598
rect 20345 28595 20411 28598
rect 20532 28656 25839 28658
rect 20532 28600 25778 28656
rect 25834 28600 25839 28656
rect 20532 28598 25839 28600
rect 0 28522 800 28552
rect 1577 28522 1643 28525
rect 0 28520 1643 28522
rect 0 28464 1582 28520
rect 1638 28464 1643 28520
rect 0 28462 1643 28464
rect 0 28432 800 28462
rect 1577 28459 1643 28462
rect 16982 28460 16988 28524
rect 17052 28522 17058 28524
rect 20532 28522 20592 28598
rect 25773 28595 25839 28598
rect 25998 28596 26004 28660
rect 26068 28658 26074 28660
rect 28352 28658 28412 28700
rect 26068 28598 28412 28658
rect 28901 28658 28967 28661
rect 29453 28660 29519 28661
rect 29310 28658 29316 28660
rect 28901 28656 29316 28658
rect 28901 28600 28906 28656
rect 28962 28600 29316 28656
rect 28901 28598 29316 28600
rect 26068 28596 26074 28598
rect 28901 28595 28967 28598
rect 29310 28596 29316 28598
rect 29380 28596 29386 28660
rect 29453 28656 29500 28660
rect 29564 28658 29570 28660
rect 29453 28600 29458 28656
rect 29453 28596 29500 28600
rect 29564 28598 29610 28658
rect 29564 28596 29570 28598
rect 29453 28595 29519 28596
rect 17052 28462 20592 28522
rect 20713 28522 20779 28525
rect 20897 28522 20963 28525
rect 21950 28522 21956 28524
rect 20713 28520 21956 28522
rect 20713 28464 20718 28520
rect 20774 28464 20902 28520
rect 20958 28464 21956 28520
rect 20713 28462 21956 28464
rect 17052 28460 17058 28462
rect 20713 28459 20779 28462
rect 20897 28459 20963 28462
rect 21950 28460 21956 28462
rect 22020 28460 22026 28524
rect 22870 28460 22876 28524
rect 22940 28522 22946 28524
rect 30373 28522 30439 28525
rect 22940 28520 30439 28522
rect 22940 28464 30378 28520
rect 30434 28464 30439 28520
rect 22940 28462 30439 28464
rect 22940 28460 22946 28462
rect 30373 28459 30439 28462
rect 30649 28522 30715 28525
rect 30649 28520 32138 28522
rect 30649 28464 30654 28520
rect 30710 28464 32138 28520
rect 30649 28462 32138 28464
rect 30649 28459 30715 28462
rect 16849 28386 16915 28389
rect 19425 28386 19491 28389
rect 23565 28386 23631 28389
rect 26233 28388 26299 28389
rect 16849 28384 23631 28386
rect 16849 28328 16854 28384
rect 16910 28328 19430 28384
rect 19486 28328 23570 28384
rect 23626 28328 23631 28384
rect 16849 28326 23631 28328
rect 16849 28323 16915 28326
rect 19425 28323 19491 28326
rect 23565 28323 23631 28326
rect 24526 28324 24532 28388
rect 24596 28386 24602 28388
rect 24894 28386 24900 28388
rect 24596 28326 24900 28386
rect 24596 28324 24602 28326
rect 24894 28324 24900 28326
rect 24964 28324 24970 28388
rect 25078 28324 25084 28388
rect 25148 28386 25154 28388
rect 25998 28386 26004 28388
rect 25148 28326 26004 28386
rect 25148 28324 25154 28326
rect 25998 28324 26004 28326
rect 26068 28324 26074 28388
rect 26182 28324 26188 28388
rect 26252 28386 26299 28388
rect 26601 28386 26667 28389
rect 28206 28386 28212 28388
rect 26252 28384 26344 28386
rect 26294 28328 26344 28384
rect 26252 28326 26344 28328
rect 26601 28384 28212 28386
rect 26601 28328 26606 28384
rect 26662 28328 28212 28384
rect 26601 28326 28212 28328
rect 26252 28324 26299 28326
rect 26233 28323 26299 28324
rect 26601 28323 26667 28326
rect 28206 28324 28212 28326
rect 28276 28324 28282 28388
rect 28441 28386 28507 28389
rect 28574 28386 28580 28388
rect 28441 28384 28580 28386
rect 28441 28328 28446 28384
rect 28502 28328 28580 28384
rect 28441 28326 28580 28328
rect 28441 28323 28507 28326
rect 28574 28324 28580 28326
rect 28644 28324 28650 28388
rect 29269 28386 29335 28389
rect 29494 28386 29500 28388
rect 29269 28384 29500 28386
rect 29269 28328 29274 28384
rect 29330 28328 29500 28384
rect 29269 28326 29500 28328
rect 29269 28323 29335 28326
rect 29494 28324 29500 28326
rect 29564 28324 29570 28388
rect 30005 28386 30071 28389
rect 31334 28386 31340 28388
rect 30005 28384 31340 28386
rect 30005 28328 30010 28384
rect 30066 28328 31340 28384
rect 30005 28326 31340 28328
rect 30005 28323 30071 28326
rect 31334 28324 31340 28326
rect 31404 28324 31410 28388
rect 32078 28386 32138 28462
rect 32206 28386 33006 28416
rect 32078 28326 33006 28386
rect 8628 28320 8944 28321
rect 8628 28256 8634 28320
rect 8698 28256 8714 28320
rect 8778 28256 8794 28320
rect 8858 28256 8874 28320
rect 8938 28256 8944 28320
rect 8628 28255 8944 28256
rect 16310 28320 16626 28321
rect 16310 28256 16316 28320
rect 16380 28256 16396 28320
rect 16460 28256 16476 28320
rect 16540 28256 16556 28320
rect 16620 28256 16626 28320
rect 16310 28255 16626 28256
rect 23992 28320 24308 28321
rect 23992 28256 23998 28320
rect 24062 28256 24078 28320
rect 24142 28256 24158 28320
rect 24222 28256 24238 28320
rect 24302 28256 24308 28320
rect 23992 28255 24308 28256
rect 31674 28320 31990 28321
rect 31674 28256 31680 28320
rect 31744 28256 31760 28320
rect 31824 28256 31840 28320
rect 31904 28256 31920 28320
rect 31984 28256 31990 28320
rect 32206 28296 33006 28326
rect 31674 28255 31990 28256
rect 14774 28188 14780 28252
rect 14844 28250 14850 28252
rect 15929 28250 15995 28253
rect 18597 28252 18663 28253
rect 14844 28248 15995 28250
rect 14844 28192 15934 28248
rect 15990 28192 15995 28248
rect 14844 28190 15995 28192
rect 14844 28188 14850 28190
rect 15929 28187 15995 28190
rect 16798 28188 16804 28252
rect 16868 28250 16874 28252
rect 18454 28250 18460 28252
rect 16868 28190 18460 28250
rect 16868 28188 16874 28190
rect 18454 28188 18460 28190
rect 18524 28188 18530 28252
rect 18597 28248 18644 28252
rect 18708 28250 18714 28252
rect 18965 28250 19031 28253
rect 22185 28250 22251 28253
rect 18597 28192 18602 28248
rect 18597 28188 18644 28192
rect 18708 28190 18754 28250
rect 18965 28248 22251 28250
rect 18965 28192 18970 28248
rect 19026 28192 22190 28248
rect 22246 28192 22251 28248
rect 18965 28190 22251 28192
rect 18708 28188 18714 28190
rect 18597 28187 18663 28188
rect 18965 28187 19031 28190
rect 22185 28187 22251 28190
rect 22318 28188 22324 28252
rect 22388 28250 22394 28252
rect 22553 28250 22619 28253
rect 23657 28252 23723 28253
rect 22388 28248 22619 28250
rect 22388 28192 22558 28248
rect 22614 28192 22619 28248
rect 22388 28190 22619 28192
rect 22388 28188 22394 28190
rect 22553 28187 22619 28190
rect 22686 28188 22692 28252
rect 22756 28250 22762 28252
rect 23606 28250 23612 28252
rect 22756 28190 23490 28250
rect 23566 28190 23612 28250
rect 23676 28248 23723 28252
rect 23718 28192 23723 28248
rect 22756 28188 22762 28190
rect 14549 28116 14615 28117
rect 14549 28112 14596 28116
rect 14660 28114 14666 28116
rect 14549 28056 14554 28112
rect 14549 28052 14596 28056
rect 14660 28054 14706 28114
rect 14660 28052 14666 28054
rect 15878 28052 15884 28116
rect 15948 28114 15954 28116
rect 22921 28114 22987 28117
rect 15948 28112 22987 28114
rect 15948 28056 22926 28112
rect 22982 28056 22987 28112
rect 15948 28054 22987 28056
rect 23430 28114 23490 28190
rect 23606 28188 23612 28190
rect 23676 28188 23723 28192
rect 23657 28187 23723 28188
rect 24577 28250 24643 28253
rect 25814 28250 25820 28252
rect 24577 28248 25820 28250
rect 24577 28192 24582 28248
rect 24638 28192 25820 28248
rect 24577 28190 25820 28192
rect 24577 28187 24643 28190
rect 25814 28188 25820 28190
rect 25884 28188 25890 28252
rect 25998 28188 26004 28252
rect 26068 28250 26074 28252
rect 26417 28250 26483 28253
rect 26068 28248 26483 28250
rect 26068 28192 26422 28248
rect 26478 28192 26483 28248
rect 26068 28190 26483 28192
rect 26068 28188 26074 28190
rect 26417 28187 26483 28190
rect 26785 28250 26851 28253
rect 29310 28250 29316 28252
rect 26785 28248 29316 28250
rect 26785 28192 26790 28248
rect 26846 28192 29316 28248
rect 26785 28190 29316 28192
rect 26785 28187 26851 28190
rect 29310 28188 29316 28190
rect 29380 28188 29386 28252
rect 23430 28054 24364 28114
rect 15948 28052 15954 28054
rect 14549 28051 14615 28052
rect 22921 28051 22987 28054
rect 24304 27981 24364 28054
rect 25630 28052 25636 28116
rect 25700 28114 25706 28116
rect 29821 28114 29887 28117
rect 25700 28112 29887 28114
rect 25700 28056 29826 28112
rect 29882 28056 29887 28112
rect 25700 28054 29887 28056
rect 25700 28052 25706 28054
rect 29821 28051 29887 28054
rect 10317 27978 10383 27981
rect 13302 27978 13308 27980
rect 10317 27976 13308 27978
rect 10317 27920 10322 27976
rect 10378 27920 13308 27976
rect 10317 27918 13308 27920
rect 10317 27915 10383 27918
rect 13302 27916 13308 27918
rect 13372 27978 13378 27980
rect 18965 27978 19031 27981
rect 13372 27976 19031 27978
rect 13372 27920 18970 27976
rect 19026 27920 19031 27976
rect 13372 27918 19031 27920
rect 13372 27916 13378 27918
rect 18965 27915 19031 27918
rect 19149 27978 19215 27981
rect 20989 27978 21055 27981
rect 22093 27978 22159 27981
rect 23565 27978 23631 27981
rect 19149 27976 23631 27978
rect 19149 27920 19154 27976
rect 19210 27920 20994 27976
rect 21050 27920 22098 27976
rect 22154 27920 23570 27976
rect 23626 27920 23631 27976
rect 19149 27918 23631 27920
rect 19149 27915 19215 27918
rect 20989 27915 21055 27918
rect 22093 27915 22159 27918
rect 23565 27915 23631 27918
rect 24301 27978 24367 27981
rect 26417 27978 26483 27981
rect 24301 27976 26483 27978
rect 24301 27920 24306 27976
rect 24362 27920 26422 27976
rect 26478 27920 26483 27976
rect 24301 27918 26483 27920
rect 24301 27915 24367 27918
rect 26417 27915 26483 27918
rect 26785 27978 26851 27981
rect 28574 27978 28580 27980
rect 26785 27976 28580 27978
rect 26785 27920 26790 27976
rect 26846 27920 28580 27976
rect 26785 27918 28580 27920
rect 26785 27915 26851 27918
rect 28574 27916 28580 27918
rect 28644 27916 28650 27980
rect 29453 27978 29519 27981
rect 32070 27978 32076 27980
rect 29453 27976 32076 27978
rect 29453 27920 29458 27976
rect 29514 27920 32076 27976
rect 29453 27918 32076 27920
rect 29453 27915 29519 27918
rect 32070 27916 32076 27918
rect 32140 27916 32146 27980
rect 13670 27780 13676 27844
rect 13740 27842 13746 27844
rect 18413 27842 18479 27845
rect 13740 27840 18479 27842
rect 13740 27784 18418 27840
rect 18474 27784 18479 27840
rect 13740 27782 18479 27784
rect 13740 27780 13746 27782
rect 18413 27779 18479 27782
rect 18597 27842 18663 27845
rect 19609 27842 19675 27845
rect 18597 27840 19675 27842
rect 18597 27784 18602 27840
rect 18658 27784 19614 27840
rect 19670 27784 19675 27840
rect 18597 27782 19675 27784
rect 18597 27779 18663 27782
rect 19609 27779 19675 27782
rect 20662 27780 20668 27844
rect 20732 27842 20738 27844
rect 20805 27842 20871 27845
rect 20732 27840 20871 27842
rect 20732 27784 20810 27840
rect 20866 27784 20871 27840
rect 20732 27782 20871 27784
rect 20732 27780 20738 27782
rect 20805 27779 20871 27782
rect 21541 27844 21607 27845
rect 21817 27844 21883 27845
rect 21541 27840 21588 27844
rect 21652 27842 21658 27844
rect 21541 27784 21546 27840
rect 21541 27780 21588 27784
rect 21652 27782 21698 27842
rect 21652 27780 21658 27782
rect 21766 27780 21772 27844
rect 21836 27842 21883 27844
rect 21836 27840 21928 27842
rect 21878 27784 21928 27840
rect 21836 27782 21928 27784
rect 21836 27780 21883 27782
rect 22134 27780 22140 27844
rect 22204 27842 22210 27844
rect 22553 27842 22619 27845
rect 22204 27840 22619 27842
rect 22204 27784 22558 27840
rect 22614 27784 22619 27840
rect 22204 27782 22619 27784
rect 22204 27780 22210 27782
rect 21541 27779 21607 27780
rect 21817 27779 21883 27780
rect 22553 27779 22619 27782
rect 22686 27780 22692 27844
rect 22756 27842 22762 27844
rect 24117 27842 24183 27845
rect 22756 27840 24183 27842
rect 22756 27784 24122 27840
rect 24178 27784 24183 27840
rect 22756 27782 24183 27784
rect 22756 27780 22762 27782
rect 24117 27779 24183 27782
rect 24669 27842 24735 27845
rect 25221 27844 25287 27845
rect 24894 27842 24900 27844
rect 24669 27840 24900 27842
rect 24669 27784 24674 27840
rect 24730 27784 24900 27840
rect 24669 27782 24900 27784
rect 24669 27779 24735 27782
rect 24894 27780 24900 27782
rect 24964 27780 24970 27844
rect 25221 27842 25268 27844
rect 25176 27840 25268 27842
rect 25176 27784 25226 27840
rect 25176 27782 25268 27784
rect 25221 27780 25268 27782
rect 25332 27780 25338 27844
rect 25405 27842 25471 27845
rect 25589 27842 25655 27845
rect 25405 27840 25655 27842
rect 25405 27784 25410 27840
rect 25466 27784 25594 27840
rect 25650 27784 25655 27840
rect 25405 27782 25655 27784
rect 25221 27779 25287 27780
rect 25405 27779 25471 27782
rect 25589 27779 25655 27782
rect 25773 27842 25839 27845
rect 26141 27842 26207 27845
rect 25773 27840 26207 27842
rect 25773 27784 25778 27840
rect 25834 27784 26146 27840
rect 26202 27784 26207 27840
rect 25773 27782 26207 27784
rect 25773 27779 25839 27782
rect 26141 27779 26207 27782
rect 26366 27780 26372 27844
rect 26436 27842 26442 27844
rect 26509 27842 26575 27845
rect 26436 27840 26575 27842
rect 26436 27784 26514 27840
rect 26570 27784 26575 27840
rect 26436 27782 26575 27784
rect 26436 27780 26442 27782
rect 26509 27779 26575 27782
rect 26785 27842 26851 27845
rect 27705 27844 27771 27845
rect 26918 27842 26924 27844
rect 26785 27840 26924 27842
rect 26785 27784 26790 27840
rect 26846 27784 26924 27840
rect 26785 27782 26924 27784
rect 26785 27779 26851 27782
rect 26918 27780 26924 27782
rect 26988 27780 26994 27844
rect 27654 27842 27660 27844
rect 27614 27782 27660 27842
rect 27724 27840 27771 27844
rect 27766 27784 27771 27840
rect 27654 27780 27660 27782
rect 27724 27780 27771 27784
rect 27705 27779 27771 27780
rect 28253 27842 28319 27845
rect 28625 27842 28691 27845
rect 28253 27840 28691 27842
rect 28253 27784 28258 27840
rect 28314 27784 28630 27840
rect 28686 27784 28691 27840
rect 28253 27782 28691 27784
rect 28253 27779 28319 27782
rect 28625 27779 28691 27782
rect 29269 27842 29335 27845
rect 29862 27842 29868 27844
rect 29269 27840 29868 27842
rect 29269 27784 29274 27840
rect 29330 27784 29868 27840
rect 29269 27782 29868 27784
rect 29269 27779 29335 27782
rect 29862 27780 29868 27782
rect 29932 27780 29938 27844
rect 4787 27776 5103 27777
rect 0 27706 800 27736
rect 4787 27712 4793 27776
rect 4857 27712 4873 27776
rect 4937 27712 4953 27776
rect 5017 27712 5033 27776
rect 5097 27712 5103 27776
rect 4787 27711 5103 27712
rect 12469 27776 12785 27777
rect 12469 27712 12475 27776
rect 12539 27712 12555 27776
rect 12619 27712 12635 27776
rect 12699 27712 12715 27776
rect 12779 27712 12785 27776
rect 12469 27711 12785 27712
rect 20151 27776 20467 27777
rect 20151 27712 20157 27776
rect 20221 27712 20237 27776
rect 20301 27712 20317 27776
rect 20381 27712 20397 27776
rect 20461 27712 20467 27776
rect 20151 27711 20467 27712
rect 27833 27776 28149 27777
rect 27833 27712 27839 27776
rect 27903 27712 27919 27776
rect 27983 27712 27999 27776
rect 28063 27712 28079 27776
rect 28143 27712 28149 27776
rect 27833 27711 28149 27712
rect 1577 27706 1643 27709
rect 18873 27706 18939 27709
rect 0 27704 1643 27706
rect 0 27648 1582 27704
rect 1638 27648 1643 27704
rect 0 27646 1643 27648
rect 0 27616 800 27646
rect 1577 27643 1643 27646
rect 12896 27704 18939 27706
rect 12896 27648 18878 27704
rect 18934 27648 18939 27704
rect 12896 27646 18939 27648
rect 12014 27508 12020 27572
rect 12084 27570 12090 27572
rect 12896 27570 12956 27646
rect 18873 27643 18939 27646
rect 19190 27644 19196 27708
rect 19260 27706 19266 27708
rect 19793 27706 19859 27709
rect 19260 27704 19859 27706
rect 19260 27648 19798 27704
rect 19854 27648 19859 27704
rect 19260 27646 19859 27648
rect 19260 27644 19266 27646
rect 19793 27643 19859 27646
rect 20846 27644 20852 27708
rect 20916 27706 20922 27708
rect 21633 27706 21699 27709
rect 20916 27704 21699 27706
rect 20916 27648 21638 27704
rect 21694 27648 21699 27704
rect 20916 27646 21699 27648
rect 20916 27644 20922 27646
rect 21633 27643 21699 27646
rect 22134 27644 22140 27708
rect 22204 27706 22210 27708
rect 22502 27706 22508 27708
rect 22204 27646 22508 27706
rect 22204 27644 22210 27646
rect 22502 27644 22508 27646
rect 22572 27644 22578 27708
rect 24577 27706 24643 27709
rect 22648 27704 24643 27706
rect 22648 27648 24582 27704
rect 24638 27648 24643 27704
rect 22648 27646 24643 27648
rect 12084 27510 12956 27570
rect 15377 27570 15443 27573
rect 15745 27570 15811 27573
rect 15377 27568 15811 27570
rect 15377 27512 15382 27568
rect 15438 27512 15750 27568
rect 15806 27512 15811 27568
rect 15377 27510 15811 27512
rect 12084 27508 12090 27510
rect 15377 27507 15443 27510
rect 15745 27507 15811 27510
rect 15929 27570 15995 27573
rect 16062 27570 16068 27572
rect 15929 27568 16068 27570
rect 15929 27512 15934 27568
rect 15990 27512 16068 27568
rect 15929 27510 16068 27512
rect 15929 27507 15995 27510
rect 16062 27508 16068 27510
rect 16132 27508 16138 27572
rect 16205 27570 16271 27573
rect 17493 27570 17559 27573
rect 16205 27568 17559 27570
rect 16205 27512 16210 27568
rect 16266 27512 17498 27568
rect 17554 27512 17559 27568
rect 16205 27510 17559 27512
rect 16205 27507 16271 27510
rect 17493 27507 17559 27510
rect 17861 27570 17927 27573
rect 18045 27570 18111 27573
rect 17861 27568 18111 27570
rect 17861 27512 17866 27568
rect 17922 27512 18050 27568
rect 18106 27512 18111 27568
rect 17861 27510 18111 27512
rect 17861 27507 17927 27510
rect 18045 27507 18111 27510
rect 18454 27508 18460 27572
rect 18524 27570 18530 27572
rect 19057 27570 19123 27573
rect 18524 27568 19123 27570
rect 18524 27512 19062 27568
rect 19118 27512 19123 27568
rect 18524 27510 19123 27512
rect 18524 27508 18530 27510
rect 19057 27507 19123 27510
rect 19190 27508 19196 27572
rect 19260 27570 19266 27572
rect 20253 27570 20319 27573
rect 21081 27570 21147 27573
rect 19260 27568 21147 27570
rect 19260 27512 20258 27568
rect 20314 27512 21086 27568
rect 21142 27512 21147 27568
rect 19260 27510 21147 27512
rect 19260 27508 19266 27510
rect 20253 27507 20319 27510
rect 21081 27507 21147 27510
rect 21214 27508 21220 27572
rect 21284 27570 21290 27572
rect 21357 27570 21423 27573
rect 21284 27568 21423 27570
rect 21284 27512 21362 27568
rect 21418 27512 21423 27568
rect 21284 27510 21423 27512
rect 21284 27508 21290 27510
rect 21357 27507 21423 27510
rect 21817 27570 21883 27573
rect 22001 27570 22067 27573
rect 22461 27572 22527 27573
rect 22461 27570 22508 27572
rect 21817 27568 22067 27570
rect 21817 27512 21822 27568
rect 21878 27512 22006 27568
rect 22062 27512 22067 27568
rect 21817 27510 22067 27512
rect 22416 27568 22508 27570
rect 22416 27512 22466 27568
rect 22416 27510 22508 27512
rect 21817 27507 21883 27510
rect 22001 27507 22067 27510
rect 22461 27508 22508 27510
rect 22572 27508 22578 27572
rect 22461 27507 22527 27508
rect 8017 27434 8083 27437
rect 14181 27434 14247 27437
rect 8017 27432 14247 27434
rect 8017 27376 8022 27432
rect 8078 27376 14186 27432
rect 14242 27376 14247 27432
rect 8017 27374 14247 27376
rect 8017 27371 8083 27374
rect 14181 27371 14247 27374
rect 14917 27434 14983 27437
rect 21081 27434 21147 27437
rect 14917 27432 21147 27434
rect 14917 27376 14922 27432
rect 14978 27376 21086 27432
rect 21142 27376 21147 27432
rect 14917 27374 21147 27376
rect 14917 27371 14983 27374
rect 21081 27371 21147 27374
rect 21214 27372 21220 27436
rect 21284 27434 21290 27436
rect 22648 27434 22708 27646
rect 24577 27643 24643 27646
rect 25313 27706 25379 27709
rect 26969 27706 27035 27709
rect 27613 27708 27679 27709
rect 27613 27706 27660 27708
rect 25313 27704 27035 27706
rect 25313 27648 25318 27704
rect 25374 27648 26974 27704
rect 27030 27648 27035 27704
rect 25313 27646 27035 27648
rect 27568 27704 27660 27706
rect 27568 27648 27618 27704
rect 27568 27646 27660 27648
rect 25313 27643 25379 27646
rect 26969 27643 27035 27646
rect 27613 27644 27660 27646
rect 27724 27644 27730 27708
rect 28252 27644 28258 27708
rect 28322 27706 28328 27708
rect 29085 27706 29151 27709
rect 28322 27704 29151 27706
rect 28322 27648 29090 27704
rect 29146 27648 29151 27704
rect 28322 27646 29151 27648
rect 28322 27644 28328 27646
rect 27613 27643 27679 27644
rect 29085 27643 29151 27646
rect 29269 27706 29335 27709
rect 29494 27706 29500 27708
rect 29269 27704 29500 27706
rect 29269 27648 29274 27704
rect 29330 27648 29500 27704
rect 29269 27646 29500 27648
rect 29269 27643 29335 27646
rect 29494 27644 29500 27646
rect 29564 27644 29570 27708
rect 29821 27706 29887 27709
rect 30649 27706 30715 27709
rect 29821 27704 30715 27706
rect 29821 27648 29826 27704
rect 29882 27648 30654 27704
rect 30710 27648 30715 27704
rect 29821 27646 30715 27648
rect 29821 27643 29887 27646
rect 30649 27643 30715 27646
rect 31201 27706 31267 27709
rect 32206 27706 33006 27736
rect 31201 27704 33006 27706
rect 31201 27648 31206 27704
rect 31262 27648 33006 27704
rect 31201 27646 33006 27648
rect 31201 27643 31267 27646
rect 32206 27616 33006 27646
rect 22829 27570 22895 27573
rect 23013 27570 23079 27573
rect 23197 27572 23263 27573
rect 23381 27572 23447 27573
rect 23197 27570 23244 27572
rect 22829 27568 23079 27570
rect 22829 27512 22834 27568
rect 22890 27512 23018 27568
rect 23074 27512 23079 27568
rect 22829 27510 23079 27512
rect 23152 27568 23244 27570
rect 23152 27512 23202 27568
rect 23152 27510 23244 27512
rect 22829 27507 22895 27510
rect 23013 27507 23079 27510
rect 23197 27508 23244 27510
rect 23308 27508 23314 27572
rect 23381 27568 23428 27572
rect 23492 27570 23498 27572
rect 23381 27512 23386 27568
rect 23381 27508 23428 27512
rect 23492 27510 23538 27570
rect 23492 27508 23498 27510
rect 23606 27508 23612 27572
rect 23676 27570 23682 27572
rect 24025 27570 24091 27573
rect 23676 27568 24091 27570
rect 23676 27512 24030 27568
rect 24086 27512 24091 27568
rect 23676 27510 24091 27512
rect 23676 27508 23682 27510
rect 23197 27507 23263 27508
rect 23381 27507 23447 27508
rect 24025 27507 24091 27510
rect 24710 27508 24716 27572
rect 24780 27570 24786 27572
rect 26233 27570 26299 27573
rect 24780 27510 25284 27570
rect 24780 27508 24786 27510
rect 21284 27374 22708 27434
rect 22921 27434 22987 27437
rect 23289 27434 23355 27437
rect 22921 27432 23355 27434
rect 22921 27376 22926 27432
rect 22982 27376 23294 27432
rect 23350 27376 23355 27432
rect 22921 27374 23355 27376
rect 21284 27372 21290 27374
rect 22921 27371 22987 27374
rect 23289 27371 23355 27374
rect 23749 27434 23815 27437
rect 24117 27434 24183 27437
rect 24669 27434 24735 27437
rect 25078 27434 25084 27436
rect 23749 27432 23858 27434
rect 23749 27376 23754 27432
rect 23810 27376 23858 27432
rect 23749 27371 23858 27376
rect 24117 27432 24456 27434
rect 24117 27376 24122 27432
rect 24178 27376 24456 27432
rect 24117 27374 24456 27376
rect 24117 27371 24183 27374
rect 12249 27298 12315 27301
rect 15653 27298 15719 27301
rect 12249 27296 15719 27298
rect 12249 27240 12254 27296
rect 12310 27240 15658 27296
rect 15714 27240 15719 27296
rect 12249 27238 15719 27240
rect 12249 27235 12315 27238
rect 15653 27235 15719 27238
rect 17350 27236 17356 27300
rect 17420 27298 17426 27300
rect 22277 27298 22343 27301
rect 17420 27296 22343 27298
rect 17420 27240 22282 27296
rect 22338 27240 22343 27296
rect 17420 27238 22343 27240
rect 17420 27236 17426 27238
rect 22277 27235 22343 27238
rect 22461 27298 22527 27301
rect 22737 27298 22803 27301
rect 22461 27296 22803 27298
rect 22461 27240 22466 27296
rect 22522 27240 22742 27296
rect 22798 27240 22803 27296
rect 22461 27238 22803 27240
rect 22461 27235 22527 27238
rect 22737 27235 22803 27238
rect 23013 27298 23079 27301
rect 23657 27298 23723 27301
rect 23013 27296 23723 27298
rect 23013 27240 23018 27296
rect 23074 27240 23662 27296
rect 23718 27240 23723 27296
rect 23013 27238 23723 27240
rect 23013 27235 23079 27238
rect 23657 27235 23723 27238
rect 8628 27232 8944 27233
rect 8628 27168 8634 27232
rect 8698 27168 8714 27232
rect 8778 27168 8794 27232
rect 8858 27168 8874 27232
rect 8938 27168 8944 27232
rect 8628 27167 8944 27168
rect 16310 27232 16626 27233
rect 16310 27168 16316 27232
rect 16380 27168 16396 27232
rect 16460 27168 16476 27232
rect 16540 27168 16556 27232
rect 16620 27168 16626 27232
rect 16310 27167 16626 27168
rect 11513 27162 11579 27165
rect 16062 27162 16068 27164
rect 11513 27160 16068 27162
rect 11513 27104 11518 27160
rect 11574 27104 16068 27160
rect 11513 27102 16068 27104
rect 11513 27099 11579 27102
rect 16062 27100 16068 27102
rect 16132 27100 16138 27164
rect 18321 27162 18387 27165
rect 23606 27162 23612 27164
rect 18321 27160 23612 27162
rect 18321 27104 18326 27160
rect 18382 27104 23612 27160
rect 18321 27102 23612 27104
rect 18321 27099 18387 27102
rect 23606 27100 23612 27102
rect 23676 27100 23682 27164
rect 23798 27029 23858 27371
rect 24396 27298 24456 27374
rect 24669 27432 25084 27434
rect 24669 27376 24674 27432
rect 24730 27376 25084 27432
rect 24669 27374 25084 27376
rect 24669 27371 24735 27374
rect 25078 27372 25084 27374
rect 25148 27372 25154 27436
rect 25224 27434 25284 27510
rect 26233 27568 26848 27570
rect 26233 27512 26238 27568
rect 26294 27512 26848 27568
rect 26233 27510 26848 27512
rect 26233 27507 26299 27510
rect 26141 27434 26207 27437
rect 25224 27432 26207 27434
rect 25224 27376 26146 27432
rect 26202 27376 26207 27432
rect 25224 27374 26207 27376
rect 26788 27434 26848 27510
rect 26918 27508 26924 27572
rect 26988 27570 26994 27572
rect 27061 27570 27127 27573
rect 26988 27568 27127 27570
rect 26988 27512 27066 27568
rect 27122 27512 27127 27568
rect 26988 27510 27127 27512
rect 26988 27508 26994 27510
rect 27061 27507 27127 27510
rect 27889 27570 27955 27573
rect 31518 27570 31524 27572
rect 27889 27568 31524 27570
rect 27889 27512 27894 27568
rect 27950 27512 31524 27568
rect 27889 27510 31524 27512
rect 27889 27507 27955 27510
rect 31518 27508 31524 27510
rect 31588 27508 31594 27572
rect 30966 27434 30972 27436
rect 26788 27374 30972 27434
rect 26141 27371 26207 27374
rect 30966 27372 30972 27374
rect 31036 27372 31042 27436
rect 26417 27298 26483 27301
rect 24396 27296 26483 27298
rect 24396 27240 26422 27296
rect 26478 27240 26483 27296
rect 24396 27238 26483 27240
rect 26417 27235 26483 27238
rect 26734 27236 26740 27300
rect 26804 27298 26810 27300
rect 29545 27298 29611 27301
rect 26804 27296 29611 27298
rect 26804 27240 29550 27296
rect 29606 27240 29611 27296
rect 26804 27238 29611 27240
rect 26804 27236 26810 27238
rect 29545 27235 29611 27238
rect 29678 27236 29684 27300
rect 29748 27298 29754 27300
rect 29821 27298 29887 27301
rect 29748 27296 29887 27298
rect 29748 27240 29826 27296
rect 29882 27240 29887 27296
rect 29748 27238 29887 27240
rect 29748 27236 29754 27238
rect 29821 27235 29887 27238
rect 30046 27236 30052 27300
rect 30116 27298 30122 27300
rect 30465 27298 30531 27301
rect 30116 27296 30531 27298
rect 30116 27240 30470 27296
rect 30526 27240 30531 27296
rect 30116 27238 30531 27240
rect 30116 27236 30122 27238
rect 30465 27235 30531 27238
rect 23992 27232 24308 27233
rect 23992 27168 23998 27232
rect 24062 27168 24078 27232
rect 24142 27168 24158 27232
rect 24222 27168 24238 27232
rect 24302 27168 24308 27232
rect 23992 27167 24308 27168
rect 31674 27232 31990 27233
rect 31674 27168 31680 27232
rect 31744 27168 31760 27232
rect 31824 27168 31840 27232
rect 31904 27168 31920 27232
rect 31984 27168 31990 27232
rect 31674 27167 31990 27168
rect 25129 27164 25195 27165
rect 25078 27100 25084 27164
rect 25148 27162 25195 27164
rect 25957 27162 26023 27165
rect 26969 27162 27035 27165
rect 27521 27162 27587 27165
rect 25148 27160 25240 27162
rect 25190 27104 25240 27160
rect 25148 27102 25240 27104
rect 25957 27160 27587 27162
rect 25957 27104 25962 27160
rect 26018 27104 26974 27160
rect 27030 27104 27526 27160
rect 27582 27104 27587 27160
rect 25957 27102 27587 27104
rect 25148 27100 25195 27102
rect 25129 27099 25195 27100
rect 25957 27099 26023 27102
rect 26969 27099 27035 27102
rect 27521 27099 27587 27102
rect 27654 27100 27660 27164
rect 27724 27162 27730 27164
rect 27981 27162 28047 27165
rect 27724 27160 28047 27162
rect 27724 27104 27986 27160
rect 28042 27104 28047 27160
rect 27724 27102 28047 27104
rect 27724 27100 27730 27102
rect 27981 27099 28047 27102
rect 28165 27162 28231 27165
rect 28901 27162 28967 27165
rect 28165 27160 28967 27162
rect 28165 27104 28170 27160
rect 28226 27104 28906 27160
rect 28962 27104 28967 27160
rect 28165 27102 28967 27104
rect 28165 27099 28231 27102
rect 28901 27099 28967 27102
rect 30097 27162 30163 27165
rect 30230 27162 30236 27164
rect 30097 27160 30236 27162
rect 30097 27104 30102 27160
rect 30158 27104 30236 27160
rect 30097 27102 30236 27104
rect 30097 27099 30163 27102
rect 30230 27100 30236 27102
rect 30300 27100 30306 27164
rect 13813 27026 13879 27029
rect 13813 27024 17602 27026
rect 13813 26968 13818 27024
rect 13874 26968 17602 27024
rect 13813 26966 17602 26968
rect 13813 26963 13879 26966
rect 0 26800 800 26920
rect 5257 26890 5323 26893
rect 16573 26890 16639 26893
rect 5257 26888 16639 26890
rect 5257 26832 5262 26888
rect 5318 26832 16578 26888
rect 16634 26832 16639 26888
rect 5257 26830 16639 26832
rect 5257 26827 5323 26830
rect 16573 26827 16639 26830
rect 17166 26828 17172 26892
rect 17236 26890 17242 26892
rect 17401 26890 17467 26893
rect 17236 26888 17467 26890
rect 17236 26832 17406 26888
rect 17462 26832 17467 26888
rect 17236 26830 17467 26832
rect 17542 26890 17602 26966
rect 18454 26964 18460 27028
rect 18524 27026 18530 27028
rect 21173 27026 21239 27029
rect 22369 27026 22435 27029
rect 18524 27024 21239 27026
rect 18524 26968 21178 27024
rect 21234 26968 21239 27024
rect 18524 26966 21239 26968
rect 18524 26964 18530 26966
rect 21173 26963 21239 26966
rect 21406 27024 22435 27026
rect 21406 26968 22374 27024
rect 22430 26968 22435 27024
rect 21406 26966 22435 26968
rect 19793 26890 19859 26893
rect 21406 26890 21466 26966
rect 22369 26963 22435 26966
rect 22921 27026 22987 27029
rect 23238 27026 23244 27028
rect 22921 27024 23244 27026
rect 22921 26968 22926 27024
rect 22982 26968 23244 27024
rect 22921 26966 23244 26968
rect 22921 26963 22987 26966
rect 23238 26964 23244 26966
rect 23308 26964 23314 27028
rect 23749 27024 23858 27029
rect 23749 26968 23754 27024
rect 23810 26968 23858 27024
rect 23749 26966 23858 26968
rect 24025 27026 24091 27029
rect 24025 27024 29884 27026
rect 24025 26968 24030 27024
rect 24086 26968 29884 27024
rect 24025 26966 29884 26968
rect 23749 26963 23815 26966
rect 24025 26963 24091 26966
rect 24301 26890 24367 26893
rect 17542 26888 19859 26890
rect 17542 26832 19798 26888
rect 19854 26832 19859 26888
rect 17542 26830 19859 26832
rect 17236 26828 17242 26830
rect 17401 26827 17467 26830
rect 19793 26827 19859 26830
rect 19934 26830 21466 26890
rect 21544 26888 24367 26890
rect 21544 26832 24306 26888
rect 24362 26832 24367 26888
rect 21544 26830 24367 26832
rect 14181 26756 14247 26757
rect 14181 26754 14228 26756
rect 14136 26752 14228 26754
rect 14136 26696 14186 26752
rect 14136 26694 14228 26696
rect 14181 26692 14228 26694
rect 14292 26692 14298 26756
rect 15142 26692 15148 26756
rect 15212 26754 15218 26756
rect 17902 26754 17908 26756
rect 15212 26694 17908 26754
rect 15212 26692 15218 26694
rect 17902 26692 17908 26694
rect 17972 26754 17978 26756
rect 18321 26754 18387 26757
rect 19934 26754 19994 26830
rect 17972 26752 18387 26754
rect 17972 26696 18326 26752
rect 18382 26696 18387 26752
rect 17972 26694 18387 26696
rect 17972 26692 17978 26694
rect 14181 26691 14247 26692
rect 18321 26691 18387 26694
rect 19244 26694 19994 26754
rect 20529 26754 20595 26757
rect 20662 26754 20668 26756
rect 20529 26752 20668 26754
rect 20529 26696 20534 26752
rect 20590 26696 20668 26752
rect 20529 26694 20668 26696
rect 4787 26688 5103 26689
rect 4787 26624 4793 26688
rect 4857 26624 4873 26688
rect 4937 26624 4953 26688
rect 5017 26624 5033 26688
rect 5097 26624 5103 26688
rect 4787 26623 5103 26624
rect 12469 26688 12785 26689
rect 12469 26624 12475 26688
rect 12539 26624 12555 26688
rect 12619 26624 12635 26688
rect 12699 26624 12715 26688
rect 12779 26624 12785 26688
rect 12469 26623 12785 26624
rect 16021 26618 16087 26621
rect 17861 26618 17927 26621
rect 19244 26618 19304 26694
rect 20529 26691 20595 26694
rect 20662 26692 20668 26694
rect 20732 26754 20738 26756
rect 21544 26754 21604 26830
rect 24301 26827 24367 26830
rect 24894 26828 24900 26892
rect 24964 26890 24970 26892
rect 25129 26890 25195 26893
rect 24964 26888 25195 26890
rect 24964 26832 25134 26888
rect 25190 26832 25195 26888
rect 24964 26830 25195 26832
rect 24964 26828 24970 26830
rect 25129 26827 25195 26830
rect 25865 26890 25931 26893
rect 26233 26890 26299 26893
rect 26693 26892 26759 26893
rect 26693 26890 26740 26892
rect 25865 26888 26299 26890
rect 25865 26832 25870 26888
rect 25926 26832 26238 26888
rect 26294 26832 26299 26888
rect 25865 26830 26299 26832
rect 26648 26888 26740 26890
rect 26648 26832 26698 26888
rect 26648 26830 26740 26832
rect 25865 26827 25931 26830
rect 26233 26827 26299 26830
rect 26693 26828 26740 26830
rect 26804 26828 26810 26892
rect 29678 26890 29684 26892
rect 26926 26830 29684 26890
rect 26693 26827 26759 26828
rect 26926 26754 26986 26830
rect 29678 26828 29684 26830
rect 29748 26828 29754 26892
rect 29824 26890 29884 26966
rect 30414 26964 30420 27028
rect 30484 27026 30490 27028
rect 31845 27026 31911 27029
rect 30484 27024 31911 27026
rect 30484 26968 31850 27024
rect 31906 26968 31911 27024
rect 30484 26966 31911 26968
rect 30484 26964 30490 26966
rect 31845 26963 31911 26966
rect 32206 26936 33006 27056
rect 29824 26830 30390 26890
rect 28809 26754 28875 26757
rect 20732 26694 21604 26754
rect 21912 26694 26986 26754
rect 28214 26752 28875 26754
rect 28214 26696 28814 26752
rect 28870 26696 28875 26752
rect 28214 26694 28875 26696
rect 20732 26692 20738 26694
rect 20151 26688 20467 26689
rect 20151 26624 20157 26688
rect 20221 26624 20237 26688
rect 20301 26624 20317 26688
rect 20381 26624 20397 26688
rect 20461 26624 20467 26688
rect 20151 26623 20467 26624
rect 19425 26620 19491 26621
rect 16021 26616 17927 26618
rect 16021 26560 16026 26616
rect 16082 26560 17866 26616
rect 17922 26560 17927 26616
rect 16021 26558 17927 26560
rect 16021 26555 16087 26558
rect 17861 26555 17927 26558
rect 18324 26558 19304 26618
rect 12801 26482 12867 26485
rect 14774 26482 14780 26484
rect 12801 26480 14780 26482
rect 12801 26424 12806 26480
rect 12862 26424 14780 26480
rect 12801 26422 14780 26424
rect 12801 26419 12867 26422
rect 14774 26420 14780 26422
rect 14844 26420 14850 26484
rect 15326 26420 15332 26484
rect 15396 26482 15402 26484
rect 16798 26482 16804 26484
rect 15396 26422 16804 26482
rect 15396 26420 15402 26422
rect 16798 26420 16804 26422
rect 16868 26420 16874 26484
rect 17493 26482 17559 26485
rect 17953 26484 18019 26485
rect 18137 26484 18203 26485
rect 17902 26482 17908 26484
rect 17493 26480 17786 26482
rect 17493 26424 17498 26480
rect 17554 26424 17786 26480
rect 17493 26422 17786 26424
rect 17862 26422 17908 26482
rect 17972 26480 18019 26484
rect 18014 26424 18019 26480
rect 17493 26419 17559 26422
rect 9305 26346 9371 26349
rect 14958 26346 14964 26348
rect 9305 26344 14964 26346
rect 9305 26288 9310 26344
rect 9366 26288 14964 26344
rect 9305 26286 14964 26288
rect 9305 26283 9371 26286
rect 14958 26284 14964 26286
rect 15028 26346 15034 26348
rect 15101 26346 15167 26349
rect 15028 26344 15167 26346
rect 15028 26288 15106 26344
rect 15162 26288 15167 26344
rect 15028 26286 15167 26288
rect 15028 26284 15034 26286
rect 15101 26283 15167 26286
rect 15694 26284 15700 26348
rect 15764 26346 15770 26348
rect 16389 26346 16455 26349
rect 15764 26344 16455 26346
rect 15764 26288 16394 26344
rect 16450 26288 16455 26344
rect 15764 26286 16455 26288
rect 15764 26284 15770 26286
rect 16389 26283 16455 26286
rect 16798 26284 16804 26348
rect 16868 26346 16874 26348
rect 17585 26346 17651 26349
rect 16868 26344 17651 26346
rect 16868 26288 17590 26344
rect 17646 26288 17651 26344
rect 16868 26286 17651 26288
rect 17726 26346 17786 26422
rect 17902 26420 17908 26422
rect 17972 26420 18019 26424
rect 18086 26420 18092 26484
rect 18156 26482 18203 26484
rect 18156 26480 18248 26482
rect 18198 26424 18248 26480
rect 18156 26422 18248 26424
rect 18156 26420 18203 26422
rect 17953 26419 18019 26420
rect 18137 26419 18203 26420
rect 18324 26349 18384 26558
rect 19374 26556 19380 26620
rect 19444 26618 19491 26620
rect 19609 26618 19675 26621
rect 19926 26618 19932 26620
rect 19444 26616 19536 26618
rect 19486 26560 19536 26616
rect 19444 26558 19536 26560
rect 19609 26616 19932 26618
rect 19609 26560 19614 26616
rect 19670 26560 19932 26616
rect 19609 26558 19932 26560
rect 19444 26556 19491 26558
rect 19425 26555 19491 26556
rect 19609 26555 19675 26558
rect 19926 26556 19932 26558
rect 19996 26556 20002 26620
rect 20713 26618 20779 26621
rect 21766 26618 21772 26620
rect 20713 26616 21772 26618
rect 20713 26560 20718 26616
rect 20774 26560 21772 26616
rect 20713 26558 21772 26560
rect 20713 26555 20779 26558
rect 21766 26556 21772 26558
rect 21836 26556 21842 26620
rect 18638 26420 18644 26484
rect 18708 26482 18714 26484
rect 18708 26422 20592 26482
rect 18708 26420 18714 26422
rect 18086 26346 18092 26348
rect 17726 26286 18092 26346
rect 16868 26284 16874 26286
rect 17585 26283 17651 26286
rect 18086 26284 18092 26286
rect 18156 26284 18162 26348
rect 18321 26344 18387 26349
rect 18321 26288 18326 26344
rect 18382 26288 18387 26344
rect 18321 26283 18387 26288
rect 18597 26346 18663 26349
rect 20253 26346 20319 26349
rect 18597 26344 20319 26346
rect 18597 26288 18602 26344
rect 18658 26288 20258 26344
rect 20314 26288 20319 26344
rect 18597 26286 20319 26288
rect 20532 26346 20592 26422
rect 20662 26420 20668 26484
rect 20732 26482 20738 26484
rect 21265 26482 21331 26485
rect 20732 26480 21331 26482
rect 20732 26424 21270 26480
rect 21326 26424 21331 26480
rect 20732 26422 21331 26424
rect 20732 26420 20738 26422
rect 21265 26419 21331 26422
rect 20532 26286 20730 26346
rect 18597 26283 18663 26286
rect 20253 26283 20319 26286
rect 9673 26210 9739 26213
rect 13670 26210 13676 26212
rect 9673 26208 13676 26210
rect 9673 26152 9678 26208
rect 9734 26152 13676 26208
rect 9673 26150 13676 26152
rect 9673 26147 9739 26150
rect 13670 26148 13676 26150
rect 13740 26148 13746 26212
rect 13905 26210 13971 26213
rect 15929 26210 15995 26213
rect 13905 26208 15995 26210
rect 13905 26152 13910 26208
rect 13966 26152 15934 26208
rect 15990 26152 15995 26208
rect 13905 26150 15995 26152
rect 13905 26147 13971 26150
rect 15929 26147 15995 26150
rect 17217 26210 17283 26213
rect 18321 26210 18387 26213
rect 20670 26210 20730 26286
rect 20846 26284 20852 26348
rect 20916 26346 20922 26348
rect 21173 26346 21239 26349
rect 21912 26346 21972 26694
rect 27833 26688 28149 26689
rect 27833 26624 27839 26688
rect 27903 26624 27919 26688
rect 27983 26624 27999 26688
rect 28063 26624 28079 26688
rect 28143 26624 28149 26688
rect 27833 26623 28149 26624
rect 22093 26616 22159 26621
rect 22093 26560 22098 26616
rect 22154 26560 22159 26616
rect 22093 26555 22159 26560
rect 22277 26618 22343 26621
rect 23657 26618 23723 26621
rect 23841 26620 23907 26621
rect 22277 26616 23723 26618
rect 22277 26560 22282 26616
rect 22338 26560 23662 26616
rect 23718 26560 23723 26616
rect 22277 26558 23723 26560
rect 22277 26555 22343 26558
rect 23657 26555 23723 26558
rect 23790 26556 23796 26620
rect 23860 26618 23907 26620
rect 24117 26618 24183 26621
rect 24710 26618 24716 26620
rect 23860 26616 23952 26618
rect 23902 26560 23952 26616
rect 23860 26558 23952 26560
rect 24117 26616 24716 26618
rect 24117 26560 24122 26616
rect 24178 26560 24716 26616
rect 24117 26558 24716 26560
rect 23860 26556 23907 26558
rect 23841 26555 23907 26556
rect 24117 26555 24183 26558
rect 24710 26556 24716 26558
rect 24780 26556 24786 26620
rect 24945 26618 25011 26621
rect 26734 26618 26740 26620
rect 24945 26616 26740 26618
rect 24945 26560 24950 26616
rect 25006 26560 26740 26616
rect 24945 26558 26740 26560
rect 24945 26555 25011 26558
rect 26734 26556 26740 26558
rect 26804 26556 26810 26620
rect 27061 26618 27127 26621
rect 27654 26618 27660 26620
rect 27061 26616 27660 26618
rect 27061 26560 27066 26616
rect 27122 26560 27660 26616
rect 27061 26558 27660 26560
rect 27061 26555 27127 26558
rect 27654 26556 27660 26558
rect 27724 26556 27730 26620
rect 20916 26286 21052 26346
rect 20916 26284 20922 26286
rect 20846 26210 20852 26212
rect 17217 26208 18387 26210
rect 17217 26152 17222 26208
rect 17278 26152 18326 26208
rect 18382 26152 18387 26208
rect 17217 26150 18387 26152
rect 17217 26147 17283 26150
rect 18321 26147 18387 26150
rect 18600 26150 20592 26210
rect 20670 26150 20852 26210
rect 8628 26144 8944 26145
rect 0 26074 800 26104
rect 8628 26080 8634 26144
rect 8698 26080 8714 26144
rect 8778 26080 8794 26144
rect 8858 26080 8874 26144
rect 8938 26080 8944 26144
rect 8628 26079 8944 26080
rect 16310 26144 16626 26145
rect 16310 26080 16316 26144
rect 16380 26080 16396 26144
rect 16460 26080 16476 26144
rect 16540 26080 16556 26144
rect 16620 26080 16626 26144
rect 16310 26079 16626 26080
rect 18600 26077 18660 26150
rect 1577 26074 1643 26077
rect 0 26072 1643 26074
rect 0 26016 1582 26072
rect 1638 26016 1643 26072
rect 0 26014 1643 26016
rect 0 25984 800 26014
rect 1577 26011 1643 26014
rect 12341 26074 12407 26077
rect 13486 26074 13492 26076
rect 12341 26072 13492 26074
rect 12341 26016 12346 26072
rect 12402 26016 13492 26072
rect 12341 26014 13492 26016
rect 12341 26011 12407 26014
rect 13486 26012 13492 26014
rect 13556 26012 13562 26076
rect 13629 26074 13695 26077
rect 14038 26074 14044 26076
rect 13629 26072 14044 26074
rect 13629 26016 13634 26072
rect 13690 26016 14044 26072
rect 13629 26014 14044 26016
rect 13629 26011 13695 26014
rect 14038 26012 14044 26014
rect 14108 26012 14114 26076
rect 15285 26074 15351 26077
rect 15745 26074 15811 26077
rect 15285 26072 15811 26074
rect 15285 26016 15290 26072
rect 15346 26016 15750 26072
rect 15806 26016 15811 26072
rect 15285 26014 15811 26016
rect 15285 26011 15351 26014
rect 15745 26011 15811 26014
rect 17166 26012 17172 26076
rect 17236 26074 17242 26076
rect 17309 26074 17375 26077
rect 18086 26074 18092 26076
rect 17236 26072 17375 26074
rect 17236 26016 17314 26072
rect 17370 26016 17375 26072
rect 17236 26014 17375 26016
rect 17236 26012 17242 26014
rect 17309 26011 17375 26014
rect 17910 26014 18092 26074
rect 14457 25938 14523 25941
rect 14590 25938 14596 25940
rect 14457 25936 14596 25938
rect 14457 25880 14462 25936
rect 14518 25880 14596 25936
rect 14457 25878 14596 25880
rect 14457 25875 14523 25878
rect 14590 25876 14596 25878
rect 14660 25938 14666 25940
rect 15285 25938 15351 25941
rect 14660 25936 15351 25938
rect 14660 25880 15290 25936
rect 15346 25880 15351 25936
rect 14660 25878 15351 25880
rect 14660 25876 14666 25878
rect 15285 25875 15351 25878
rect 15561 25938 15627 25941
rect 17910 25938 17970 26014
rect 18086 26012 18092 26014
rect 18156 26012 18162 26076
rect 18229 26074 18295 26077
rect 18413 26074 18479 26077
rect 18229 26072 18479 26074
rect 18229 26016 18234 26072
rect 18290 26016 18418 26072
rect 18474 26016 18479 26072
rect 18229 26014 18479 26016
rect 18229 26011 18295 26014
rect 18413 26011 18479 26014
rect 18597 26072 18663 26077
rect 18597 26016 18602 26072
rect 18658 26016 18663 26072
rect 18597 26011 18663 26016
rect 19057 26074 19123 26077
rect 20532 26074 20592 26150
rect 20846 26148 20852 26150
rect 20916 26148 20922 26212
rect 20662 26074 20668 26076
rect 19057 26072 20132 26074
rect 19057 26016 19062 26072
rect 19118 26016 20132 26072
rect 19057 26014 20132 26016
rect 20532 26014 20668 26074
rect 19057 26011 19123 26014
rect 15561 25936 17970 25938
rect 15561 25880 15566 25936
rect 15622 25880 17970 25936
rect 15561 25878 17970 25880
rect 18413 25938 18479 25941
rect 19926 25938 19932 25940
rect 18413 25936 19932 25938
rect 18413 25880 18418 25936
rect 18474 25880 19932 25936
rect 18413 25878 19932 25880
rect 15561 25875 15627 25878
rect 18413 25875 18479 25878
rect 19926 25876 19932 25878
rect 19996 25876 20002 25940
rect 20072 25938 20132 26014
rect 20662 26012 20668 26014
rect 20732 26012 20738 26076
rect 20992 26074 21052 26286
rect 21173 26344 21972 26346
rect 21173 26288 21178 26344
rect 21234 26288 21972 26344
rect 21173 26286 21972 26288
rect 22096 26346 22156 26555
rect 22369 26482 22435 26485
rect 28214 26482 28274 26694
rect 28809 26691 28875 26694
rect 28349 26618 28415 26621
rect 28758 26618 28764 26620
rect 28349 26616 28764 26618
rect 28349 26560 28354 26616
rect 28410 26560 28764 26616
rect 28349 26558 28764 26560
rect 28349 26555 28415 26558
rect 28758 26556 28764 26558
rect 28828 26556 28834 26620
rect 29494 26618 29500 26620
rect 28904 26558 29500 26618
rect 28904 26485 28964 26558
rect 29494 26556 29500 26558
rect 29564 26556 29570 26620
rect 29686 26618 29746 26828
rect 30330 26754 30390 26830
rect 32765 26754 32831 26757
rect 30330 26752 32831 26754
rect 30330 26696 32770 26752
rect 32826 26696 32831 26752
rect 30330 26694 32831 26696
rect 32765 26691 32831 26694
rect 30046 26618 30052 26620
rect 29686 26558 30052 26618
rect 30046 26556 30052 26558
rect 30116 26556 30122 26620
rect 30598 26618 30604 26620
rect 30284 26558 30604 26618
rect 22369 26480 28274 26482
rect 22369 26424 22374 26480
rect 22430 26424 28274 26480
rect 22369 26422 28274 26424
rect 22369 26419 22435 26422
rect 28390 26420 28396 26484
rect 28460 26482 28466 26484
rect 28533 26482 28599 26485
rect 28460 26480 28599 26482
rect 28460 26424 28538 26480
rect 28594 26424 28599 26480
rect 28460 26422 28599 26424
rect 28460 26420 28466 26422
rect 28533 26419 28599 26422
rect 28901 26480 28967 26485
rect 28901 26424 28906 26480
rect 28962 26424 28967 26480
rect 28901 26419 28967 26424
rect 29085 26482 29151 26485
rect 29494 26482 29500 26484
rect 29085 26480 29500 26482
rect 29085 26424 29090 26480
rect 29146 26424 29500 26480
rect 29085 26422 29500 26424
rect 29085 26419 29151 26422
rect 29494 26420 29500 26422
rect 29564 26420 29570 26484
rect 30097 26482 30163 26485
rect 30284 26482 30344 26558
rect 30598 26556 30604 26558
rect 30668 26556 30674 26620
rect 32121 26618 32187 26621
rect 30974 26616 32187 26618
rect 30974 26560 32126 26616
rect 32182 26560 32187 26616
rect 30974 26558 32187 26560
rect 30097 26480 30344 26482
rect 30097 26424 30102 26480
rect 30158 26424 30344 26480
rect 30097 26422 30344 26424
rect 30097 26419 30163 26422
rect 30414 26420 30420 26484
rect 30484 26482 30490 26484
rect 30833 26482 30899 26485
rect 30484 26480 30899 26482
rect 30484 26424 30838 26480
rect 30894 26424 30899 26480
rect 30484 26422 30899 26424
rect 30484 26420 30490 26422
rect 30833 26419 30899 26422
rect 24209 26346 24275 26349
rect 24710 26346 24716 26348
rect 22096 26286 22938 26346
rect 21173 26283 21239 26286
rect 21173 26212 21239 26213
rect 21173 26210 21220 26212
rect 21128 26208 21220 26210
rect 21128 26152 21178 26208
rect 21128 26150 21220 26152
rect 21173 26148 21220 26150
rect 21284 26148 21290 26212
rect 21357 26210 21423 26213
rect 22185 26210 22251 26213
rect 21357 26208 22251 26210
rect 21357 26152 21362 26208
rect 21418 26152 22190 26208
rect 22246 26152 22251 26208
rect 21357 26150 22251 26152
rect 21173 26147 21239 26148
rect 21357 26147 21423 26150
rect 22185 26147 22251 26150
rect 22369 26074 22435 26077
rect 20808 26072 22435 26074
rect 20808 26016 22374 26072
rect 22430 26016 22435 26072
rect 20808 26014 22435 26016
rect 20808 25938 20868 26014
rect 22369 26011 22435 26014
rect 22553 26074 22619 26077
rect 22878 26074 22938 26286
rect 24209 26344 24716 26346
rect 24209 26288 24214 26344
rect 24270 26288 24716 26344
rect 24209 26286 24716 26288
rect 24209 26283 24275 26286
rect 24710 26284 24716 26286
rect 24780 26284 24786 26348
rect 24894 26284 24900 26348
rect 24964 26346 24970 26348
rect 25037 26346 25103 26349
rect 24964 26344 25103 26346
rect 24964 26288 25042 26344
rect 25098 26288 25103 26344
rect 24964 26286 25103 26288
rect 24964 26284 24970 26286
rect 25037 26283 25103 26286
rect 25446 26284 25452 26348
rect 25516 26346 25522 26348
rect 27286 26346 27292 26348
rect 25516 26286 27292 26346
rect 25516 26284 25522 26286
rect 27286 26284 27292 26286
rect 27356 26346 27362 26348
rect 27521 26346 27587 26349
rect 27356 26344 27587 26346
rect 27356 26288 27526 26344
rect 27582 26288 27587 26344
rect 27356 26286 27587 26288
rect 27356 26284 27362 26286
rect 27521 26283 27587 26286
rect 27889 26346 27955 26349
rect 28717 26348 28783 26349
rect 28206 26346 28212 26348
rect 27889 26344 28212 26346
rect 27889 26288 27894 26344
rect 27950 26288 28212 26344
rect 27889 26286 28212 26288
rect 27889 26283 27955 26286
rect 28206 26284 28212 26286
rect 28276 26284 28282 26348
rect 28717 26346 28764 26348
rect 28672 26344 28764 26346
rect 28672 26288 28722 26344
rect 28672 26286 28764 26288
rect 28717 26284 28764 26286
rect 28828 26284 28834 26348
rect 29085 26346 29151 26349
rect 29678 26346 29684 26348
rect 29085 26344 29684 26346
rect 29085 26288 29090 26344
rect 29146 26288 29684 26344
rect 29085 26286 29684 26288
rect 28717 26283 28783 26284
rect 29085 26283 29151 26286
rect 29678 26284 29684 26286
rect 29748 26284 29754 26348
rect 30833 26346 30899 26349
rect 30974 26346 31034 26558
rect 32121 26555 32187 26558
rect 30833 26344 31034 26346
rect 30833 26288 30838 26344
rect 30894 26288 31034 26344
rect 30833 26286 31034 26288
rect 32029 26346 32095 26349
rect 32206 26346 33006 26376
rect 32029 26344 33006 26346
rect 32029 26288 32034 26344
rect 32090 26288 33006 26344
rect 32029 26286 33006 26288
rect 30833 26283 30899 26286
rect 32029 26283 32095 26286
rect 32206 26256 33006 26286
rect 23054 26148 23060 26212
rect 23124 26210 23130 26212
rect 23790 26210 23796 26212
rect 23124 26150 23796 26210
rect 23124 26148 23130 26150
rect 23790 26148 23796 26150
rect 23860 26148 23866 26212
rect 25497 26210 25563 26213
rect 25681 26210 25747 26213
rect 25497 26208 25747 26210
rect 25497 26152 25502 26208
rect 25558 26152 25686 26208
rect 25742 26152 25747 26208
rect 25497 26150 25747 26152
rect 25497 26147 25563 26150
rect 25681 26147 25747 26150
rect 26785 26210 26851 26213
rect 31017 26210 31083 26213
rect 26785 26208 31083 26210
rect 26785 26152 26790 26208
rect 26846 26152 31022 26208
rect 31078 26152 31083 26208
rect 26785 26150 31083 26152
rect 26785 26147 26851 26150
rect 31017 26147 31083 26150
rect 23992 26144 24308 26145
rect 23992 26080 23998 26144
rect 24062 26080 24078 26144
rect 24142 26080 24158 26144
rect 24222 26080 24238 26144
rect 24302 26080 24308 26144
rect 23992 26079 24308 26080
rect 31674 26144 31990 26145
rect 31674 26080 31680 26144
rect 31744 26080 31760 26144
rect 31824 26080 31840 26144
rect 31904 26080 31920 26144
rect 31984 26080 31990 26144
rect 31674 26079 31990 26080
rect 23054 26074 23060 26076
rect 22553 26072 22754 26074
rect 22553 26016 22558 26072
rect 22614 26016 22754 26072
rect 22553 26014 22754 26016
rect 22878 26014 23060 26074
rect 22553 26011 22619 26014
rect 21265 25940 21331 25941
rect 20072 25878 20868 25938
rect 21214 25876 21220 25940
rect 21284 25938 21331 25940
rect 21817 25938 21883 25941
rect 22461 25938 22527 25941
rect 21284 25936 21376 25938
rect 21326 25880 21376 25936
rect 21284 25878 21376 25880
rect 21817 25936 22527 25938
rect 21817 25880 21822 25936
rect 21878 25880 22466 25936
rect 22522 25880 22527 25936
rect 21817 25878 22527 25880
rect 22694 25938 22754 26014
rect 23054 26012 23060 26014
rect 23124 26012 23130 26076
rect 24761 26074 24827 26077
rect 24894 26074 24900 26076
rect 24761 26072 24900 26074
rect 24761 26016 24766 26072
rect 24822 26016 24900 26072
rect 24761 26014 24900 26016
rect 24761 26011 24827 26014
rect 24894 26012 24900 26014
rect 24964 26012 24970 26076
rect 25865 26074 25931 26077
rect 28390 26074 28396 26076
rect 25865 26072 28396 26074
rect 25865 26016 25870 26072
rect 25926 26016 28396 26072
rect 25865 26014 28396 26016
rect 25865 26011 25931 26014
rect 28390 26012 28396 26014
rect 28460 26012 28466 26076
rect 29269 26074 29335 26077
rect 28996 26072 29335 26074
rect 28996 26016 29274 26072
rect 29330 26016 29335 26072
rect 28996 26014 29335 26016
rect 24388 25938 24394 25940
rect 22694 25878 24394 25938
rect 21284 25876 21331 25878
rect 21265 25875 21331 25876
rect 21817 25875 21883 25878
rect 22461 25875 22527 25878
rect 24388 25876 24394 25878
rect 24458 25938 24464 25940
rect 25589 25938 25655 25941
rect 24458 25936 25655 25938
rect 24458 25880 25594 25936
rect 25650 25880 25655 25936
rect 24458 25878 25655 25880
rect 24458 25876 24464 25878
rect 25589 25875 25655 25878
rect 25865 25938 25931 25941
rect 25998 25938 26004 25940
rect 25865 25936 26004 25938
rect 25865 25880 25870 25936
rect 25926 25880 26004 25936
rect 25865 25878 26004 25880
rect 25865 25875 25931 25878
rect 25998 25876 26004 25878
rect 26068 25876 26074 25940
rect 28165 25938 28231 25941
rect 28996 25938 29056 26014
rect 29269 26011 29335 26014
rect 29821 26074 29887 26077
rect 30782 26074 30788 26076
rect 29821 26072 30788 26074
rect 29821 26016 29826 26072
rect 29882 26016 30788 26072
rect 29821 26014 30788 26016
rect 29821 26011 29887 26014
rect 30782 26012 30788 26014
rect 30852 26012 30858 26076
rect 26374 25936 29056 25938
rect 26374 25880 28170 25936
rect 28226 25880 29056 25936
rect 26374 25878 29056 25880
rect 29177 25938 29243 25941
rect 29177 25936 29562 25938
rect 29177 25880 29182 25936
rect 29238 25880 29562 25936
rect 29177 25878 29562 25880
rect 8385 25802 8451 25805
rect 13629 25802 13695 25805
rect 19793 25802 19859 25805
rect 8385 25800 13554 25802
rect 8385 25744 8390 25800
rect 8446 25744 13554 25800
rect 8385 25742 13554 25744
rect 8385 25739 8451 25742
rect 13494 25666 13554 25742
rect 13629 25800 19859 25802
rect 13629 25744 13634 25800
rect 13690 25744 19798 25800
rect 19854 25744 19859 25800
rect 13629 25742 19859 25744
rect 13629 25739 13695 25742
rect 19793 25739 19859 25742
rect 20069 25802 20135 25805
rect 21357 25802 21423 25805
rect 24209 25802 24275 25805
rect 20069 25800 20730 25802
rect 20069 25744 20074 25800
rect 20130 25744 20730 25800
rect 20069 25742 20730 25744
rect 20069 25739 20135 25742
rect 17534 25666 17540 25668
rect 13494 25606 17540 25666
rect 17534 25604 17540 25606
rect 17604 25666 17610 25668
rect 17677 25666 17743 25669
rect 17604 25664 17743 25666
rect 17604 25608 17682 25664
rect 17738 25608 17743 25664
rect 17604 25606 17743 25608
rect 17604 25604 17610 25606
rect 17677 25603 17743 25606
rect 18873 25666 18939 25669
rect 19190 25666 19196 25668
rect 18873 25664 19196 25666
rect 18873 25608 18878 25664
rect 18934 25608 19196 25664
rect 18873 25606 19196 25608
rect 18873 25603 18939 25606
rect 19190 25604 19196 25606
rect 19260 25604 19266 25668
rect 20670 25666 20730 25742
rect 21357 25800 24275 25802
rect 21357 25744 21362 25800
rect 21418 25744 24214 25800
rect 24270 25744 24275 25800
rect 21357 25742 24275 25744
rect 21357 25739 21423 25742
rect 24209 25739 24275 25742
rect 25078 25740 25084 25804
rect 25148 25802 25154 25804
rect 26374 25802 26434 25878
rect 28165 25875 28231 25878
rect 29177 25875 29243 25878
rect 25148 25742 26434 25802
rect 26509 25802 26575 25805
rect 27521 25802 27587 25805
rect 26509 25800 27587 25802
rect 26509 25744 26514 25800
rect 26570 25744 27526 25800
rect 27582 25744 27587 25800
rect 26509 25742 27587 25744
rect 25148 25740 25154 25742
rect 26509 25739 26575 25742
rect 27521 25739 27587 25742
rect 27654 25740 27660 25804
rect 27724 25802 27730 25804
rect 29361 25802 29427 25805
rect 27724 25800 29427 25802
rect 27724 25744 29366 25800
rect 29422 25744 29427 25800
rect 27724 25742 29427 25744
rect 29502 25802 29562 25878
rect 29862 25876 29868 25940
rect 29932 25938 29938 25940
rect 30373 25938 30439 25941
rect 32489 25938 32555 25941
rect 29932 25936 30439 25938
rect 29932 25880 30378 25936
rect 30434 25880 30439 25936
rect 29932 25878 30439 25880
rect 29932 25876 29938 25878
rect 30373 25875 30439 25878
rect 30560 25936 32555 25938
rect 30560 25880 32494 25936
rect 32550 25880 32555 25936
rect 30560 25878 32555 25880
rect 30560 25802 30620 25878
rect 32489 25875 32555 25878
rect 29502 25742 30620 25802
rect 27724 25740 27730 25742
rect 29361 25739 29427 25742
rect 24945 25666 25011 25669
rect 20670 25664 25011 25666
rect 20670 25608 24950 25664
rect 25006 25608 25011 25664
rect 20670 25606 25011 25608
rect 24945 25603 25011 25606
rect 26509 25666 26575 25669
rect 27429 25666 27495 25669
rect 27654 25666 27660 25668
rect 26509 25664 27495 25666
rect 26509 25608 26514 25664
rect 26570 25608 27434 25664
rect 27490 25608 27495 25664
rect 26509 25606 27495 25608
rect 26509 25603 26575 25606
rect 27429 25603 27495 25606
rect 27616 25604 27660 25666
rect 27724 25604 27730 25668
rect 29126 25604 29132 25668
rect 29196 25666 29202 25668
rect 29637 25666 29703 25669
rect 29196 25664 29703 25666
rect 29196 25608 29642 25664
rect 29698 25608 29703 25664
rect 29196 25606 29703 25608
rect 29196 25604 29202 25606
rect 4787 25600 5103 25601
rect 4787 25536 4793 25600
rect 4857 25536 4873 25600
rect 4937 25536 4953 25600
rect 5017 25536 5033 25600
rect 5097 25536 5103 25600
rect 4787 25535 5103 25536
rect 12469 25600 12785 25601
rect 12469 25536 12475 25600
rect 12539 25536 12555 25600
rect 12619 25536 12635 25600
rect 12699 25536 12715 25600
rect 12779 25536 12785 25600
rect 12469 25535 12785 25536
rect 20151 25600 20467 25601
rect 20151 25536 20157 25600
rect 20221 25536 20237 25600
rect 20301 25536 20317 25600
rect 20381 25536 20397 25600
rect 20461 25536 20467 25600
rect 20151 25535 20467 25536
rect 27616 25533 27676 25604
rect 29637 25603 29703 25606
rect 29821 25666 29887 25669
rect 30598 25666 30604 25668
rect 29821 25664 30604 25666
rect 29821 25608 29826 25664
rect 29882 25608 30604 25664
rect 29821 25606 30604 25608
rect 29821 25603 29887 25606
rect 30598 25604 30604 25606
rect 30668 25604 30674 25668
rect 31293 25666 31359 25669
rect 32206 25666 33006 25696
rect 31293 25664 33006 25666
rect 31293 25608 31298 25664
rect 31354 25608 33006 25664
rect 31293 25606 33006 25608
rect 31293 25603 31359 25606
rect 27833 25600 28149 25601
rect 27833 25536 27839 25600
rect 27903 25536 27919 25600
rect 27983 25536 27999 25600
rect 28063 25536 28079 25600
rect 28143 25536 28149 25600
rect 32206 25576 33006 25606
rect 27833 25535 28149 25536
rect 5390 25468 5396 25532
rect 5460 25530 5466 25532
rect 12014 25530 12020 25532
rect 5460 25470 12020 25530
rect 5460 25468 5466 25470
rect 12014 25468 12020 25470
rect 12084 25468 12090 25532
rect 12893 25530 12959 25533
rect 13721 25530 13787 25533
rect 14273 25532 14339 25533
rect 12893 25528 13787 25530
rect 12893 25472 12898 25528
rect 12954 25472 13726 25528
rect 13782 25472 13787 25528
rect 12893 25470 13787 25472
rect 12893 25467 12959 25470
rect 13721 25467 13787 25470
rect 14222 25468 14228 25532
rect 14292 25530 14339 25532
rect 14292 25528 14384 25530
rect 14334 25472 14384 25528
rect 14292 25470 14384 25472
rect 14292 25468 14339 25470
rect 14590 25468 14596 25532
rect 14660 25530 14666 25532
rect 14733 25530 14799 25533
rect 14660 25528 14799 25530
rect 14660 25472 14738 25528
rect 14794 25472 14799 25528
rect 14660 25470 14799 25472
rect 14660 25468 14666 25470
rect 14273 25467 14339 25468
rect 14733 25467 14799 25470
rect 15929 25530 15995 25533
rect 16757 25530 16823 25533
rect 15929 25528 16823 25530
rect 15929 25472 15934 25528
rect 15990 25472 16762 25528
rect 16818 25472 16823 25528
rect 15929 25470 16823 25472
rect 15929 25467 15995 25470
rect 16757 25467 16823 25470
rect 17125 25530 17191 25533
rect 17350 25530 17356 25532
rect 17125 25528 17356 25530
rect 17125 25472 17130 25528
rect 17186 25472 17356 25528
rect 17125 25470 17356 25472
rect 17125 25467 17191 25470
rect 17350 25468 17356 25470
rect 17420 25468 17426 25532
rect 17493 25530 17559 25533
rect 17493 25528 19810 25530
rect 17493 25472 17498 25528
rect 17554 25472 19810 25528
rect 17493 25470 19810 25472
rect 17493 25467 17559 25470
rect 9489 25394 9555 25397
rect 19333 25394 19399 25397
rect 9489 25392 19399 25394
rect 9489 25336 9494 25392
rect 9550 25336 19338 25392
rect 19394 25336 19399 25392
rect 9489 25334 19399 25336
rect 9489 25331 9555 25334
rect 19333 25331 19399 25334
rect 19517 25396 19583 25397
rect 19517 25392 19564 25396
rect 19628 25394 19634 25396
rect 19750 25394 19810 25470
rect 20662 25468 20668 25532
rect 20732 25530 20738 25532
rect 24117 25530 24183 25533
rect 20732 25528 24183 25530
rect 20732 25472 24122 25528
rect 24178 25472 24183 25528
rect 20732 25470 24183 25472
rect 20732 25468 20738 25470
rect 24117 25467 24183 25470
rect 24485 25530 24551 25533
rect 25262 25530 25268 25532
rect 24485 25528 25268 25530
rect 24485 25472 24490 25528
rect 24546 25472 25268 25528
rect 24485 25470 25268 25472
rect 24485 25467 24551 25470
rect 25262 25468 25268 25470
rect 25332 25530 25338 25532
rect 27429 25530 27495 25533
rect 25332 25528 27495 25530
rect 25332 25472 27434 25528
rect 27490 25472 27495 25528
rect 25332 25470 27495 25472
rect 25332 25468 25338 25470
rect 27429 25467 27495 25470
rect 27613 25528 27679 25533
rect 27613 25472 27618 25528
rect 27674 25472 27679 25528
rect 27613 25467 27679 25472
rect 28257 25530 28323 25533
rect 29126 25530 29132 25532
rect 28257 25528 29132 25530
rect 28257 25472 28262 25528
rect 28318 25472 29132 25528
rect 28257 25470 29132 25472
rect 28257 25467 28323 25470
rect 29126 25468 29132 25470
rect 29196 25468 29202 25532
rect 29637 25530 29703 25533
rect 32070 25530 32076 25532
rect 29637 25528 32076 25530
rect 29637 25472 29642 25528
rect 29698 25472 32076 25528
rect 29637 25470 32076 25472
rect 29637 25467 29703 25470
rect 32070 25468 32076 25470
rect 32140 25468 32146 25532
rect 21909 25394 21975 25397
rect 19517 25336 19522 25392
rect 19517 25332 19564 25336
rect 19628 25334 19674 25394
rect 19750 25392 21975 25394
rect 19750 25336 21914 25392
rect 21970 25336 21975 25392
rect 19750 25334 21975 25336
rect 19628 25332 19634 25334
rect 19517 25331 19583 25332
rect 21909 25331 21975 25334
rect 22185 25394 22251 25397
rect 23381 25394 23447 25397
rect 23657 25396 23723 25397
rect 23606 25394 23612 25396
rect 22185 25392 23447 25394
rect 22185 25336 22190 25392
rect 22246 25336 23386 25392
rect 23442 25336 23447 25392
rect 22185 25334 23447 25336
rect 23566 25334 23612 25394
rect 23676 25392 23723 25396
rect 23718 25336 23723 25392
rect 22185 25331 22251 25334
rect 23381 25331 23447 25334
rect 23606 25332 23612 25334
rect 23676 25332 23723 25336
rect 23657 25331 23723 25332
rect 24301 25394 24367 25397
rect 24526 25394 24532 25396
rect 24301 25392 24532 25394
rect 24301 25336 24306 25392
rect 24362 25336 24532 25392
rect 24301 25334 24532 25336
rect 24301 25331 24367 25334
rect 24526 25332 24532 25334
rect 24596 25332 24602 25396
rect 24761 25394 24827 25397
rect 30925 25394 30991 25397
rect 24761 25392 30991 25394
rect 24761 25336 24766 25392
rect 24822 25336 30930 25392
rect 30986 25336 30991 25392
rect 24761 25334 30991 25336
rect 24761 25331 24827 25334
rect 30925 25331 30991 25334
rect 31150 25332 31156 25396
rect 31220 25394 31226 25396
rect 31293 25394 31359 25397
rect 32489 25396 32555 25397
rect 32438 25394 32444 25396
rect 31220 25392 31359 25394
rect 31220 25336 31298 25392
rect 31354 25336 31359 25392
rect 31220 25334 31359 25336
rect 32398 25334 32444 25394
rect 32508 25392 32555 25396
rect 32550 25336 32555 25392
rect 31220 25332 31226 25334
rect 31293 25331 31359 25334
rect 32438 25332 32444 25334
rect 32508 25332 32555 25336
rect 32489 25331 32555 25332
rect 0 25258 800 25288
rect 1577 25258 1643 25261
rect 0 25256 1643 25258
rect 0 25200 1582 25256
rect 1638 25200 1643 25256
rect 0 25198 1643 25200
rect 0 25168 800 25198
rect 1577 25195 1643 25198
rect 12157 25258 12223 25261
rect 14457 25258 14523 25261
rect 14590 25258 14596 25260
rect 12157 25256 14596 25258
rect 12157 25200 12162 25256
rect 12218 25200 14462 25256
rect 14518 25200 14596 25256
rect 12157 25198 14596 25200
rect 12157 25195 12223 25198
rect 14457 25195 14523 25198
rect 14590 25196 14596 25198
rect 14660 25196 14666 25260
rect 14774 25196 14780 25260
rect 14844 25258 14850 25260
rect 15929 25258 15995 25261
rect 14844 25256 15995 25258
rect 14844 25200 15934 25256
rect 15990 25200 15995 25256
rect 14844 25198 15995 25200
rect 14844 25196 14850 25198
rect 15929 25195 15995 25198
rect 17585 25258 17651 25261
rect 20069 25258 20135 25261
rect 21357 25258 21423 25261
rect 22553 25258 22619 25261
rect 23565 25258 23631 25261
rect 17585 25256 22432 25258
rect 17585 25200 17590 25256
rect 17646 25200 20074 25256
rect 20130 25200 21362 25256
rect 21418 25200 22432 25256
rect 17585 25198 22432 25200
rect 17585 25195 17651 25198
rect 20069 25195 20135 25198
rect 21357 25195 21423 25198
rect 10225 25122 10291 25125
rect 14089 25122 14155 25125
rect 15929 25122 15995 25125
rect 10225 25120 14155 25122
rect 10225 25064 10230 25120
rect 10286 25064 14094 25120
rect 14150 25064 14155 25120
rect 10225 25062 14155 25064
rect 10225 25059 10291 25062
rect 14089 25059 14155 25062
rect 14782 25120 15995 25122
rect 14782 25064 15934 25120
rect 15990 25064 15995 25120
rect 14782 25062 15995 25064
rect 8628 25056 8944 25057
rect 8628 24992 8634 25056
rect 8698 24992 8714 25056
rect 8778 24992 8794 25056
rect 8858 24992 8874 25056
rect 8938 24992 8944 25056
rect 8628 24991 8944 24992
rect 12801 24986 12867 24989
rect 13261 24986 13327 24989
rect 14782 24986 14842 25062
rect 15929 25059 15995 25062
rect 17534 25060 17540 25124
rect 17604 25122 17610 25124
rect 17769 25122 17835 25125
rect 17604 25120 17835 25122
rect 17604 25064 17774 25120
rect 17830 25064 17835 25120
rect 17604 25062 17835 25064
rect 17604 25060 17610 25062
rect 17769 25059 17835 25062
rect 17953 25122 18019 25125
rect 20662 25122 20668 25124
rect 17953 25120 20668 25122
rect 17953 25064 17958 25120
rect 18014 25064 20668 25120
rect 17953 25062 20668 25064
rect 17953 25059 18019 25062
rect 20662 25060 20668 25062
rect 20732 25060 20738 25124
rect 21725 25122 21791 25125
rect 21544 25120 21791 25122
rect 21544 25064 21730 25120
rect 21786 25064 21791 25120
rect 21544 25062 21791 25064
rect 16310 25056 16626 25057
rect 16310 24992 16316 25056
rect 16380 24992 16396 25056
rect 16460 24992 16476 25056
rect 16540 24992 16556 25056
rect 16620 24992 16626 25056
rect 16310 24991 16626 24992
rect 21544 24989 21604 25062
rect 21725 25059 21791 25062
rect 21909 25122 21975 25125
rect 22372 25122 22432 25198
rect 22553 25256 23631 25258
rect 22553 25200 22558 25256
rect 22614 25200 23570 25256
rect 23626 25200 23631 25256
rect 22553 25198 23631 25200
rect 22553 25195 22619 25198
rect 23565 25195 23631 25198
rect 24025 25258 24091 25261
rect 24485 25258 24551 25261
rect 24025 25256 24551 25258
rect 24025 25200 24030 25256
rect 24086 25200 24490 25256
rect 24546 25200 24551 25256
rect 24025 25198 24551 25200
rect 24025 25195 24091 25198
rect 24485 25195 24551 25198
rect 25262 25196 25268 25260
rect 25332 25258 25338 25260
rect 29729 25258 29795 25261
rect 25332 25256 29795 25258
rect 25332 25200 29734 25256
rect 29790 25200 29795 25256
rect 25332 25198 29795 25200
rect 25332 25196 25338 25198
rect 29729 25195 29795 25198
rect 30598 25196 30604 25260
rect 30668 25258 30674 25260
rect 32622 25258 32628 25260
rect 30668 25198 32628 25258
rect 30668 25196 30674 25198
rect 32622 25196 32628 25198
rect 32692 25196 32698 25260
rect 24393 25122 24459 25125
rect 25773 25122 25839 25125
rect 21909 25120 22202 25122
rect 21909 25064 21914 25120
rect 21970 25064 22202 25120
rect 21909 25062 22202 25064
rect 22372 25062 23490 25122
rect 21909 25059 21975 25062
rect 12801 24984 14842 24986
rect 12801 24928 12806 24984
rect 12862 24928 13266 24984
rect 13322 24928 14842 24984
rect 12801 24926 14842 24928
rect 14917 24986 14983 24989
rect 15878 24986 15884 24988
rect 14917 24984 15884 24986
rect 14917 24928 14922 24984
rect 14978 24928 15884 24984
rect 14917 24926 15884 24928
rect 12801 24923 12867 24926
rect 13261 24923 13327 24926
rect 14917 24923 14983 24926
rect 15878 24924 15884 24926
rect 15948 24924 15954 24988
rect 16757 24986 16823 24989
rect 18638 24986 18644 24988
rect 16757 24984 18644 24986
rect 16757 24928 16762 24984
rect 16818 24928 18644 24984
rect 16757 24926 18644 24928
rect 16757 24923 16823 24926
rect 18638 24924 18644 24926
rect 18708 24924 18714 24988
rect 18781 24986 18847 24989
rect 19057 24986 19123 24989
rect 18781 24984 19123 24986
rect 18781 24928 18786 24984
rect 18842 24928 19062 24984
rect 19118 24928 19123 24984
rect 18781 24926 19123 24928
rect 18781 24923 18847 24926
rect 19057 24923 19123 24926
rect 19425 24986 19491 24989
rect 20345 24986 20411 24989
rect 20524 24986 20530 24988
rect 19425 24984 20530 24986
rect 19425 24928 19430 24984
rect 19486 24928 20350 24984
rect 20406 24928 20530 24984
rect 19425 24926 20530 24928
rect 19425 24923 19491 24926
rect 20345 24923 20411 24926
rect 20524 24924 20530 24926
rect 20594 24924 20600 24988
rect 21081 24986 21147 24989
rect 21398 24986 21404 24988
rect 21081 24984 21404 24986
rect 21081 24928 21086 24984
rect 21142 24928 21404 24984
rect 21081 24926 21404 24928
rect 21081 24923 21147 24926
rect 21398 24924 21404 24926
rect 21468 24924 21474 24988
rect 21541 24984 21607 24989
rect 21541 24928 21546 24984
rect 21602 24928 21607 24984
rect 21541 24923 21607 24928
rect 21766 24924 21772 24988
rect 21836 24986 21842 24988
rect 22001 24986 22067 24989
rect 21836 24984 22067 24986
rect 21836 24928 22006 24984
rect 22062 24928 22067 24984
rect 21836 24926 22067 24928
rect 22142 24986 22202 25062
rect 22686 24986 22692 24988
rect 22142 24926 22692 24986
rect 21836 24924 21842 24926
rect 22001 24923 22067 24926
rect 22686 24924 22692 24926
rect 22756 24924 22762 24988
rect 9213 24850 9279 24853
rect 13905 24850 13971 24853
rect 9213 24848 13971 24850
rect 9213 24792 9218 24848
rect 9274 24792 13910 24848
rect 13966 24792 13971 24848
rect 9213 24790 13971 24792
rect 9213 24787 9279 24790
rect 13905 24787 13971 24790
rect 14733 24850 14799 24853
rect 15510 24850 15516 24852
rect 14733 24848 15516 24850
rect 14733 24792 14738 24848
rect 14794 24792 15516 24848
rect 14733 24790 15516 24792
rect 14733 24787 14799 24790
rect 15510 24788 15516 24790
rect 15580 24850 15586 24852
rect 17125 24850 17191 24853
rect 15580 24848 17191 24850
rect 15580 24792 17130 24848
rect 17186 24792 17191 24848
rect 15580 24790 17191 24792
rect 15580 24788 15586 24790
rect 17125 24787 17191 24790
rect 17309 24850 17375 24853
rect 22001 24850 22067 24853
rect 22185 24850 22251 24853
rect 17309 24848 22251 24850
rect 17309 24792 17314 24848
rect 17370 24792 22006 24848
rect 22062 24792 22190 24848
rect 22246 24792 22251 24848
rect 17309 24790 22251 24792
rect 23430 24850 23490 25062
rect 24393 25120 25839 25122
rect 24393 25064 24398 25120
rect 24454 25064 25778 25120
rect 25834 25064 25839 25120
rect 24393 25062 25839 25064
rect 24393 25059 24459 25062
rect 25773 25059 25839 25062
rect 26550 25060 26556 25124
rect 26620 25122 26626 25124
rect 26693 25122 26759 25125
rect 26620 25120 26759 25122
rect 26620 25064 26698 25120
rect 26754 25064 26759 25120
rect 26620 25062 26759 25064
rect 26620 25060 26626 25062
rect 26693 25059 26759 25062
rect 26969 25122 27035 25125
rect 30925 25122 30991 25125
rect 26969 25120 30991 25122
rect 26969 25064 26974 25120
rect 27030 25064 30930 25120
rect 30986 25064 30991 25120
rect 26969 25062 30991 25064
rect 26969 25059 27035 25062
rect 30925 25059 30991 25062
rect 23992 25056 24308 25057
rect 23992 24992 23998 25056
rect 24062 24992 24078 25056
rect 24142 24992 24158 25056
rect 24222 24992 24238 25056
rect 24302 24992 24308 25056
rect 23992 24991 24308 24992
rect 31674 25056 31990 25057
rect 31674 24992 31680 25056
rect 31744 24992 31760 25056
rect 31824 24992 31840 25056
rect 31904 24992 31920 25056
rect 31984 24992 31990 25056
rect 31674 24991 31990 24992
rect 23565 24988 23631 24989
rect 23565 24984 23612 24988
rect 23676 24986 23682 24988
rect 24393 24986 24459 24989
rect 25078 24986 25084 24988
rect 23565 24928 23570 24984
rect 23565 24924 23612 24928
rect 23676 24926 23722 24986
rect 24393 24984 25084 24986
rect 24393 24928 24398 24984
rect 24454 24928 25084 24984
rect 24393 24926 25084 24928
rect 23676 24924 23682 24926
rect 23565 24923 23631 24924
rect 24393 24923 24459 24926
rect 25078 24924 25084 24926
rect 25148 24924 25154 24988
rect 26417 24986 26483 24989
rect 31109 24988 31175 24989
rect 29862 24986 29868 24988
rect 26417 24984 29868 24986
rect 26417 24928 26422 24984
rect 26478 24928 29868 24984
rect 26417 24926 29868 24928
rect 26417 24923 26483 24926
rect 29824 24924 29868 24926
rect 29932 24986 29938 24988
rect 29932 24926 30014 24986
rect 31109 24984 31156 24988
rect 31220 24986 31226 24988
rect 31109 24928 31114 24984
rect 29932 24924 29938 24926
rect 31109 24924 31156 24928
rect 31220 24926 31266 24986
rect 31220 24924 31226 24926
rect 29824 24853 29884 24924
rect 31109 24923 31175 24924
rect 32206 24896 33006 25016
rect 25957 24850 26023 24853
rect 26366 24850 26372 24852
rect 23430 24790 24962 24850
rect 17309 24787 17375 24790
rect 22001 24787 22067 24790
rect 22185 24787 22251 24790
rect 5993 24714 6059 24717
rect 6862 24714 6868 24716
rect 5993 24712 6868 24714
rect 5993 24656 5998 24712
rect 6054 24656 6868 24712
rect 5993 24654 6868 24656
rect 5993 24651 6059 24654
rect 6862 24652 6868 24654
rect 6932 24714 6938 24716
rect 14774 24714 14780 24716
rect 6932 24654 14780 24714
rect 6932 24652 6938 24654
rect 14774 24652 14780 24654
rect 14844 24652 14850 24716
rect 15377 24714 15443 24717
rect 15510 24714 15516 24716
rect 15377 24712 15516 24714
rect 15377 24656 15382 24712
rect 15438 24656 15516 24712
rect 15377 24654 15516 24656
rect 15377 24651 15443 24654
rect 15510 24652 15516 24654
rect 15580 24652 15586 24716
rect 15929 24714 15995 24717
rect 16062 24714 16068 24716
rect 15929 24712 16068 24714
rect 15929 24656 15934 24712
rect 15990 24656 16068 24712
rect 15929 24654 16068 24656
rect 15929 24651 15995 24654
rect 16062 24652 16068 24654
rect 16132 24652 16138 24716
rect 16389 24714 16455 24717
rect 16849 24714 16915 24717
rect 16389 24712 16915 24714
rect 16389 24656 16394 24712
rect 16450 24656 16854 24712
rect 16910 24656 16915 24712
rect 16389 24654 16915 24656
rect 16389 24651 16455 24654
rect 16849 24651 16915 24654
rect 17350 24652 17356 24716
rect 17420 24714 17426 24716
rect 17493 24714 17559 24717
rect 17420 24712 17559 24714
rect 17420 24656 17498 24712
rect 17554 24656 17559 24712
rect 17420 24654 17559 24656
rect 17420 24652 17426 24654
rect 17493 24651 17559 24654
rect 17953 24714 18019 24717
rect 24761 24714 24827 24717
rect 17953 24712 24827 24714
rect 17953 24656 17958 24712
rect 18014 24656 24766 24712
rect 24822 24656 24827 24712
rect 17953 24654 24827 24656
rect 24902 24714 24962 24790
rect 25957 24848 26372 24850
rect 25957 24792 25962 24848
rect 26018 24792 26372 24848
rect 25957 24790 26372 24792
rect 25957 24787 26023 24790
rect 26366 24788 26372 24790
rect 26436 24788 26442 24852
rect 26734 24788 26740 24852
rect 26804 24850 26810 24852
rect 27429 24850 27495 24853
rect 29085 24852 29151 24853
rect 29085 24850 29132 24852
rect 26804 24848 27495 24850
rect 26804 24792 27434 24848
rect 27490 24792 27495 24848
rect 26804 24790 27495 24792
rect 26804 24788 26810 24790
rect 27429 24787 27495 24790
rect 27570 24790 28412 24850
rect 29040 24848 29132 24850
rect 29040 24792 29090 24848
rect 29040 24790 29132 24792
rect 25865 24714 25931 24717
rect 27570 24714 27630 24790
rect 28352 24714 28412 24790
rect 29085 24788 29132 24790
rect 29196 24788 29202 24852
rect 29821 24848 29887 24853
rect 29821 24792 29826 24848
rect 29882 24792 29887 24848
rect 29085 24787 29151 24788
rect 29821 24787 29887 24792
rect 30925 24714 30991 24717
rect 24902 24712 27630 24714
rect 24902 24656 25870 24712
rect 25926 24656 27630 24712
rect 24902 24654 27630 24656
rect 27708 24654 28274 24714
rect 28352 24712 30991 24714
rect 28352 24656 30930 24712
rect 30986 24656 30991 24712
rect 28352 24654 30991 24656
rect 17953 24651 18019 24654
rect 24761 24651 24827 24654
rect 25865 24651 25931 24654
rect 13854 24516 13860 24580
rect 13924 24578 13930 24580
rect 14825 24578 14891 24581
rect 15377 24580 15443 24581
rect 15326 24578 15332 24580
rect 13924 24576 14891 24578
rect 13924 24520 14830 24576
rect 14886 24520 14891 24576
rect 13924 24518 14891 24520
rect 15250 24518 15332 24578
rect 15396 24578 15443 24580
rect 18597 24578 18663 24581
rect 15396 24576 18663 24578
rect 15438 24520 18602 24576
rect 18658 24520 18663 24576
rect 13924 24516 13930 24518
rect 14825 24515 14891 24518
rect 15326 24516 15332 24518
rect 15396 24518 18663 24520
rect 15396 24516 15443 24518
rect 15377 24515 15443 24516
rect 18597 24515 18663 24518
rect 18873 24578 18939 24581
rect 19425 24578 19491 24581
rect 18873 24576 19491 24578
rect 18873 24520 18878 24576
rect 18934 24520 19430 24576
rect 19486 24520 19491 24576
rect 18873 24518 19491 24520
rect 18873 24515 18939 24518
rect 19425 24515 19491 24518
rect 19609 24578 19675 24581
rect 19885 24578 19951 24581
rect 25037 24578 25103 24581
rect 19609 24576 19951 24578
rect 19609 24520 19614 24576
rect 19670 24520 19890 24576
rect 19946 24520 19951 24576
rect 19609 24518 19951 24520
rect 19609 24515 19675 24518
rect 19885 24515 19951 24518
rect 20670 24576 25103 24578
rect 20670 24520 25042 24576
rect 25098 24520 25103 24576
rect 20670 24518 25103 24520
rect 4787 24512 5103 24513
rect 0 24352 800 24472
rect 4787 24448 4793 24512
rect 4857 24448 4873 24512
rect 4937 24448 4953 24512
rect 5017 24448 5033 24512
rect 5097 24448 5103 24512
rect 4787 24447 5103 24448
rect 12469 24512 12785 24513
rect 12469 24448 12475 24512
rect 12539 24448 12555 24512
rect 12619 24448 12635 24512
rect 12699 24448 12715 24512
rect 12779 24448 12785 24512
rect 12469 24447 12785 24448
rect 20151 24512 20467 24513
rect 20151 24448 20157 24512
rect 20221 24448 20237 24512
rect 20301 24448 20317 24512
rect 20381 24448 20397 24512
rect 20461 24448 20467 24512
rect 20151 24447 20467 24448
rect 14038 24380 14044 24444
rect 14108 24442 14114 24444
rect 14733 24442 14799 24445
rect 14108 24440 14799 24442
rect 14108 24384 14738 24440
rect 14794 24384 14799 24440
rect 14108 24382 14799 24384
rect 14108 24380 14114 24382
rect 14733 24379 14799 24382
rect 15561 24442 15627 24445
rect 16798 24442 16804 24444
rect 15561 24440 16804 24442
rect 15561 24384 15566 24440
rect 15622 24384 16804 24440
rect 15561 24382 16804 24384
rect 15561 24379 15627 24382
rect 16798 24380 16804 24382
rect 16868 24380 16874 24444
rect 17401 24442 17467 24445
rect 19517 24444 19583 24445
rect 19006 24442 19012 24444
rect 17401 24440 19012 24442
rect 17401 24384 17406 24440
rect 17462 24384 19012 24440
rect 17401 24382 19012 24384
rect 17401 24379 17467 24382
rect 19006 24380 19012 24382
rect 19076 24442 19082 24444
rect 19076 24382 19212 24442
rect 19076 24380 19082 24382
rect 6913 24306 6979 24309
rect 7046 24306 7052 24308
rect 6913 24304 7052 24306
rect 6913 24248 6918 24304
rect 6974 24248 7052 24304
rect 6913 24246 7052 24248
rect 6913 24243 6979 24246
rect 7046 24244 7052 24246
rect 7116 24244 7122 24308
rect 12157 24306 12223 24309
rect 7238 24304 12223 24306
rect 7238 24248 12162 24304
rect 12218 24248 12223 24304
rect 7238 24246 12223 24248
rect 5809 24170 5875 24173
rect 7238 24170 7298 24246
rect 12157 24243 12223 24246
rect 12433 24306 12499 24309
rect 13261 24306 13327 24309
rect 12433 24304 13327 24306
rect 12433 24248 12438 24304
rect 12494 24248 13266 24304
rect 13322 24248 13327 24304
rect 12433 24246 13327 24248
rect 12433 24243 12499 24246
rect 13261 24243 13327 24246
rect 14089 24306 14155 24309
rect 15326 24306 15332 24308
rect 14089 24304 15332 24306
rect 14089 24248 14094 24304
rect 14150 24248 15332 24304
rect 14089 24246 15332 24248
rect 14089 24243 14155 24246
rect 15326 24244 15332 24246
rect 15396 24244 15402 24308
rect 15745 24306 15811 24309
rect 16573 24306 16639 24309
rect 15745 24304 16639 24306
rect 15745 24248 15750 24304
rect 15806 24248 16578 24304
rect 16634 24248 16639 24304
rect 15745 24246 16639 24248
rect 15745 24243 15811 24246
rect 16573 24243 16639 24246
rect 16849 24306 16915 24309
rect 17493 24306 17559 24309
rect 18137 24306 18203 24309
rect 16849 24304 18203 24306
rect 16849 24248 16854 24304
rect 16910 24248 17498 24304
rect 17554 24248 18142 24304
rect 18198 24248 18203 24304
rect 16849 24246 18203 24248
rect 16849 24243 16915 24246
rect 17493 24243 17559 24246
rect 18137 24243 18203 24246
rect 18413 24306 18479 24309
rect 18873 24306 18939 24309
rect 18413 24304 18939 24306
rect 18413 24248 18418 24304
rect 18474 24248 18878 24304
rect 18934 24248 18939 24304
rect 18413 24246 18939 24248
rect 19152 24306 19212 24382
rect 19517 24440 19564 24444
rect 19628 24442 19634 24444
rect 19793 24442 19859 24445
rect 19977 24442 20043 24445
rect 19517 24384 19522 24440
rect 19517 24380 19564 24384
rect 19628 24382 19674 24442
rect 19793 24440 20043 24442
rect 19793 24384 19798 24440
rect 19854 24384 19982 24440
rect 20038 24384 20043 24440
rect 19793 24382 20043 24384
rect 19628 24380 19634 24382
rect 19517 24379 19583 24380
rect 19793 24379 19859 24382
rect 19977 24379 20043 24382
rect 20670 24306 20730 24518
rect 25037 24515 25103 24518
rect 25221 24578 25287 24581
rect 26693 24578 26759 24581
rect 26969 24578 27035 24581
rect 25221 24576 26204 24578
rect 25221 24520 25226 24576
rect 25282 24520 26204 24576
rect 25221 24518 26204 24520
rect 25221 24515 25287 24518
rect 20989 24442 21055 24445
rect 21541 24444 21607 24445
rect 21398 24442 21404 24444
rect 20989 24440 21404 24442
rect 20989 24384 20994 24440
rect 21050 24384 21404 24440
rect 20989 24382 21404 24384
rect 20989 24379 21055 24382
rect 21398 24380 21404 24382
rect 21468 24380 21474 24444
rect 21541 24440 21588 24444
rect 21652 24442 21658 24444
rect 22185 24442 22251 24445
rect 22369 24442 22435 24445
rect 23473 24442 23539 24445
rect 25589 24442 25655 24445
rect 25865 24444 25931 24445
rect 21541 24384 21546 24440
rect 21541 24380 21588 24384
rect 21652 24382 21698 24442
rect 22185 24440 23122 24442
rect 22185 24384 22190 24440
rect 22246 24384 22374 24440
rect 22430 24384 23122 24440
rect 22185 24382 23122 24384
rect 21652 24380 21658 24382
rect 21541 24379 21607 24380
rect 22185 24379 22251 24382
rect 22369 24379 22435 24382
rect 19152 24246 20730 24306
rect 21081 24306 21147 24309
rect 22870 24306 22876 24308
rect 21081 24304 22876 24306
rect 21081 24248 21086 24304
rect 21142 24248 22876 24304
rect 21081 24246 22876 24248
rect 18413 24243 18479 24246
rect 18873 24243 18939 24246
rect 21081 24243 21147 24246
rect 22870 24244 22876 24246
rect 22940 24244 22946 24308
rect 23062 24306 23122 24382
rect 23473 24440 25655 24442
rect 23473 24384 23478 24440
rect 23534 24384 25594 24440
rect 25650 24384 25655 24440
rect 23473 24382 25655 24384
rect 23473 24379 23539 24382
rect 25589 24379 25655 24382
rect 25814 24380 25820 24444
rect 25884 24442 25931 24444
rect 26144 24442 26204 24518
rect 26693 24576 27035 24578
rect 26693 24520 26698 24576
rect 26754 24520 26974 24576
rect 27030 24520 27035 24576
rect 26693 24518 27035 24520
rect 26693 24515 26759 24518
rect 26969 24515 27035 24518
rect 27102 24516 27108 24580
rect 27172 24578 27178 24580
rect 27708 24578 27768 24654
rect 27172 24518 27768 24578
rect 28214 24578 28274 24654
rect 30925 24651 30991 24654
rect 31477 24714 31543 24717
rect 32254 24714 32260 24716
rect 31477 24712 32260 24714
rect 31477 24656 31482 24712
rect 31538 24656 32260 24712
rect 31477 24654 32260 24656
rect 31477 24651 31543 24654
rect 32254 24652 32260 24654
rect 32324 24652 32330 24716
rect 30833 24578 30899 24581
rect 28214 24576 30899 24578
rect 28214 24520 30838 24576
rect 30894 24520 30899 24576
rect 28214 24518 30899 24520
rect 27172 24516 27178 24518
rect 30833 24515 30899 24518
rect 27833 24512 28149 24513
rect 27833 24448 27839 24512
rect 27903 24448 27919 24512
rect 27983 24448 27999 24512
rect 28063 24448 28079 24512
rect 28143 24448 28149 24512
rect 27833 24447 28149 24448
rect 28993 24442 29059 24445
rect 29862 24442 29868 24444
rect 25884 24440 25976 24442
rect 25926 24384 25976 24440
rect 25884 24382 25976 24384
rect 26144 24382 27170 24442
rect 25884 24380 25931 24382
rect 25865 24379 25931 24380
rect 27110 24306 27170 24382
rect 28993 24440 29868 24442
rect 28993 24384 28998 24440
rect 29054 24384 29868 24440
rect 28993 24382 29868 24384
rect 28993 24379 29059 24382
rect 29862 24380 29868 24382
rect 29932 24380 29938 24444
rect 32029 24442 32095 24445
rect 30192 24440 32095 24442
rect 30192 24384 32034 24440
rect 32090 24384 32095 24440
rect 30192 24382 32095 24384
rect 29821 24306 29887 24309
rect 30046 24306 30052 24308
rect 23062 24246 26986 24306
rect 27110 24246 29194 24306
rect 5809 24168 7298 24170
rect 5809 24112 5814 24168
rect 5870 24112 7298 24168
rect 5809 24110 7298 24112
rect 11421 24170 11487 24173
rect 13537 24170 13603 24173
rect 13905 24172 13971 24173
rect 11421 24168 13603 24170
rect 11421 24112 11426 24168
rect 11482 24112 13542 24168
rect 13598 24112 13603 24168
rect 11421 24110 13603 24112
rect 5809 24107 5875 24110
rect 11421 24107 11487 24110
rect 13537 24107 13603 24110
rect 13854 24108 13860 24172
rect 13924 24170 13971 24172
rect 14641 24170 14707 24173
rect 20989 24170 21055 24173
rect 21766 24170 21772 24172
rect 13924 24168 14016 24170
rect 13966 24112 14016 24168
rect 13924 24110 14016 24112
rect 14641 24168 21055 24170
rect 14641 24112 14646 24168
rect 14702 24112 20994 24168
rect 21050 24112 21055 24168
rect 14641 24110 21055 24112
rect 13924 24108 13971 24110
rect 13905 24107 13971 24108
rect 14641 24107 14707 24110
rect 20989 24107 21055 24110
rect 21176 24110 21772 24170
rect 13997 24034 14063 24037
rect 13997 24032 14796 24034
rect 13997 23976 14002 24032
rect 14058 23976 14796 24032
rect 13997 23974 14796 23976
rect 13997 23971 14063 23974
rect 8628 23968 8944 23969
rect 8628 23904 8634 23968
rect 8698 23904 8714 23968
rect 8778 23904 8794 23968
rect 8858 23904 8874 23968
rect 8938 23904 8944 23968
rect 8628 23903 8944 23904
rect 11881 23898 11947 23901
rect 14549 23898 14615 23901
rect 11881 23896 14615 23898
rect 11881 23840 11886 23896
rect 11942 23840 14554 23896
rect 14610 23840 14615 23896
rect 11881 23838 14615 23840
rect 14736 23898 14796 23974
rect 15142 23972 15148 24036
rect 15212 24034 15218 24036
rect 16113 24034 16179 24037
rect 15212 24032 16179 24034
rect 15212 23976 16118 24032
rect 16174 23976 16179 24032
rect 15212 23974 16179 23976
rect 15212 23972 15218 23974
rect 16113 23971 16179 23974
rect 16757 24036 16823 24037
rect 16757 24032 16804 24036
rect 16868 24034 16874 24036
rect 16757 23976 16762 24032
rect 16757 23972 16804 23976
rect 16868 23974 16914 24034
rect 16868 23972 16874 23974
rect 17534 23972 17540 24036
rect 17604 24034 17610 24036
rect 17953 24034 18019 24037
rect 17604 24032 18019 24034
rect 17604 23976 17958 24032
rect 18014 23976 18019 24032
rect 17604 23974 18019 23976
rect 17604 23972 17610 23974
rect 16757 23971 16823 23972
rect 17953 23971 18019 23974
rect 18137 24034 18203 24037
rect 19057 24034 19123 24037
rect 21176 24034 21236 24110
rect 21766 24108 21772 24110
rect 21836 24108 21842 24172
rect 22461 24170 22527 24173
rect 22686 24170 22692 24172
rect 22461 24168 22692 24170
rect 22461 24112 22466 24168
rect 22522 24112 22692 24168
rect 22461 24110 22692 24112
rect 22461 24107 22527 24110
rect 22686 24108 22692 24110
rect 22756 24108 22762 24172
rect 22921 24170 22987 24173
rect 25681 24170 25747 24173
rect 26785 24170 26851 24173
rect 22921 24168 26851 24170
rect 22921 24112 22926 24168
rect 22982 24112 25686 24168
rect 25742 24112 26790 24168
rect 26846 24112 26851 24168
rect 22921 24110 26851 24112
rect 26926 24170 26986 24246
rect 28993 24170 29059 24173
rect 26926 24168 29059 24170
rect 26926 24112 28998 24168
rect 29054 24112 29059 24168
rect 26926 24110 29059 24112
rect 29134 24170 29194 24246
rect 29821 24304 30052 24306
rect 29821 24248 29826 24304
rect 29882 24248 30052 24304
rect 29821 24246 30052 24248
rect 29821 24243 29887 24246
rect 30046 24244 30052 24246
rect 30116 24244 30122 24308
rect 29269 24170 29335 24173
rect 30192 24170 30252 24382
rect 32029 24379 32095 24382
rect 31569 24306 31635 24309
rect 32206 24306 33006 24336
rect 31569 24304 33006 24306
rect 31569 24248 31574 24304
rect 31630 24248 33006 24304
rect 31569 24246 33006 24248
rect 31569 24243 31635 24246
rect 32206 24216 33006 24246
rect 29134 24168 30252 24170
rect 29134 24112 29274 24168
rect 29330 24112 30252 24168
rect 29134 24110 30252 24112
rect 22921 24107 22987 24110
rect 25681 24107 25747 24110
rect 26785 24107 26851 24110
rect 28993 24107 29059 24110
rect 29269 24107 29335 24110
rect 18137 24032 21236 24034
rect 18137 23976 18142 24032
rect 18198 23976 19062 24032
rect 19118 23976 21236 24032
rect 18137 23974 21236 23976
rect 21449 24034 21515 24037
rect 22645 24034 22711 24037
rect 21449 24032 22711 24034
rect 21449 23976 21454 24032
rect 21510 23976 22650 24032
rect 22706 23976 22711 24032
rect 21449 23974 22711 23976
rect 18137 23971 18203 23974
rect 19057 23971 19123 23974
rect 21449 23971 21515 23974
rect 22645 23971 22711 23974
rect 22829 24034 22895 24037
rect 23381 24034 23447 24037
rect 23841 24034 23907 24037
rect 22829 24032 23907 24034
rect 22829 23976 22834 24032
rect 22890 23976 23386 24032
rect 23442 23976 23846 24032
rect 23902 23976 23907 24032
rect 22829 23974 23907 23976
rect 22829 23971 22895 23974
rect 23381 23971 23447 23974
rect 23841 23971 23907 23974
rect 25497 24034 25563 24037
rect 27245 24034 27311 24037
rect 25497 24032 27311 24034
rect 25497 23976 25502 24032
rect 25558 23976 27250 24032
rect 27306 23976 27311 24032
rect 25497 23974 27311 23976
rect 25497 23971 25563 23974
rect 27245 23971 27311 23974
rect 27470 23972 27476 24036
rect 27540 24034 27546 24036
rect 30833 24034 30899 24037
rect 27540 24032 30899 24034
rect 27540 23976 30838 24032
rect 30894 23976 30899 24032
rect 27540 23974 30899 23976
rect 27540 23972 27546 23974
rect 30833 23971 30899 23974
rect 16310 23968 16626 23969
rect 16310 23904 16316 23968
rect 16380 23904 16396 23968
rect 16460 23904 16476 23968
rect 16540 23904 16556 23968
rect 16620 23904 16626 23968
rect 16310 23903 16626 23904
rect 23992 23968 24308 23969
rect 23992 23904 23998 23968
rect 24062 23904 24078 23968
rect 24142 23904 24158 23968
rect 24222 23904 24238 23968
rect 24302 23904 24308 23968
rect 23992 23903 24308 23904
rect 31674 23968 31990 23969
rect 31674 23904 31680 23968
rect 31744 23904 31760 23968
rect 31824 23904 31840 23968
rect 31904 23904 31920 23968
rect 31984 23904 31990 23968
rect 31674 23903 31990 23904
rect 15285 23898 15351 23901
rect 14736 23896 15351 23898
rect 14736 23840 15290 23896
rect 15346 23840 15351 23896
rect 14736 23838 15351 23840
rect 11881 23835 11947 23838
rect 14549 23835 14615 23838
rect 15285 23835 15351 23838
rect 17166 23836 17172 23900
rect 17236 23898 17242 23900
rect 17309 23898 17375 23901
rect 17585 23900 17651 23901
rect 17534 23898 17540 23900
rect 17236 23896 17375 23898
rect 17236 23840 17314 23896
rect 17370 23840 17375 23896
rect 17236 23838 17375 23840
rect 17494 23838 17540 23898
rect 17604 23896 17651 23900
rect 17646 23840 17651 23896
rect 17236 23836 17242 23838
rect 17309 23835 17375 23838
rect 17534 23836 17540 23838
rect 17604 23836 17651 23840
rect 17718 23836 17724 23900
rect 17788 23898 17794 23900
rect 18137 23898 18203 23901
rect 17788 23896 18203 23898
rect 17788 23840 18142 23896
rect 18198 23840 18203 23896
rect 17788 23838 18203 23840
rect 17788 23836 17794 23838
rect 17585 23835 17651 23836
rect 18137 23835 18203 23838
rect 18321 23898 18387 23901
rect 19701 23898 19767 23901
rect 22737 23898 22803 23901
rect 18321 23896 19626 23898
rect 18321 23840 18326 23896
rect 18382 23840 19626 23896
rect 18321 23838 19626 23840
rect 18321 23835 18387 23838
rect 9673 23762 9739 23765
rect 12065 23762 12131 23765
rect 12341 23762 12407 23765
rect 14590 23762 14596 23764
rect 9673 23760 14596 23762
rect 9673 23704 9678 23760
rect 9734 23704 12070 23760
rect 12126 23704 12346 23760
rect 12402 23704 14596 23760
rect 9673 23702 14596 23704
rect 9673 23699 9739 23702
rect 12065 23699 12131 23702
rect 12341 23699 12407 23702
rect 14590 23700 14596 23702
rect 14660 23700 14666 23764
rect 14917 23762 14983 23765
rect 15745 23762 15811 23765
rect 19241 23762 19307 23765
rect 14917 23760 19307 23762
rect 14917 23704 14922 23760
rect 14978 23704 15750 23760
rect 15806 23704 19246 23760
rect 19302 23704 19307 23760
rect 14917 23702 19307 23704
rect 19566 23762 19626 23838
rect 19701 23896 22803 23898
rect 19701 23840 19706 23896
rect 19762 23840 22742 23896
rect 22798 23840 22803 23896
rect 19701 23838 22803 23840
rect 19701 23835 19767 23838
rect 22737 23835 22803 23838
rect 23197 23898 23263 23901
rect 23565 23898 23631 23901
rect 23197 23896 23631 23898
rect 23197 23840 23202 23896
rect 23258 23840 23570 23896
rect 23626 23840 23631 23896
rect 23197 23838 23631 23840
rect 23197 23835 23263 23838
rect 23565 23835 23631 23838
rect 23749 23900 23815 23901
rect 23749 23896 23796 23900
rect 23860 23898 23866 23900
rect 24485 23898 24551 23901
rect 26601 23898 26667 23901
rect 23749 23840 23754 23896
rect 23749 23836 23796 23840
rect 23860 23838 23906 23898
rect 24485 23896 30252 23898
rect 24485 23840 24490 23896
rect 24546 23840 26606 23896
rect 26662 23840 30252 23896
rect 24485 23838 30252 23840
rect 23860 23836 23866 23838
rect 23749 23835 23815 23836
rect 24485 23835 24551 23838
rect 26601 23835 26667 23838
rect 30192 23765 30252 23838
rect 21449 23762 21515 23765
rect 19566 23760 21515 23762
rect 19566 23704 21454 23760
rect 21510 23704 21515 23760
rect 19566 23702 21515 23704
rect 14917 23699 14983 23702
rect 15745 23699 15811 23702
rect 19241 23699 19307 23702
rect 21449 23699 21515 23702
rect 22093 23762 22159 23765
rect 22502 23762 22508 23764
rect 22093 23760 22508 23762
rect 22093 23704 22098 23760
rect 22154 23704 22508 23760
rect 22093 23702 22508 23704
rect 22093 23699 22159 23702
rect 22502 23700 22508 23702
rect 22572 23700 22578 23764
rect 22737 23762 22803 23765
rect 25221 23762 25287 23765
rect 22737 23760 25287 23762
rect 22737 23704 22742 23760
rect 22798 23704 25226 23760
rect 25282 23704 25287 23760
rect 22737 23702 25287 23704
rect 22737 23699 22803 23702
rect 25221 23699 25287 23702
rect 25681 23762 25747 23765
rect 26693 23764 26759 23765
rect 26693 23762 26740 23764
rect 25681 23760 26740 23762
rect 25681 23704 25686 23760
rect 25742 23704 26698 23760
rect 25681 23702 26740 23704
rect 25681 23699 25747 23702
rect 26693 23700 26740 23702
rect 26804 23700 26810 23764
rect 26877 23762 26943 23765
rect 30005 23762 30071 23765
rect 26877 23760 30071 23762
rect 26877 23704 26882 23760
rect 26938 23704 30010 23760
rect 30066 23704 30071 23760
rect 26877 23702 30071 23704
rect 26693 23699 26759 23700
rect 26877 23699 26943 23702
rect 30005 23699 30071 23702
rect 30189 23760 30255 23765
rect 30189 23704 30194 23760
rect 30250 23704 30255 23760
rect 30189 23699 30255 23704
rect 0 23626 800 23656
rect 1577 23626 1643 23629
rect 0 23624 1643 23626
rect 0 23568 1582 23624
rect 1638 23568 1643 23624
rect 0 23566 1643 23568
rect 0 23536 800 23566
rect 1577 23563 1643 23566
rect 9765 23626 9831 23629
rect 12157 23626 12223 23629
rect 9765 23624 12223 23626
rect 9765 23568 9770 23624
rect 9826 23568 12162 23624
rect 12218 23568 12223 23624
rect 9765 23566 12223 23568
rect 9765 23563 9831 23566
rect 12157 23563 12223 23566
rect 12985 23626 13051 23629
rect 12985 23624 15440 23626
rect 12985 23568 12990 23624
rect 13046 23568 15440 23624
rect 12985 23566 15440 23568
rect 12985 23563 13051 23566
rect 6310 23428 6316 23492
rect 6380 23490 6386 23492
rect 6821 23490 6887 23493
rect 6380 23488 6887 23490
rect 6380 23432 6826 23488
rect 6882 23432 6887 23488
rect 6380 23430 6887 23432
rect 6380 23428 6386 23430
rect 6821 23427 6887 23430
rect 11605 23490 11671 23493
rect 12341 23490 12407 23493
rect 11605 23488 12407 23490
rect 11605 23432 11610 23488
rect 11666 23432 12346 23488
rect 12402 23432 12407 23488
rect 11605 23430 12407 23432
rect 11605 23427 11671 23430
rect 12341 23427 12407 23430
rect 13261 23490 13327 23493
rect 13486 23490 13492 23492
rect 13261 23488 13492 23490
rect 13261 23432 13266 23488
rect 13322 23432 13492 23488
rect 13261 23430 13492 23432
rect 13261 23427 13327 23430
rect 13486 23428 13492 23430
rect 13556 23428 13562 23492
rect 14917 23490 14983 23493
rect 14644 23488 14983 23490
rect 14644 23432 14922 23488
rect 14978 23432 14983 23488
rect 14644 23430 14983 23432
rect 15380 23490 15440 23566
rect 15510 23564 15516 23628
rect 15580 23626 15586 23628
rect 23473 23626 23539 23629
rect 25865 23626 25931 23629
rect 15580 23624 23539 23626
rect 15580 23568 23478 23624
rect 23534 23568 23539 23624
rect 15580 23566 23539 23568
rect 15580 23564 15586 23566
rect 23473 23563 23539 23566
rect 23614 23624 25931 23626
rect 23614 23568 25870 23624
rect 25926 23568 25931 23624
rect 23614 23566 25931 23568
rect 17534 23490 17540 23492
rect 15380 23430 17540 23490
rect 4787 23424 5103 23425
rect 4787 23360 4793 23424
rect 4857 23360 4873 23424
rect 4937 23360 4953 23424
rect 5017 23360 5033 23424
rect 5097 23360 5103 23424
rect 4787 23359 5103 23360
rect 12469 23424 12785 23425
rect 12469 23360 12475 23424
rect 12539 23360 12555 23424
rect 12619 23360 12635 23424
rect 12699 23360 12715 23424
rect 12779 23360 12785 23424
rect 12469 23359 12785 23360
rect 8477 23354 8543 23357
rect 9254 23354 9260 23356
rect 8477 23352 9260 23354
rect 8477 23296 8482 23352
rect 8538 23296 9260 23352
rect 8477 23294 9260 23296
rect 8477 23291 8543 23294
rect 9254 23292 9260 23294
rect 9324 23354 9330 23356
rect 11053 23354 11119 23357
rect 13353 23356 13419 23357
rect 13302 23354 13308 23356
rect 9324 23352 11119 23354
rect 9324 23296 11058 23352
rect 11114 23296 11119 23352
rect 9324 23294 11119 23296
rect 13262 23294 13308 23354
rect 13372 23352 13419 23356
rect 13414 23296 13419 23352
rect 9324 23292 9330 23294
rect 11053 23291 11119 23294
rect 13302 23292 13308 23294
rect 13372 23292 13419 23296
rect 13353 23291 13419 23292
rect 13537 23354 13603 23357
rect 13905 23354 13971 23357
rect 13537 23352 13971 23354
rect 13537 23296 13542 23352
rect 13598 23296 13910 23352
rect 13966 23296 13971 23352
rect 13537 23294 13971 23296
rect 13537 23291 13603 23294
rect 13905 23291 13971 23294
rect 14089 23354 14155 23357
rect 14644 23354 14704 23430
rect 14917 23427 14983 23430
rect 17534 23428 17540 23430
rect 17604 23428 17610 23492
rect 19425 23490 19491 23493
rect 19742 23490 19748 23492
rect 17680 23430 19258 23490
rect 14825 23356 14891 23357
rect 14089 23352 14704 23354
rect 14089 23296 14094 23352
rect 14150 23296 14704 23352
rect 14089 23294 14704 23296
rect 14089 23291 14155 23294
rect 14774 23292 14780 23356
rect 14844 23354 14891 23356
rect 14844 23352 14936 23354
rect 14886 23296 14936 23352
rect 14844 23294 14936 23296
rect 14844 23292 14891 23294
rect 15142 23292 15148 23356
rect 15212 23354 15218 23356
rect 16205 23354 16271 23357
rect 15212 23352 16271 23354
rect 15212 23296 16210 23352
rect 16266 23296 16271 23352
rect 15212 23294 16271 23296
rect 15212 23292 15218 23294
rect 14825 23291 14891 23292
rect 16205 23291 16271 23294
rect 16389 23354 16455 23357
rect 16982 23354 16988 23356
rect 16389 23352 16988 23354
rect 16389 23296 16394 23352
rect 16450 23296 16988 23352
rect 16389 23294 16988 23296
rect 16389 23291 16455 23294
rect 16982 23292 16988 23294
rect 17052 23292 17058 23356
rect 17125 23354 17191 23357
rect 17680 23354 17740 23430
rect 17125 23352 17740 23354
rect 17125 23296 17130 23352
rect 17186 23296 17740 23352
rect 17125 23294 17740 23296
rect 18321 23354 18387 23357
rect 19057 23354 19123 23357
rect 18321 23352 19123 23354
rect 18321 23296 18326 23352
rect 18382 23296 19062 23352
rect 19118 23296 19123 23352
rect 18321 23294 19123 23296
rect 19198 23354 19258 23430
rect 19425 23488 19748 23490
rect 19425 23432 19430 23488
rect 19486 23432 19748 23488
rect 19425 23430 19748 23432
rect 19425 23427 19491 23430
rect 19742 23428 19748 23430
rect 19812 23428 19818 23492
rect 20529 23488 20595 23493
rect 20529 23432 20534 23488
rect 20590 23432 20595 23488
rect 20529 23427 20595 23432
rect 20662 23428 20668 23492
rect 20732 23490 20738 23492
rect 21081 23490 21147 23493
rect 20732 23488 21147 23490
rect 20732 23432 21086 23488
rect 21142 23432 21147 23488
rect 20732 23430 21147 23432
rect 20732 23428 20738 23430
rect 21081 23427 21147 23430
rect 21357 23490 21423 23493
rect 23473 23490 23539 23493
rect 21357 23488 23539 23490
rect 21357 23432 21362 23488
rect 21418 23432 23478 23488
rect 23534 23432 23539 23488
rect 21357 23430 23539 23432
rect 21357 23427 21423 23430
rect 23473 23427 23539 23430
rect 20151 23424 20467 23425
rect 20151 23360 20157 23424
rect 20221 23360 20237 23424
rect 20301 23360 20317 23424
rect 20381 23360 20397 23424
rect 20461 23360 20467 23424
rect 20151 23359 20467 23360
rect 19701 23354 19767 23357
rect 19198 23352 19767 23354
rect 19198 23296 19706 23352
rect 19762 23296 19767 23352
rect 19198 23294 19767 23296
rect 20532 23354 20592 23427
rect 20662 23354 20668 23356
rect 20532 23294 20668 23354
rect 17125 23291 17191 23294
rect 18321 23291 18387 23294
rect 19057 23291 19123 23294
rect 19701 23291 19767 23294
rect 20662 23292 20668 23294
rect 20732 23292 20738 23356
rect 20846 23292 20852 23356
rect 20916 23354 20922 23356
rect 23614 23354 23674 23566
rect 25865 23563 25931 23566
rect 26325 23626 26391 23629
rect 27153 23626 27219 23629
rect 26325 23624 27219 23626
rect 26325 23568 26330 23624
rect 26386 23568 27158 23624
rect 27214 23568 27219 23624
rect 26325 23566 27219 23568
rect 26325 23563 26391 23566
rect 27153 23563 27219 23566
rect 27286 23564 27292 23628
rect 27356 23626 27362 23628
rect 29821 23626 29887 23629
rect 27356 23624 29887 23626
rect 27356 23568 29826 23624
rect 29882 23568 29887 23624
rect 27356 23566 29887 23568
rect 27356 23564 27362 23566
rect 29821 23563 29887 23566
rect 30281 23626 30347 23629
rect 32206 23626 33006 23656
rect 30281 23624 33006 23626
rect 30281 23568 30286 23624
rect 30342 23568 33006 23624
rect 30281 23566 33006 23568
rect 30281 23563 30347 23566
rect 32206 23536 33006 23566
rect 24526 23428 24532 23492
rect 24596 23490 24602 23492
rect 26509 23490 26575 23493
rect 24596 23488 26575 23490
rect 24596 23432 26514 23488
rect 26570 23432 26575 23488
rect 24596 23430 26575 23432
rect 24596 23428 24602 23430
rect 26509 23427 26575 23430
rect 26734 23428 26740 23492
rect 26804 23490 26810 23492
rect 27429 23490 27495 23493
rect 26804 23488 27495 23490
rect 26804 23432 27434 23488
rect 27490 23432 27495 23488
rect 26804 23430 27495 23432
rect 26804 23428 26810 23430
rect 27429 23427 27495 23430
rect 28390 23428 28396 23492
rect 28460 23490 28466 23492
rect 28533 23490 28599 23493
rect 28460 23488 28599 23490
rect 28460 23432 28538 23488
rect 28594 23432 28599 23488
rect 28460 23430 28599 23432
rect 28460 23428 28466 23430
rect 28533 23427 28599 23430
rect 28717 23490 28783 23493
rect 29085 23490 29151 23493
rect 28717 23488 29151 23490
rect 28717 23432 28722 23488
rect 28778 23432 29090 23488
rect 29146 23432 29151 23488
rect 28717 23430 29151 23432
rect 28717 23427 28783 23430
rect 29085 23427 29151 23430
rect 27833 23424 28149 23425
rect 27833 23360 27839 23424
rect 27903 23360 27919 23424
rect 27983 23360 27999 23424
rect 28063 23360 28079 23424
rect 28143 23360 28149 23424
rect 27833 23359 28149 23360
rect 20916 23294 23674 23354
rect 24393 23354 24459 23357
rect 27705 23356 27771 23357
rect 28441 23356 28507 23357
rect 28809 23356 28875 23357
rect 27102 23354 27108 23356
rect 24393 23352 27108 23354
rect 24393 23296 24398 23352
rect 24454 23296 27108 23352
rect 24393 23294 27108 23296
rect 20916 23292 20922 23294
rect 24393 23291 24459 23294
rect 27102 23292 27108 23294
rect 27172 23292 27178 23356
rect 27654 23354 27660 23356
rect 27614 23294 27660 23354
rect 27724 23352 27771 23356
rect 27766 23296 27771 23352
rect 27654 23292 27660 23294
rect 27724 23292 27771 23296
rect 28390 23292 28396 23356
rect 28460 23354 28507 23356
rect 28460 23352 28552 23354
rect 28502 23296 28552 23352
rect 28460 23294 28552 23296
rect 28460 23292 28507 23294
rect 28758 23292 28764 23356
rect 28828 23354 28875 23356
rect 30097 23354 30163 23357
rect 30230 23354 30236 23356
rect 28828 23352 28920 23354
rect 28870 23296 28920 23352
rect 28828 23294 28920 23296
rect 30097 23352 30236 23354
rect 30097 23296 30102 23352
rect 30158 23296 30236 23352
rect 30097 23294 30236 23296
rect 28828 23292 28875 23294
rect 27705 23291 27771 23292
rect 28441 23291 28507 23292
rect 28809 23291 28875 23292
rect 30097 23291 30163 23294
rect 30230 23292 30236 23294
rect 30300 23292 30306 23356
rect 31334 23292 31340 23356
rect 31404 23354 31410 23356
rect 32397 23354 32463 23357
rect 31404 23352 32463 23354
rect 31404 23296 32402 23352
rect 32458 23296 32463 23352
rect 31404 23294 32463 23296
rect 31404 23292 31410 23294
rect 32397 23291 32463 23294
rect 8845 23218 8911 23221
rect 12709 23218 12775 23221
rect 8845 23216 12775 23218
rect 8845 23160 8850 23216
rect 8906 23160 12714 23216
rect 12770 23160 12775 23216
rect 8845 23158 12775 23160
rect 8845 23155 8911 23158
rect 12709 23155 12775 23158
rect 13445 23218 13511 23221
rect 17769 23218 17835 23221
rect 13445 23216 17835 23218
rect 13445 23160 13450 23216
rect 13506 23160 17774 23216
rect 17830 23160 17835 23216
rect 13445 23158 17835 23160
rect 13445 23155 13511 23158
rect 17769 23155 17835 23158
rect 17902 23156 17908 23220
rect 17972 23218 17978 23220
rect 21817 23218 21883 23221
rect 17972 23216 21883 23218
rect 17972 23160 21822 23216
rect 21878 23160 21883 23216
rect 17972 23158 21883 23160
rect 17972 23156 17978 23158
rect 21817 23155 21883 23158
rect 22001 23218 22067 23221
rect 25405 23218 25471 23221
rect 22001 23216 25471 23218
rect 22001 23160 22006 23216
rect 22062 23160 25410 23216
rect 25466 23160 25471 23216
rect 22001 23158 25471 23160
rect 22001 23155 22067 23158
rect 25405 23155 25471 23158
rect 25589 23218 25655 23221
rect 31017 23218 31083 23221
rect 25589 23216 31083 23218
rect 25589 23160 25594 23216
rect 25650 23160 31022 23216
rect 31078 23160 31083 23216
rect 25589 23158 31083 23160
rect 25589 23155 25655 23158
rect 31017 23155 31083 23158
rect 8201 23082 8267 23085
rect 12801 23082 12867 23085
rect 28625 23082 28691 23085
rect 8201 23080 12680 23082
rect 8201 23024 8206 23080
rect 8262 23024 12680 23080
rect 8201 23022 12680 23024
rect 8201 23019 8267 23022
rect 12620 22949 12680 23022
rect 12801 23080 28691 23082
rect 12801 23024 12806 23080
rect 12862 23024 28630 23080
rect 28686 23024 28691 23080
rect 12801 23022 28691 23024
rect 12801 23019 12867 23022
rect 28625 23019 28691 23022
rect 28809 23082 28875 23085
rect 29821 23082 29887 23085
rect 28809 23080 29887 23082
rect 28809 23024 28814 23080
rect 28870 23024 29826 23080
rect 29882 23024 29887 23080
rect 28809 23022 29887 23024
rect 28809 23019 28875 23022
rect 29821 23019 29887 23022
rect 11881 22946 11947 22949
rect 12157 22946 12223 22949
rect 11881 22944 12223 22946
rect 11881 22888 11886 22944
rect 11942 22888 12162 22944
rect 12218 22888 12223 22944
rect 11881 22886 12223 22888
rect 11881 22883 11947 22886
rect 12157 22883 12223 22886
rect 12617 22946 12683 22949
rect 13486 22946 13492 22948
rect 12617 22944 13492 22946
rect 12617 22888 12622 22944
rect 12678 22888 13492 22944
rect 12617 22886 13492 22888
rect 12617 22883 12683 22886
rect 13486 22884 13492 22886
rect 13556 22884 13562 22948
rect 13721 22946 13787 22949
rect 16021 22946 16087 22949
rect 17401 22946 17467 22949
rect 17769 22948 17835 22949
rect 13721 22944 16087 22946
rect 13721 22888 13726 22944
rect 13782 22888 16026 22944
rect 16082 22888 16087 22944
rect 13721 22886 16087 22888
rect 13721 22883 13787 22886
rect 16021 22883 16087 22886
rect 16760 22944 17467 22946
rect 16760 22888 17406 22944
rect 17462 22888 17467 22944
rect 16760 22886 17467 22888
rect 8628 22880 8944 22881
rect 0 22810 800 22840
rect 8628 22816 8634 22880
rect 8698 22816 8714 22880
rect 8778 22816 8794 22880
rect 8858 22816 8874 22880
rect 8938 22816 8944 22880
rect 8628 22815 8944 22816
rect 16310 22880 16626 22881
rect 16310 22816 16316 22880
rect 16380 22816 16396 22880
rect 16460 22816 16476 22880
rect 16540 22816 16556 22880
rect 16620 22816 16626 22880
rect 16310 22815 16626 22816
rect 1577 22810 1643 22813
rect 8201 22812 8267 22813
rect 0 22808 1643 22810
rect 0 22752 1582 22808
rect 1638 22752 1643 22808
rect 0 22750 1643 22752
rect 0 22720 800 22750
rect 1577 22747 1643 22750
rect 8150 22748 8156 22812
rect 8220 22810 8267 22812
rect 11237 22810 11303 22813
rect 14641 22810 14707 22813
rect 15837 22810 15903 22813
rect 8220 22808 8312 22810
rect 8262 22752 8312 22808
rect 8220 22750 8312 22752
rect 11237 22808 14060 22810
rect 11237 22752 11242 22808
rect 11298 22752 14060 22808
rect 11237 22750 14060 22752
rect 8220 22748 8267 22750
rect 8201 22747 8267 22748
rect 11237 22747 11303 22750
rect 10501 22674 10567 22677
rect 11421 22676 11487 22677
rect 11421 22674 11468 22676
rect 10501 22672 11468 22674
rect 10501 22616 10506 22672
rect 10562 22616 11426 22672
rect 10501 22614 11468 22616
rect 10501 22611 10567 22614
rect 11421 22612 11468 22614
rect 11532 22612 11538 22676
rect 11697 22674 11763 22677
rect 13854 22674 13860 22676
rect 11697 22672 13860 22674
rect 11697 22616 11702 22672
rect 11758 22616 13860 22672
rect 11697 22614 13860 22616
rect 11421 22611 11487 22612
rect 11697 22611 11763 22614
rect 13854 22612 13860 22614
rect 13924 22612 13930 22676
rect 14000 22674 14060 22750
rect 14641 22808 15903 22810
rect 14641 22752 14646 22808
rect 14702 22752 15842 22808
rect 15898 22752 15903 22808
rect 14641 22750 15903 22752
rect 14641 22747 14707 22750
rect 15837 22747 15903 22750
rect 16760 22674 16820 22886
rect 17401 22883 17467 22886
rect 17718 22884 17724 22948
rect 17788 22946 17835 22948
rect 17788 22944 17880 22946
rect 17830 22888 17880 22944
rect 17788 22886 17880 22888
rect 17788 22884 17835 22886
rect 18270 22884 18276 22948
rect 18340 22946 18346 22948
rect 18413 22946 18479 22949
rect 18340 22944 18479 22946
rect 18340 22888 18418 22944
rect 18474 22888 18479 22944
rect 18340 22886 18479 22888
rect 18340 22884 18346 22886
rect 17769 22883 17835 22884
rect 18413 22883 18479 22886
rect 18638 22884 18644 22948
rect 18708 22946 18714 22948
rect 22001 22946 22067 22949
rect 18708 22944 22067 22946
rect 18708 22888 22006 22944
rect 22062 22888 22067 22944
rect 18708 22886 22067 22888
rect 18708 22884 18714 22886
rect 22001 22883 22067 22886
rect 22369 22946 22435 22949
rect 23606 22946 23612 22948
rect 22369 22944 23612 22946
rect 22369 22888 22374 22944
rect 22430 22888 23612 22944
rect 22369 22886 23612 22888
rect 22369 22883 22435 22886
rect 23606 22884 23612 22886
rect 23676 22884 23682 22948
rect 24577 22946 24643 22949
rect 27153 22946 27219 22949
rect 29637 22946 29703 22949
rect 24577 22944 29703 22946
rect 24577 22888 24582 22944
rect 24638 22888 27158 22944
rect 27214 22888 29642 22944
rect 29698 22888 29703 22944
rect 24577 22886 29703 22888
rect 24577 22883 24643 22886
rect 27153 22883 27219 22886
rect 29637 22883 29703 22886
rect 23992 22880 24308 22881
rect 23992 22816 23998 22880
rect 24062 22816 24078 22880
rect 24142 22816 24158 22880
rect 24222 22816 24238 22880
rect 24302 22816 24308 22880
rect 23992 22815 24308 22816
rect 31674 22880 31990 22881
rect 31674 22816 31680 22880
rect 31744 22816 31760 22880
rect 31824 22816 31840 22880
rect 31904 22816 31920 22880
rect 31984 22816 31990 22880
rect 32206 22856 33006 22976
rect 31674 22815 31990 22816
rect 17166 22748 17172 22812
rect 17236 22810 17242 22812
rect 17309 22810 17375 22813
rect 17236 22808 17375 22810
rect 17236 22752 17314 22808
rect 17370 22752 17375 22808
rect 17236 22750 17375 22752
rect 17236 22748 17242 22750
rect 17309 22747 17375 22750
rect 17861 22810 17927 22813
rect 18413 22810 18479 22813
rect 19333 22810 19399 22813
rect 23422 22810 23428 22812
rect 17861 22808 18479 22810
rect 17861 22752 17866 22808
rect 17922 22752 18418 22808
rect 18474 22752 18479 22808
rect 17861 22750 18479 22752
rect 17861 22747 17927 22750
rect 18413 22747 18479 22750
rect 18876 22750 19212 22810
rect 14000 22614 16820 22674
rect 16982 22612 16988 22676
rect 17052 22674 17058 22676
rect 17217 22674 17283 22677
rect 17052 22672 17283 22674
rect 17052 22616 17222 22672
rect 17278 22616 17283 22672
rect 17052 22614 17283 22616
rect 17052 22612 17058 22614
rect 17217 22611 17283 22614
rect 17718 22612 17724 22676
rect 17788 22674 17794 22676
rect 18876 22674 18936 22750
rect 17788 22614 18936 22674
rect 19152 22674 19212 22750
rect 19333 22808 23428 22810
rect 19333 22752 19338 22808
rect 19394 22752 23428 22808
rect 19333 22750 23428 22752
rect 19333 22747 19399 22750
rect 23422 22748 23428 22750
rect 23492 22748 23498 22812
rect 24710 22748 24716 22812
rect 24780 22810 24786 22812
rect 28073 22810 28139 22813
rect 24780 22808 28139 22810
rect 24780 22752 28078 22808
rect 28134 22752 28139 22808
rect 24780 22750 28139 22752
rect 24780 22748 24786 22750
rect 28073 22747 28139 22750
rect 28257 22810 28323 22813
rect 29729 22810 29795 22813
rect 29862 22810 29868 22812
rect 28257 22808 29868 22810
rect 28257 22752 28262 22808
rect 28318 22752 29734 22808
rect 29790 22752 29868 22808
rect 28257 22750 29868 22752
rect 28257 22747 28323 22750
rect 29729 22747 29795 22750
rect 29862 22748 29868 22750
rect 29932 22748 29938 22812
rect 30230 22748 30236 22812
rect 30300 22810 30306 22812
rect 31293 22810 31359 22813
rect 30300 22808 31359 22810
rect 30300 22752 31298 22808
rect 31354 22752 31359 22808
rect 30300 22750 31359 22752
rect 30300 22748 30306 22750
rect 31293 22747 31359 22750
rect 21030 22674 21036 22676
rect 19152 22614 21036 22674
rect 17788 22612 17794 22614
rect 21030 22612 21036 22614
rect 21100 22674 21106 22676
rect 21265 22674 21331 22677
rect 21100 22672 21331 22674
rect 21100 22616 21270 22672
rect 21326 22616 21331 22672
rect 21100 22614 21331 22616
rect 21100 22612 21106 22614
rect 21265 22611 21331 22614
rect 21398 22612 21404 22676
rect 21468 22674 21474 22676
rect 21633 22674 21699 22677
rect 22737 22674 22803 22677
rect 31293 22674 31359 22677
rect 21468 22672 21699 22674
rect 21468 22616 21638 22672
rect 21694 22616 21699 22672
rect 21468 22614 21699 22616
rect 21468 22612 21474 22614
rect 21633 22611 21699 22614
rect 21774 22672 22803 22674
rect 21774 22616 22742 22672
rect 22798 22616 22803 22672
rect 21774 22614 22803 22616
rect 10593 22538 10659 22541
rect 13445 22538 13511 22541
rect 18270 22538 18276 22540
rect 10593 22536 18276 22538
rect 10593 22480 10598 22536
rect 10654 22480 13450 22536
rect 13506 22480 18276 22536
rect 10593 22478 18276 22480
rect 10593 22475 10659 22478
rect 13445 22475 13511 22478
rect 18270 22476 18276 22478
rect 18340 22476 18346 22540
rect 19701 22538 19767 22541
rect 20897 22538 20963 22541
rect 19701 22536 20963 22538
rect 19701 22480 19706 22536
rect 19762 22480 20902 22536
rect 20958 22480 20963 22536
rect 19701 22478 20963 22480
rect 19701 22475 19767 22478
rect 20897 22475 20963 22478
rect 21030 22476 21036 22540
rect 21100 22538 21106 22540
rect 21582 22538 21588 22540
rect 21100 22478 21588 22538
rect 21100 22476 21106 22478
rect 21582 22476 21588 22478
rect 21652 22476 21658 22540
rect 8201 22402 8267 22405
rect 12157 22402 12223 22405
rect 8201 22400 12223 22402
rect 8201 22344 8206 22400
rect 8262 22344 12162 22400
rect 12218 22344 12223 22400
rect 8201 22342 12223 22344
rect 8201 22339 8267 22342
rect 12157 22339 12223 22342
rect 13261 22404 13327 22405
rect 13261 22400 13308 22404
rect 13372 22402 13378 22404
rect 15837 22402 15903 22405
rect 18597 22402 18663 22405
rect 19793 22402 19859 22405
rect 13261 22344 13266 22400
rect 13261 22340 13308 22344
rect 13372 22342 13418 22402
rect 15837 22400 19859 22402
rect 15837 22344 15842 22400
rect 15898 22344 18602 22400
rect 18658 22344 19798 22400
rect 19854 22344 19859 22400
rect 15837 22342 19859 22344
rect 13372 22340 13378 22342
rect 13261 22339 13327 22340
rect 15837 22339 15903 22342
rect 18597 22339 18663 22342
rect 19793 22339 19859 22342
rect 20805 22402 20871 22405
rect 21774 22402 21834 22614
rect 22737 22611 22803 22614
rect 22878 22672 31359 22674
rect 22878 22616 31298 22672
rect 31354 22616 31359 22672
rect 22878 22614 31359 22616
rect 21950 22476 21956 22540
rect 22020 22538 22026 22540
rect 22878 22538 22938 22614
rect 31293 22611 31359 22614
rect 22020 22478 22938 22538
rect 23473 22538 23539 22541
rect 26366 22538 26372 22540
rect 23473 22536 26372 22538
rect 23473 22480 23478 22536
rect 23534 22480 26372 22536
rect 23473 22478 26372 22480
rect 22020 22476 22026 22478
rect 23473 22475 23539 22478
rect 26366 22476 26372 22478
rect 26436 22476 26442 22540
rect 26601 22538 26667 22541
rect 27245 22538 27311 22541
rect 27521 22540 27587 22541
rect 27470 22538 27476 22540
rect 26601 22536 27311 22538
rect 26601 22480 26606 22536
rect 26662 22480 27250 22536
rect 27306 22480 27311 22536
rect 26601 22478 27311 22480
rect 27430 22478 27476 22538
rect 27540 22536 27587 22540
rect 27582 22480 27587 22536
rect 26601 22475 26667 22478
rect 27245 22475 27311 22478
rect 27470 22476 27476 22478
rect 27540 22476 27587 22480
rect 27654 22476 27660 22540
rect 27724 22538 27730 22540
rect 28441 22538 28507 22541
rect 27724 22536 28507 22538
rect 27724 22480 28446 22536
rect 28502 22480 28507 22536
rect 27724 22478 28507 22480
rect 27724 22476 27730 22478
rect 27521 22475 27587 22476
rect 28441 22475 28507 22478
rect 20805 22400 21834 22402
rect 20805 22344 20810 22400
rect 20866 22344 21834 22400
rect 20805 22342 21834 22344
rect 20805 22339 20871 22342
rect 22134 22340 22140 22404
rect 22204 22402 22210 22404
rect 22921 22402 22987 22405
rect 22204 22400 22987 22402
rect 22204 22344 22926 22400
rect 22982 22344 22987 22400
rect 22204 22342 22987 22344
rect 22204 22340 22210 22342
rect 22921 22339 22987 22342
rect 23105 22402 23171 22405
rect 25078 22402 25084 22404
rect 23105 22400 25084 22402
rect 23105 22344 23110 22400
rect 23166 22344 25084 22400
rect 23105 22342 25084 22344
rect 23105 22339 23171 22342
rect 25078 22340 25084 22342
rect 25148 22340 25154 22404
rect 25221 22402 25287 22405
rect 27613 22402 27679 22405
rect 25221 22400 27679 22402
rect 25221 22344 25226 22400
rect 25282 22344 27618 22400
rect 27674 22344 27679 22400
rect 25221 22342 27679 22344
rect 25221 22339 25287 22342
rect 27613 22339 27679 22342
rect 28349 22402 28415 22405
rect 30925 22402 30991 22405
rect 28349 22400 30991 22402
rect 28349 22344 28354 22400
rect 28410 22344 30930 22400
rect 30986 22344 30991 22400
rect 28349 22342 30991 22344
rect 28349 22339 28415 22342
rect 30925 22339 30991 22342
rect 4787 22336 5103 22337
rect 4787 22272 4793 22336
rect 4857 22272 4873 22336
rect 4937 22272 4953 22336
rect 5017 22272 5033 22336
rect 5097 22272 5103 22336
rect 4787 22271 5103 22272
rect 12469 22336 12785 22337
rect 12469 22272 12475 22336
rect 12539 22272 12555 22336
rect 12619 22272 12635 22336
rect 12699 22272 12715 22336
rect 12779 22272 12785 22336
rect 12469 22271 12785 22272
rect 20151 22336 20467 22337
rect 20151 22272 20157 22336
rect 20221 22272 20237 22336
rect 20301 22272 20317 22336
rect 20381 22272 20397 22336
rect 20461 22272 20467 22336
rect 20151 22271 20467 22272
rect 27833 22336 28149 22337
rect 27833 22272 27839 22336
rect 27903 22272 27919 22336
rect 27983 22272 27999 22336
rect 28063 22272 28079 22336
rect 28143 22272 28149 22336
rect 27833 22271 28149 22272
rect 11973 22268 12039 22269
rect 11973 22266 12020 22268
rect 11928 22264 12020 22266
rect 11928 22208 11978 22264
rect 11928 22206 12020 22208
rect 11973 22204 12020 22206
rect 12084 22204 12090 22268
rect 12893 22266 12959 22269
rect 13721 22266 13787 22269
rect 12893 22264 13787 22266
rect 12893 22208 12898 22264
rect 12954 22208 13726 22264
rect 13782 22208 13787 22264
rect 12893 22206 13787 22208
rect 11973 22203 12039 22204
rect 12893 22203 12959 22206
rect 13721 22203 13787 22206
rect 13854 22204 13860 22268
rect 13924 22266 13930 22268
rect 16665 22266 16731 22269
rect 13924 22264 16731 22266
rect 13924 22208 16670 22264
rect 16726 22208 16731 22264
rect 13924 22206 16731 22208
rect 13924 22204 13930 22206
rect 16665 22203 16731 22206
rect 16798 22204 16804 22268
rect 16868 22266 16874 22268
rect 16941 22266 17007 22269
rect 16868 22264 17007 22266
rect 16868 22208 16946 22264
rect 17002 22208 17007 22264
rect 16868 22206 17007 22208
rect 16868 22204 16874 22206
rect 16941 22203 17007 22206
rect 17677 22266 17743 22269
rect 18638 22266 18644 22268
rect 17677 22264 18644 22266
rect 17677 22208 17682 22264
rect 17738 22208 18644 22264
rect 17677 22206 18644 22208
rect 17677 22203 17743 22206
rect 18638 22204 18644 22206
rect 18708 22204 18714 22268
rect 18781 22266 18847 22269
rect 19374 22266 19380 22268
rect 18781 22264 19380 22266
rect 18781 22208 18786 22264
rect 18842 22208 19380 22264
rect 18781 22206 19380 22208
rect 18781 22203 18847 22206
rect 19374 22204 19380 22206
rect 19444 22266 19450 22268
rect 19977 22266 20043 22269
rect 19444 22264 20043 22266
rect 19444 22208 19982 22264
rect 20038 22208 20043 22264
rect 19444 22206 20043 22208
rect 19444 22204 19450 22206
rect 19977 22203 20043 22206
rect 20662 22204 20668 22268
rect 20732 22266 20738 22268
rect 23933 22266 23999 22269
rect 28349 22268 28415 22269
rect 20732 22264 23999 22266
rect 20732 22208 23938 22264
rect 23994 22208 23999 22264
rect 20732 22206 23999 22208
rect 20732 22204 20738 22206
rect 23933 22203 23999 22206
rect 24902 22206 27538 22266
rect 7833 22130 7899 22133
rect 11145 22130 11211 22133
rect 12801 22130 12867 22133
rect 14365 22130 14431 22133
rect 17217 22130 17283 22133
rect 18413 22130 18479 22133
rect 7790 22128 12220 22130
rect 7790 22072 7838 22128
rect 7894 22072 11150 22128
rect 11206 22072 12220 22128
rect 7790 22070 12220 22072
rect 7790 22067 7899 22070
rect 11145 22067 11211 22070
rect 0 21904 800 22024
rect 4705 21994 4771 21997
rect 7790 21994 7850 22067
rect 4705 21992 7850 21994
rect 4705 21936 4710 21992
rect 4766 21936 7850 21992
rect 4705 21934 7850 21936
rect 8753 21994 8819 21997
rect 10174 21994 10180 21996
rect 8753 21992 10180 21994
rect 8753 21936 8758 21992
rect 8814 21936 10180 21992
rect 8753 21934 10180 21936
rect 4705 21931 4771 21934
rect 8753 21931 8819 21934
rect 10174 21932 10180 21934
rect 10244 21932 10250 21996
rect 12160 21994 12220 22070
rect 12801 22128 17050 22130
rect 12801 22072 12806 22128
rect 12862 22072 14370 22128
rect 14426 22072 17050 22128
rect 12801 22070 17050 22072
rect 12801 22067 12867 22070
rect 14365 22067 14431 22070
rect 15285 21994 15351 21997
rect 12160 21992 16912 21994
rect 12160 21936 15290 21992
rect 15346 21936 16912 21992
rect 12160 21934 16912 21936
rect 15285 21931 15351 21934
rect 6729 21858 6795 21861
rect 6862 21858 6868 21860
rect 6729 21856 6868 21858
rect 6729 21800 6734 21856
rect 6790 21800 6868 21856
rect 6729 21798 6868 21800
rect 6729 21795 6795 21798
rect 6862 21796 6868 21798
rect 6932 21796 6938 21860
rect 9029 21858 9095 21861
rect 12617 21858 12683 21861
rect 13118 21858 13124 21860
rect 9029 21856 13124 21858
rect 9029 21800 9034 21856
rect 9090 21800 12622 21856
rect 12678 21800 13124 21856
rect 9029 21798 13124 21800
rect 9029 21795 9095 21798
rect 12617 21795 12683 21798
rect 13118 21796 13124 21798
rect 13188 21858 13194 21860
rect 14641 21858 14707 21861
rect 13188 21856 14707 21858
rect 13188 21800 14646 21856
rect 14702 21800 14707 21856
rect 13188 21798 14707 21800
rect 13188 21796 13194 21798
rect 14641 21795 14707 21798
rect 15469 21858 15535 21861
rect 15878 21858 15884 21860
rect 15469 21856 15884 21858
rect 15469 21800 15474 21856
rect 15530 21800 15884 21856
rect 15469 21798 15884 21800
rect 15469 21795 15535 21798
rect 15878 21796 15884 21798
rect 15948 21858 15954 21860
rect 16113 21858 16179 21861
rect 15948 21856 16179 21858
rect 15948 21800 16118 21856
rect 16174 21800 16179 21856
rect 15948 21798 16179 21800
rect 15948 21796 15954 21798
rect 16113 21795 16179 21798
rect 8628 21792 8944 21793
rect 8628 21728 8634 21792
rect 8698 21728 8714 21792
rect 8778 21728 8794 21792
rect 8858 21728 8874 21792
rect 8938 21728 8944 21792
rect 8628 21727 8944 21728
rect 16310 21792 16626 21793
rect 16310 21728 16316 21792
rect 16380 21728 16396 21792
rect 16460 21728 16476 21792
rect 16540 21728 16556 21792
rect 16620 21728 16626 21792
rect 16310 21727 16626 21728
rect 12249 21724 12315 21725
rect 12198 21722 12204 21724
rect 12158 21662 12204 21722
rect 12268 21720 12315 21724
rect 12310 21664 12315 21720
rect 12198 21660 12204 21662
rect 12268 21660 12315 21664
rect 12249 21659 12315 21660
rect 12433 21722 12499 21725
rect 14181 21724 14247 21725
rect 14181 21722 14228 21724
rect 12433 21720 13554 21722
rect 12433 21664 12438 21720
rect 12494 21664 13554 21720
rect 12433 21662 13554 21664
rect 14100 21720 14228 21722
rect 14292 21722 14298 21724
rect 16113 21722 16179 21725
rect 14292 21720 16179 21722
rect 14100 21664 14186 21720
rect 14292 21664 16118 21720
rect 16174 21664 16179 21720
rect 14100 21662 14228 21664
rect 12433 21659 12499 21662
rect 9765 21586 9831 21589
rect 13353 21586 13419 21589
rect 9765 21584 13419 21586
rect 9765 21528 9770 21584
rect 9826 21528 13358 21584
rect 13414 21528 13419 21584
rect 9765 21526 13419 21528
rect 13494 21586 13554 21662
rect 14181 21660 14228 21662
rect 14292 21662 16179 21664
rect 16852 21722 16912 21934
rect 16990 21858 17050 22070
rect 17217 22128 18479 22130
rect 17217 22072 17222 22128
rect 17278 22072 18418 22128
rect 18474 22072 18479 22128
rect 17217 22070 18479 22072
rect 17217 22067 17283 22070
rect 18413 22067 18479 22070
rect 18638 22068 18644 22132
rect 18708 22130 18714 22132
rect 21357 22130 21423 22133
rect 18708 22128 21423 22130
rect 18708 22072 21362 22128
rect 21418 22072 21423 22128
rect 18708 22070 21423 22072
rect 18708 22068 18714 22070
rect 21357 22067 21423 22070
rect 22001 22130 22067 22133
rect 24902 22130 24962 22206
rect 22001 22128 24962 22130
rect 22001 22072 22006 22128
rect 22062 22072 24962 22128
rect 22001 22070 24962 22072
rect 25313 22130 25379 22133
rect 26141 22132 26207 22133
rect 25630 22130 25636 22132
rect 25313 22128 25636 22130
rect 25313 22072 25318 22128
rect 25374 22072 25636 22128
rect 25313 22070 25636 22072
rect 22001 22067 22067 22070
rect 25313 22067 25379 22070
rect 25630 22068 25636 22070
rect 25700 22068 25706 22132
rect 26141 22130 26188 22132
rect 26096 22128 26188 22130
rect 26096 22072 26146 22128
rect 26096 22070 26188 22072
rect 26141 22068 26188 22070
rect 26252 22068 26258 22132
rect 26366 22068 26372 22132
rect 26436 22130 26442 22132
rect 26969 22130 27035 22133
rect 26436 22128 27035 22130
rect 26436 22072 26974 22128
rect 27030 22072 27035 22128
rect 26436 22070 27035 22072
rect 27478 22130 27538 22206
rect 28349 22264 28396 22268
rect 28460 22266 28466 22268
rect 28349 22208 28354 22264
rect 28349 22204 28396 22208
rect 28460 22206 28506 22266
rect 28460 22204 28466 22206
rect 28942 22204 28948 22268
rect 29012 22266 29018 22268
rect 32206 22266 33006 22296
rect 29012 22206 33006 22266
rect 29012 22204 29018 22206
rect 28349 22203 28415 22204
rect 32206 22176 33006 22206
rect 30005 22130 30071 22133
rect 27478 22128 30071 22130
rect 27478 22072 30010 22128
rect 30066 22072 30071 22128
rect 27478 22070 30071 22072
rect 26436 22068 26442 22070
rect 26141 22067 26207 22068
rect 26969 22067 27035 22070
rect 30005 22067 30071 22070
rect 17125 21994 17191 21997
rect 17677 21994 17743 21997
rect 17953 21996 18019 21997
rect 17902 21994 17908 21996
rect 17125 21992 17743 21994
rect 17125 21936 17130 21992
rect 17186 21936 17682 21992
rect 17738 21936 17743 21992
rect 17125 21934 17743 21936
rect 17862 21934 17908 21994
rect 17972 21992 18019 21996
rect 30281 21994 30347 21997
rect 18014 21936 18019 21992
rect 17125 21931 17191 21934
rect 17677 21931 17743 21934
rect 17902 21932 17908 21934
rect 17972 21932 18019 21936
rect 17953 21931 18019 21932
rect 18416 21992 30347 21994
rect 18416 21936 30286 21992
rect 30342 21936 30347 21992
rect 18416 21934 30347 21936
rect 17718 21858 17724 21860
rect 16990 21798 17724 21858
rect 17718 21796 17724 21798
rect 17788 21796 17794 21860
rect 18045 21858 18111 21861
rect 18416 21858 18476 21934
rect 30281 21931 30347 21934
rect 30649 21994 30715 21997
rect 30966 21994 30972 21996
rect 30649 21992 30972 21994
rect 30649 21936 30654 21992
rect 30710 21936 30972 21992
rect 30649 21934 30972 21936
rect 30649 21931 30715 21934
rect 30966 21932 30972 21934
rect 31036 21932 31042 21996
rect 18045 21856 18476 21858
rect 18045 21800 18050 21856
rect 18106 21800 18476 21856
rect 18045 21798 18476 21800
rect 18045 21795 18111 21798
rect 18822 21796 18828 21860
rect 18892 21858 18898 21860
rect 21633 21858 21699 21861
rect 18892 21856 21699 21858
rect 18892 21800 21638 21856
rect 21694 21800 21699 21856
rect 18892 21798 21699 21800
rect 18892 21796 18898 21798
rect 21633 21795 21699 21798
rect 21766 21796 21772 21860
rect 21836 21858 21842 21860
rect 22686 21858 22692 21860
rect 21836 21798 22692 21858
rect 21836 21796 21842 21798
rect 22686 21796 22692 21798
rect 22756 21796 22762 21860
rect 24669 21858 24735 21861
rect 26550 21858 26556 21860
rect 24669 21856 26556 21858
rect 24669 21800 24674 21856
rect 24730 21800 26556 21856
rect 24669 21798 26556 21800
rect 24669 21795 24735 21798
rect 26550 21796 26556 21798
rect 26620 21796 26626 21860
rect 28993 21858 29059 21861
rect 26742 21856 29059 21858
rect 26742 21800 28998 21856
rect 29054 21800 29059 21856
rect 26742 21798 29059 21800
rect 23992 21792 24308 21793
rect 23992 21728 23998 21792
rect 24062 21728 24078 21792
rect 24142 21728 24158 21792
rect 24222 21728 24238 21792
rect 24302 21728 24308 21792
rect 23992 21727 24308 21728
rect 17350 21722 17356 21724
rect 16852 21662 17356 21722
rect 14292 21660 14298 21662
rect 14181 21659 14247 21660
rect 16113 21659 16179 21662
rect 17350 21660 17356 21662
rect 17420 21660 17426 21724
rect 18086 21660 18092 21724
rect 18156 21722 18162 21724
rect 18229 21722 18295 21725
rect 18505 21724 18571 21725
rect 18156 21720 18295 21722
rect 18156 21664 18234 21720
rect 18290 21664 18295 21720
rect 18156 21662 18295 21664
rect 18156 21660 18162 21662
rect 18229 21659 18295 21662
rect 18454 21660 18460 21724
rect 18524 21722 18571 21724
rect 18689 21722 18755 21725
rect 18873 21722 18939 21725
rect 18524 21720 18616 21722
rect 18566 21664 18616 21720
rect 18524 21662 18616 21664
rect 18689 21720 18939 21722
rect 18689 21664 18694 21720
rect 18750 21664 18878 21720
rect 18934 21664 18939 21720
rect 18689 21662 18939 21664
rect 18524 21660 18571 21662
rect 18505 21659 18571 21660
rect 18689 21659 18755 21662
rect 18873 21659 18939 21662
rect 19057 21722 19123 21725
rect 19374 21722 19380 21724
rect 19057 21720 19380 21722
rect 19057 21664 19062 21720
rect 19118 21664 19380 21720
rect 19057 21662 19380 21664
rect 19057 21659 19123 21662
rect 19374 21660 19380 21662
rect 19444 21660 19450 21724
rect 19609 21722 19675 21725
rect 22185 21722 22251 21725
rect 19609 21720 22251 21722
rect 19609 21664 19614 21720
rect 19670 21664 22190 21720
rect 22246 21664 22251 21720
rect 19609 21662 22251 21664
rect 19609 21659 19675 21662
rect 22185 21659 22251 21662
rect 24577 21722 24643 21725
rect 26742 21722 26802 21798
rect 28993 21795 29059 21798
rect 29126 21796 29132 21860
rect 29196 21858 29202 21860
rect 29545 21858 29611 21861
rect 29196 21856 29611 21858
rect 29196 21800 29550 21856
rect 29606 21800 29611 21856
rect 29196 21798 29611 21800
rect 29196 21796 29202 21798
rect 29545 21795 29611 21798
rect 29913 21858 29979 21861
rect 30966 21858 30972 21860
rect 29913 21856 30972 21858
rect 29913 21800 29918 21856
rect 29974 21800 30972 21856
rect 29913 21798 30972 21800
rect 29913 21795 29979 21798
rect 30966 21796 30972 21798
rect 31036 21796 31042 21860
rect 31674 21792 31990 21793
rect 31674 21728 31680 21792
rect 31744 21728 31760 21792
rect 31824 21728 31840 21792
rect 31904 21728 31920 21792
rect 31984 21728 31990 21792
rect 31674 21727 31990 21728
rect 24577 21720 26802 21722
rect 24577 21664 24582 21720
rect 24638 21664 26802 21720
rect 24577 21662 26802 21664
rect 26969 21722 27035 21725
rect 29729 21722 29795 21725
rect 26969 21720 29795 21722
rect 26969 21664 26974 21720
rect 27030 21664 29734 21720
rect 29790 21664 29795 21720
rect 26969 21662 29795 21664
rect 24577 21659 24643 21662
rect 26969 21659 27035 21662
rect 29729 21659 29795 21662
rect 29913 21722 29979 21725
rect 30414 21722 30420 21724
rect 29913 21720 30420 21722
rect 29913 21664 29918 21720
rect 29974 21664 30420 21720
rect 29913 21662 30420 21664
rect 29913 21659 29979 21662
rect 30414 21660 30420 21662
rect 30484 21660 30490 21724
rect 31150 21660 31156 21724
rect 31220 21722 31226 21724
rect 31220 21662 31402 21722
rect 31220 21660 31226 21662
rect 14457 21586 14523 21589
rect 13494 21584 14523 21586
rect 13494 21528 14462 21584
rect 14518 21528 14523 21584
rect 13494 21526 14523 21528
rect 9765 21523 9831 21526
rect 13353 21523 13419 21526
rect 14457 21523 14523 21526
rect 15285 21586 15351 21589
rect 17166 21586 17172 21588
rect 15285 21584 17172 21586
rect 15285 21528 15290 21584
rect 15346 21528 17172 21584
rect 15285 21526 17172 21528
rect 15285 21523 15351 21526
rect 17166 21524 17172 21526
rect 17236 21524 17242 21588
rect 17309 21586 17375 21589
rect 17534 21586 17540 21588
rect 17309 21584 17540 21586
rect 17309 21528 17314 21584
rect 17370 21528 17540 21584
rect 17309 21526 17540 21528
rect 17309 21523 17375 21526
rect 17534 21524 17540 21526
rect 17604 21524 17610 21588
rect 17769 21586 17835 21589
rect 31109 21586 31175 21589
rect 17769 21584 31175 21586
rect 17769 21528 17774 21584
rect 17830 21528 31114 21584
rect 31170 21528 31175 21584
rect 17769 21526 31175 21528
rect 31342 21586 31402 21662
rect 32206 21586 33006 21616
rect 31342 21526 33006 21586
rect 17769 21523 17835 21526
rect 31109 21523 31175 21526
rect 32206 21496 33006 21526
rect 9673 21450 9739 21453
rect 12341 21450 12407 21453
rect 9673 21448 12407 21450
rect 9673 21392 9678 21448
rect 9734 21392 12346 21448
rect 12402 21392 12407 21448
rect 9673 21390 12407 21392
rect 9673 21387 9739 21390
rect 12341 21387 12407 21390
rect 12525 21450 12591 21453
rect 12934 21450 12940 21452
rect 12525 21448 12940 21450
rect 12525 21392 12530 21448
rect 12586 21392 12940 21448
rect 12525 21390 12940 21392
rect 12525 21387 12591 21390
rect 12934 21388 12940 21390
rect 13004 21388 13010 21452
rect 14733 21450 14799 21453
rect 17534 21450 17540 21452
rect 14733 21448 17540 21450
rect 14733 21392 14738 21448
rect 14794 21392 17540 21448
rect 14733 21390 17540 21392
rect 14733 21387 14799 21390
rect 17534 21388 17540 21390
rect 17604 21388 17610 21452
rect 17861 21450 17927 21453
rect 28809 21450 28875 21453
rect 17861 21448 28875 21450
rect 17861 21392 17866 21448
rect 17922 21392 28814 21448
rect 28870 21392 28875 21448
rect 17861 21390 28875 21392
rect 17861 21387 17927 21390
rect 28809 21387 28875 21390
rect 28993 21450 29059 21453
rect 30833 21452 30899 21453
rect 30598 21450 30604 21452
rect 28993 21448 30604 21450
rect 28993 21392 28998 21448
rect 29054 21392 30604 21448
rect 28993 21390 30604 21392
rect 28993 21387 29059 21390
rect 30598 21388 30604 21390
rect 30668 21388 30674 21452
rect 30782 21388 30788 21452
rect 30852 21450 30899 21452
rect 30852 21448 30944 21450
rect 30894 21392 30944 21448
rect 30852 21390 30944 21392
rect 30852 21388 30899 21390
rect 30833 21387 30899 21388
rect 13302 21252 13308 21316
rect 13372 21314 13378 21316
rect 19977 21314 20043 21317
rect 13372 21312 20043 21314
rect 13372 21256 19982 21312
rect 20038 21256 20043 21312
rect 13372 21254 20043 21256
rect 13372 21252 13378 21254
rect 19977 21251 20043 21254
rect 20529 21314 20595 21317
rect 21081 21314 21147 21317
rect 20529 21312 21147 21314
rect 20529 21256 20534 21312
rect 20590 21256 21086 21312
rect 21142 21256 21147 21312
rect 20529 21254 21147 21256
rect 20529 21251 20595 21254
rect 21081 21251 21147 21254
rect 21817 21314 21883 21317
rect 23565 21314 23631 21317
rect 21817 21312 23631 21314
rect 21817 21256 21822 21312
rect 21878 21256 23570 21312
rect 23626 21256 23631 21312
rect 21817 21254 23631 21256
rect 21817 21251 21883 21254
rect 23565 21251 23631 21254
rect 24485 21314 24551 21317
rect 26417 21314 26483 21317
rect 24485 21312 26483 21314
rect 24485 21256 24490 21312
rect 24546 21256 26422 21312
rect 26478 21256 26483 21312
rect 24485 21254 26483 21256
rect 24485 21251 24551 21254
rect 26417 21251 26483 21254
rect 26550 21252 26556 21316
rect 26620 21314 26626 21316
rect 27613 21314 27679 21317
rect 26620 21312 27679 21314
rect 26620 21256 27618 21312
rect 27674 21256 27679 21312
rect 26620 21254 27679 21256
rect 26620 21252 26626 21254
rect 27613 21251 27679 21254
rect 28993 21314 29059 21317
rect 30833 21314 30899 21317
rect 28993 21312 30899 21314
rect 28993 21256 28998 21312
rect 29054 21256 30838 21312
rect 30894 21256 30899 21312
rect 28993 21254 30899 21256
rect 28993 21251 29059 21254
rect 30833 21251 30899 21254
rect 4787 21248 5103 21249
rect 0 21178 800 21208
rect 4787 21184 4793 21248
rect 4857 21184 4873 21248
rect 4937 21184 4953 21248
rect 5017 21184 5033 21248
rect 5097 21184 5103 21248
rect 4787 21183 5103 21184
rect 12469 21248 12785 21249
rect 12469 21184 12475 21248
rect 12539 21184 12555 21248
rect 12619 21184 12635 21248
rect 12699 21184 12715 21248
rect 12779 21184 12785 21248
rect 12469 21183 12785 21184
rect 20151 21248 20467 21249
rect 20151 21184 20157 21248
rect 20221 21184 20237 21248
rect 20301 21184 20317 21248
rect 20381 21184 20397 21248
rect 20461 21184 20467 21248
rect 20151 21183 20467 21184
rect 27833 21248 28149 21249
rect 27833 21184 27839 21248
rect 27903 21184 27919 21248
rect 27983 21184 27999 21248
rect 28063 21184 28079 21248
rect 28143 21184 28149 21248
rect 27833 21183 28149 21184
rect 1577 21178 1643 21181
rect 0 21176 1643 21178
rect 0 21120 1582 21176
rect 1638 21120 1643 21176
rect 0 21118 1643 21120
rect 0 21088 800 21118
rect 1577 21115 1643 21118
rect 7741 21178 7807 21181
rect 12014 21178 12020 21180
rect 7741 21176 12020 21178
rect 7741 21120 7746 21176
rect 7802 21120 12020 21176
rect 7741 21118 12020 21120
rect 7741 21115 7807 21118
rect 12014 21116 12020 21118
rect 12084 21178 12090 21180
rect 12341 21178 12407 21181
rect 12084 21176 12407 21178
rect 12084 21120 12346 21176
rect 12402 21120 12407 21176
rect 12084 21118 12407 21120
rect 12084 21116 12090 21118
rect 12341 21115 12407 21118
rect 13629 21178 13695 21181
rect 16021 21178 16087 21181
rect 13629 21176 16087 21178
rect 13629 21120 13634 21176
rect 13690 21120 16026 21176
rect 16082 21120 16087 21176
rect 13629 21118 16087 21120
rect 13629 21115 13695 21118
rect 16021 21115 16087 21118
rect 16389 21178 16455 21181
rect 16982 21178 16988 21180
rect 16389 21176 16988 21178
rect 16389 21120 16394 21176
rect 16450 21120 16988 21176
rect 16389 21118 16988 21120
rect 16389 21115 16455 21118
rect 16982 21116 16988 21118
rect 17052 21178 17058 21180
rect 19558 21178 19564 21180
rect 17052 21118 19564 21178
rect 17052 21116 17058 21118
rect 19558 21116 19564 21118
rect 19628 21116 19634 21180
rect 20662 21116 20668 21180
rect 20732 21178 20738 21180
rect 22185 21178 22251 21181
rect 20732 21176 22251 21178
rect 20732 21120 22190 21176
rect 22246 21120 22251 21176
rect 20732 21118 22251 21120
rect 20732 21116 20738 21118
rect 22185 21115 22251 21118
rect 22318 21116 22324 21180
rect 22388 21178 22394 21180
rect 28257 21178 28323 21181
rect 28390 21178 28396 21180
rect 22388 21118 27676 21178
rect 22388 21116 22394 21118
rect 8293 21042 8359 21045
rect 12065 21042 12131 21045
rect 16665 21042 16731 21045
rect 25221 21042 25287 21045
rect 8293 21040 11898 21042
rect 8293 20984 8298 21040
rect 8354 20984 11898 21040
rect 8293 20982 11898 20984
rect 8293 20979 8402 20982
rect 8342 20637 8402 20979
rect 11838 20906 11898 20982
rect 12065 21040 16590 21042
rect 12065 20984 12070 21040
rect 12126 20984 16590 21040
rect 12065 20982 16590 20984
rect 12065 20979 12131 20982
rect 12525 20906 12591 20909
rect 15009 20906 15075 20909
rect 11838 20904 12591 20906
rect 11838 20848 12530 20904
rect 12586 20848 12591 20904
rect 11838 20846 12591 20848
rect 12525 20843 12591 20846
rect 13126 20904 15075 20906
rect 13126 20848 15014 20904
rect 15070 20848 15075 20904
rect 13126 20846 15075 20848
rect 10869 20772 10935 20773
rect 10869 20768 10916 20772
rect 10980 20770 10986 20772
rect 11421 20770 11487 20773
rect 11646 20770 11652 20772
rect 10869 20712 10874 20768
rect 10869 20708 10916 20712
rect 10980 20710 11026 20770
rect 11421 20768 11652 20770
rect 11421 20712 11426 20768
rect 11482 20712 11652 20768
rect 11421 20710 11652 20712
rect 10980 20708 10986 20710
rect 10869 20707 10935 20708
rect 11421 20707 11487 20710
rect 11646 20708 11652 20710
rect 11716 20708 11722 20772
rect 12065 20770 12131 20773
rect 12198 20770 12204 20772
rect 12065 20768 12204 20770
rect 12065 20712 12070 20768
rect 12126 20712 12204 20768
rect 12065 20710 12204 20712
rect 12065 20707 12131 20710
rect 12198 20708 12204 20710
rect 12268 20708 12274 20772
rect 12341 20770 12407 20773
rect 13126 20770 13186 20846
rect 15009 20843 15075 20846
rect 15285 20906 15351 20909
rect 16297 20906 16363 20909
rect 15285 20904 16363 20906
rect 15285 20848 15290 20904
rect 15346 20848 16302 20904
rect 16358 20848 16363 20904
rect 15285 20846 16363 20848
rect 16530 20906 16590 20982
rect 16665 21040 25287 21042
rect 16665 20984 16670 21040
rect 16726 20984 25226 21040
rect 25282 20984 25287 21040
rect 16665 20982 25287 20984
rect 16665 20979 16731 20982
rect 25221 20979 25287 20982
rect 25773 21042 25839 21045
rect 26693 21042 26759 21045
rect 25773 21040 26759 21042
rect 25773 20984 25778 21040
rect 25834 20984 26698 21040
rect 26754 20984 26759 21040
rect 25773 20982 26759 20984
rect 25773 20979 25839 20982
rect 26693 20979 26759 20982
rect 26918 20980 26924 21044
rect 26988 21042 26994 21044
rect 27245 21042 27311 21045
rect 27429 21044 27495 21045
rect 27429 21042 27476 21044
rect 26988 21040 27311 21042
rect 26988 20984 27250 21040
rect 27306 20984 27311 21040
rect 26988 20982 27311 20984
rect 27384 21040 27476 21042
rect 27384 20984 27434 21040
rect 27384 20982 27476 20984
rect 26988 20980 26994 20982
rect 27245 20979 27311 20982
rect 27429 20980 27476 20982
rect 27540 20980 27546 21044
rect 27616 21042 27676 21118
rect 28257 21176 28396 21178
rect 28257 21120 28262 21176
rect 28318 21120 28396 21176
rect 28257 21118 28396 21120
rect 28257 21115 28323 21118
rect 28390 21116 28396 21118
rect 28460 21116 28466 21180
rect 28625 21178 28691 21181
rect 31109 21178 31175 21181
rect 28625 21176 31175 21178
rect 28625 21120 28630 21176
rect 28686 21120 31114 21176
rect 31170 21120 31175 21176
rect 28625 21118 31175 21120
rect 28625 21115 28691 21118
rect 31109 21115 31175 21118
rect 29637 21042 29703 21045
rect 27616 21040 29703 21042
rect 27616 20984 29642 21040
rect 29698 20984 29703 21040
rect 27616 20982 29703 20984
rect 27429 20979 27495 20980
rect 29637 20979 29703 20982
rect 29821 21042 29887 21045
rect 30046 21042 30052 21044
rect 29821 21040 30052 21042
rect 29821 20984 29826 21040
rect 29882 20984 30052 21040
rect 29821 20982 30052 20984
rect 29821 20979 29887 20982
rect 30046 20980 30052 20982
rect 30116 20980 30122 21044
rect 17309 20906 17375 20909
rect 16530 20904 17375 20906
rect 16530 20848 17314 20904
rect 17370 20848 17375 20904
rect 16530 20846 17375 20848
rect 15285 20843 15351 20846
rect 16297 20843 16363 20846
rect 17309 20843 17375 20846
rect 17534 20844 17540 20908
rect 17604 20906 17610 20908
rect 17677 20906 17743 20909
rect 20897 20906 20963 20909
rect 17604 20904 20963 20906
rect 17604 20848 17682 20904
rect 17738 20848 20902 20904
rect 20958 20848 20963 20904
rect 17604 20846 20963 20848
rect 17604 20844 17610 20846
rect 17677 20843 17743 20846
rect 20897 20843 20963 20846
rect 21633 20906 21699 20909
rect 29085 20906 29151 20909
rect 21633 20904 29151 20906
rect 21633 20848 21638 20904
rect 21694 20848 29090 20904
rect 29146 20848 29151 20904
rect 21633 20846 29151 20848
rect 21633 20843 21699 20846
rect 29085 20843 29151 20846
rect 29678 20844 29684 20908
rect 29748 20906 29754 20908
rect 30005 20906 30071 20909
rect 29748 20904 30071 20906
rect 29748 20848 30010 20904
rect 30066 20848 30071 20904
rect 29748 20846 30071 20848
rect 29748 20844 29754 20846
rect 30005 20843 30071 20846
rect 30189 20906 30255 20909
rect 30414 20906 30420 20908
rect 30189 20904 30420 20906
rect 30189 20848 30194 20904
rect 30250 20848 30420 20904
rect 30189 20846 30420 20848
rect 30189 20843 30255 20846
rect 30414 20844 30420 20846
rect 30484 20844 30490 20908
rect 31201 20906 31267 20909
rect 32206 20906 33006 20936
rect 31201 20904 33006 20906
rect 31201 20848 31206 20904
rect 31262 20848 33006 20904
rect 31201 20846 33006 20848
rect 31201 20843 31267 20846
rect 32206 20816 33006 20846
rect 12341 20768 13186 20770
rect 12341 20712 12346 20768
rect 12402 20712 13186 20768
rect 12341 20710 13186 20712
rect 13261 20770 13327 20773
rect 13445 20770 13511 20773
rect 15653 20770 15719 20773
rect 13261 20768 15719 20770
rect 13261 20712 13266 20768
rect 13322 20712 13450 20768
rect 13506 20712 15658 20768
rect 15714 20712 15719 20768
rect 13261 20710 15719 20712
rect 12341 20707 12407 20710
rect 13261 20707 13327 20710
rect 13445 20707 13511 20710
rect 15653 20707 15719 20710
rect 17166 20708 17172 20772
rect 17236 20770 17242 20772
rect 18137 20770 18203 20773
rect 22461 20770 22527 20773
rect 17236 20768 22527 20770
rect 17236 20712 18142 20768
rect 18198 20712 22466 20768
rect 22522 20712 22527 20768
rect 17236 20710 22527 20712
rect 17236 20708 17242 20710
rect 18137 20707 18203 20710
rect 22461 20707 22527 20710
rect 25078 20708 25084 20772
rect 25148 20770 25154 20772
rect 26233 20770 26299 20773
rect 25148 20768 26299 20770
rect 25148 20712 26238 20768
rect 26294 20712 26299 20768
rect 25148 20710 26299 20712
rect 25148 20708 25154 20710
rect 26233 20707 26299 20710
rect 26417 20770 26483 20773
rect 29453 20770 29519 20773
rect 26417 20768 29519 20770
rect 26417 20712 26422 20768
rect 26478 20712 29458 20768
rect 29514 20712 29519 20768
rect 26417 20710 29519 20712
rect 26417 20707 26483 20710
rect 29453 20707 29519 20710
rect 29637 20772 29703 20773
rect 29637 20768 29684 20772
rect 29748 20770 29754 20772
rect 29913 20770 29979 20773
rect 30373 20770 30439 20773
rect 29637 20712 29642 20768
rect 29637 20708 29684 20712
rect 29748 20710 29794 20770
rect 29913 20768 30439 20770
rect 29913 20712 29918 20768
rect 29974 20712 30378 20768
rect 30434 20712 30439 20768
rect 29913 20710 30439 20712
rect 29748 20708 29754 20710
rect 29637 20707 29703 20708
rect 29913 20707 29979 20710
rect 30373 20707 30439 20710
rect 31150 20708 31156 20772
rect 31220 20770 31226 20772
rect 31293 20770 31359 20773
rect 31220 20768 31359 20770
rect 31220 20712 31298 20768
rect 31354 20712 31359 20768
rect 31220 20710 31359 20712
rect 31220 20708 31226 20710
rect 31293 20707 31359 20710
rect 8628 20704 8944 20705
rect 8628 20640 8634 20704
rect 8698 20640 8714 20704
rect 8778 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8944 20704
rect 8628 20639 8944 20640
rect 16310 20704 16626 20705
rect 16310 20640 16316 20704
rect 16380 20640 16396 20704
rect 16460 20640 16476 20704
rect 16540 20640 16556 20704
rect 16620 20640 16626 20704
rect 16310 20639 16626 20640
rect 23992 20704 24308 20705
rect 23992 20640 23998 20704
rect 24062 20640 24078 20704
rect 24142 20640 24158 20704
rect 24222 20640 24238 20704
rect 24302 20640 24308 20704
rect 23992 20639 24308 20640
rect 31674 20704 31990 20705
rect 31674 20640 31680 20704
rect 31744 20640 31760 20704
rect 31824 20640 31840 20704
rect 31904 20640 31920 20704
rect 31984 20640 31990 20704
rect 31674 20639 31990 20640
rect 8342 20632 8451 20637
rect 8342 20576 8390 20632
rect 8446 20576 8451 20632
rect 8342 20574 8451 20576
rect 8385 20571 8451 20574
rect 9029 20634 9095 20637
rect 12341 20634 12407 20637
rect 9029 20632 12407 20634
rect 9029 20576 9034 20632
rect 9090 20576 12346 20632
rect 12402 20576 12407 20632
rect 9029 20574 12407 20576
rect 9029 20571 9095 20574
rect 12341 20571 12407 20574
rect 12893 20634 12959 20637
rect 13537 20634 13603 20637
rect 12893 20632 13603 20634
rect 12893 20576 12898 20632
rect 12954 20576 13542 20632
rect 13598 20576 13603 20632
rect 12893 20574 13603 20576
rect 12893 20571 12959 20574
rect 13537 20571 13603 20574
rect 14590 20572 14596 20636
rect 14660 20634 14666 20636
rect 16113 20634 16179 20637
rect 14660 20632 16179 20634
rect 14660 20576 16118 20632
rect 16174 20576 16179 20632
rect 14660 20574 16179 20576
rect 14660 20572 14666 20574
rect 16113 20571 16179 20574
rect 16757 20634 16823 20637
rect 18873 20634 18939 20637
rect 16757 20632 18939 20634
rect 16757 20576 16762 20632
rect 16818 20576 18878 20632
rect 18934 20576 18939 20632
rect 16757 20574 18939 20576
rect 16757 20571 16823 20574
rect 18873 20571 18939 20574
rect 19190 20572 19196 20636
rect 19260 20634 19266 20636
rect 21633 20634 21699 20637
rect 19260 20632 21699 20634
rect 19260 20576 21638 20632
rect 21694 20576 21699 20632
rect 19260 20574 21699 20576
rect 19260 20572 19266 20574
rect 21633 20571 21699 20574
rect 25497 20634 25563 20637
rect 26734 20634 26740 20636
rect 25497 20632 26740 20634
rect 25497 20576 25502 20632
rect 25558 20576 26740 20632
rect 25497 20574 26740 20576
rect 25497 20571 25563 20574
rect 26734 20572 26740 20574
rect 26804 20634 26810 20636
rect 27286 20634 27292 20636
rect 26804 20574 27292 20634
rect 26804 20572 26810 20574
rect 27286 20572 27292 20574
rect 27356 20572 27362 20636
rect 27521 20634 27587 20637
rect 30281 20634 30347 20637
rect 27521 20632 30347 20634
rect 27521 20576 27526 20632
rect 27582 20576 30286 20632
rect 30342 20576 30347 20632
rect 27521 20574 30347 20576
rect 27521 20571 27587 20574
rect 30281 20571 30347 20574
rect 10409 20498 10475 20501
rect 22277 20498 22343 20501
rect 10409 20496 22343 20498
rect 10409 20440 10414 20496
rect 10470 20440 22282 20496
rect 22338 20440 22343 20496
rect 10409 20438 22343 20440
rect 10409 20435 10475 20438
rect 22277 20435 22343 20438
rect 23054 20436 23060 20500
rect 23124 20498 23130 20500
rect 29729 20498 29795 20501
rect 23124 20496 29795 20498
rect 23124 20440 29734 20496
rect 29790 20440 29795 20496
rect 23124 20438 29795 20440
rect 23124 20436 23130 20438
rect 29729 20435 29795 20438
rect 29913 20498 29979 20501
rect 30230 20498 30236 20500
rect 29913 20496 30236 20498
rect 29913 20440 29918 20496
rect 29974 20440 30236 20496
rect 29913 20438 30236 20440
rect 29913 20435 29979 20438
rect 30230 20436 30236 20438
rect 30300 20436 30306 20500
rect 0 20362 800 20392
rect 1577 20362 1643 20365
rect 0 20360 1643 20362
rect 0 20304 1582 20360
rect 1638 20304 1643 20360
rect 0 20302 1643 20304
rect 0 20272 800 20302
rect 1577 20299 1643 20302
rect 3969 20362 4035 20365
rect 9673 20362 9739 20365
rect 22001 20362 22067 20365
rect 26417 20362 26483 20365
rect 26693 20362 26759 20365
rect 3969 20360 9506 20362
rect 3969 20304 3974 20360
rect 4030 20304 9506 20360
rect 3969 20302 9506 20304
rect 3969 20299 4035 20302
rect 9446 20226 9506 20302
rect 9673 20360 22067 20362
rect 9673 20304 9678 20360
rect 9734 20304 22006 20360
rect 22062 20304 22067 20360
rect 9673 20302 22067 20304
rect 9673 20299 9739 20302
rect 22001 20299 22067 20302
rect 22142 20360 26759 20362
rect 22142 20304 26422 20360
rect 26478 20304 26698 20360
rect 26754 20304 26759 20360
rect 22142 20302 26759 20304
rect 11237 20226 11303 20229
rect 9446 20224 11303 20226
rect 9446 20168 11242 20224
rect 11298 20168 11303 20224
rect 9446 20166 11303 20168
rect 11237 20163 11303 20166
rect 15193 20226 15259 20229
rect 18137 20226 18203 20229
rect 18413 20226 18479 20229
rect 19885 20226 19951 20229
rect 15193 20224 19951 20226
rect 15193 20168 15198 20224
rect 15254 20168 18142 20224
rect 18198 20168 18418 20224
rect 18474 20168 19890 20224
rect 19946 20168 19951 20224
rect 15193 20166 19951 20168
rect 15193 20163 15259 20166
rect 18137 20163 18203 20166
rect 18413 20163 18479 20166
rect 19885 20163 19951 20166
rect 20621 20226 20687 20229
rect 22142 20226 22202 20302
rect 26417 20299 26483 20302
rect 26693 20299 26759 20302
rect 26877 20362 26943 20365
rect 27102 20362 27108 20364
rect 26877 20360 27108 20362
rect 26877 20304 26882 20360
rect 26938 20304 27108 20360
rect 26877 20302 27108 20304
rect 26877 20299 26943 20302
rect 27102 20300 27108 20302
rect 27172 20300 27178 20364
rect 27286 20300 27292 20364
rect 27356 20362 27362 20364
rect 27797 20362 27863 20365
rect 27356 20360 27863 20362
rect 27356 20304 27802 20360
rect 27858 20304 27863 20360
rect 27356 20302 27863 20304
rect 27356 20300 27362 20302
rect 27797 20299 27863 20302
rect 28390 20300 28396 20364
rect 28460 20362 28466 20364
rect 28809 20362 28875 20365
rect 28460 20360 28875 20362
rect 28460 20304 28814 20360
rect 28870 20304 28875 20360
rect 28460 20302 28875 20304
rect 28460 20300 28466 20302
rect 28809 20299 28875 20302
rect 28993 20362 29059 20365
rect 30465 20362 30531 20365
rect 28993 20360 30531 20362
rect 28993 20304 28998 20360
rect 29054 20304 30470 20360
rect 30526 20304 30531 20360
rect 28993 20302 30531 20304
rect 28993 20299 29059 20302
rect 30465 20299 30531 20302
rect 20621 20224 22202 20226
rect 20621 20168 20626 20224
rect 20682 20168 22202 20224
rect 20621 20166 22202 20168
rect 22369 20226 22435 20229
rect 27654 20226 27660 20228
rect 22369 20224 27660 20226
rect 22369 20168 22374 20224
rect 22430 20168 27660 20224
rect 22369 20166 27660 20168
rect 20621 20163 20687 20166
rect 22369 20163 22435 20166
rect 27654 20164 27660 20166
rect 27724 20164 27730 20228
rect 28625 20226 28691 20229
rect 30046 20226 30052 20228
rect 28625 20224 30052 20226
rect 28625 20168 28630 20224
rect 28686 20168 30052 20224
rect 28625 20166 30052 20168
rect 28625 20163 28691 20166
rect 30046 20164 30052 20166
rect 30116 20164 30122 20228
rect 31477 20226 31543 20229
rect 32206 20226 33006 20256
rect 31477 20224 33006 20226
rect 31477 20168 31482 20224
rect 31538 20168 33006 20224
rect 31477 20166 33006 20168
rect 31477 20163 31543 20166
rect 4787 20160 5103 20161
rect 4787 20096 4793 20160
rect 4857 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5103 20160
rect 4787 20095 5103 20096
rect 12469 20160 12785 20161
rect 12469 20096 12475 20160
rect 12539 20096 12555 20160
rect 12619 20096 12635 20160
rect 12699 20096 12715 20160
rect 12779 20096 12785 20160
rect 12469 20095 12785 20096
rect 20151 20160 20467 20161
rect 20151 20096 20157 20160
rect 20221 20096 20237 20160
rect 20301 20096 20317 20160
rect 20381 20096 20397 20160
rect 20461 20096 20467 20160
rect 20151 20095 20467 20096
rect 27833 20160 28149 20161
rect 27833 20096 27839 20160
rect 27903 20096 27919 20160
rect 27983 20096 27999 20160
rect 28063 20096 28079 20160
rect 28143 20096 28149 20160
rect 32206 20136 33006 20166
rect 27833 20095 28149 20096
rect 10593 20090 10659 20093
rect 12249 20090 12315 20093
rect 10593 20088 12315 20090
rect 10593 20032 10598 20088
rect 10654 20032 12254 20088
rect 12310 20032 12315 20088
rect 10593 20030 12315 20032
rect 10593 20027 10659 20030
rect 12249 20027 12315 20030
rect 12934 20028 12940 20092
rect 13004 20090 13010 20092
rect 13813 20090 13879 20093
rect 13004 20088 13879 20090
rect 13004 20032 13818 20088
rect 13874 20032 13879 20088
rect 13004 20030 13879 20032
rect 13004 20028 13010 20030
rect 13813 20027 13879 20030
rect 14825 20090 14891 20093
rect 15377 20090 15443 20093
rect 18045 20090 18111 20093
rect 18229 20090 18295 20093
rect 14825 20088 18295 20090
rect 14825 20032 14830 20088
rect 14886 20032 15382 20088
rect 15438 20032 18050 20088
rect 18106 20032 18234 20088
rect 18290 20032 18295 20088
rect 14825 20030 18295 20032
rect 14825 20027 14891 20030
rect 15377 20027 15443 20030
rect 18045 20027 18111 20030
rect 18229 20027 18295 20030
rect 18413 20090 18479 20093
rect 19006 20090 19012 20092
rect 18413 20088 19012 20090
rect 18413 20032 18418 20088
rect 18474 20032 19012 20088
rect 18413 20030 19012 20032
rect 18413 20027 18479 20030
rect 19006 20028 19012 20030
rect 19076 20028 19082 20092
rect 19374 20028 19380 20092
rect 19444 20090 19450 20092
rect 19609 20090 19675 20093
rect 25998 20090 26004 20092
rect 19444 20088 19675 20090
rect 19444 20032 19614 20088
rect 19670 20032 19675 20088
rect 19444 20030 19675 20032
rect 19444 20028 19450 20030
rect 19609 20027 19675 20030
rect 22142 20030 26004 20090
rect 11053 19954 11119 19957
rect 17166 19954 17172 19956
rect 11053 19952 17172 19954
rect 11053 19896 11058 19952
rect 11114 19896 17172 19952
rect 11053 19894 17172 19896
rect 11053 19891 11119 19894
rect 17166 19892 17172 19894
rect 17236 19892 17242 19956
rect 17401 19954 17467 19957
rect 18229 19954 18295 19957
rect 17401 19952 18295 19954
rect 17401 19896 17406 19952
rect 17462 19896 18234 19952
rect 18290 19896 18295 19952
rect 17401 19894 18295 19896
rect 17401 19891 17467 19894
rect 18229 19891 18295 19894
rect 18454 19892 18460 19956
rect 18524 19954 18530 19956
rect 19241 19954 19307 19957
rect 22001 19954 22067 19957
rect 18524 19894 18890 19954
rect 18524 19892 18530 19894
rect 18830 19821 18890 19894
rect 19241 19952 22067 19954
rect 19241 19896 19246 19952
rect 19302 19896 22006 19952
rect 22062 19896 22067 19952
rect 19241 19894 22067 19896
rect 19241 19891 19307 19894
rect 22001 19891 22067 19894
rect 12801 19818 12867 19821
rect 18689 19818 18755 19821
rect 12801 19816 18755 19818
rect 12801 19760 12806 19816
rect 12862 19760 18694 19816
rect 18750 19760 18755 19816
rect 12801 19758 18755 19760
rect 18830 19816 18939 19821
rect 18830 19760 18878 19816
rect 18934 19760 18939 19816
rect 18830 19758 18939 19760
rect 12801 19755 12867 19758
rect 18689 19755 18755 19758
rect 18873 19755 18939 19758
rect 19149 19818 19215 19821
rect 22142 19818 22202 20030
rect 25998 20028 26004 20030
rect 26068 20028 26074 20092
rect 26141 20090 26207 20093
rect 26366 20090 26372 20092
rect 26141 20088 26372 20090
rect 26141 20032 26146 20088
rect 26202 20032 26372 20088
rect 26141 20030 26372 20032
rect 26141 20027 26207 20030
rect 26366 20028 26372 20030
rect 26436 20028 26442 20092
rect 27245 20090 27311 20093
rect 27429 20090 27495 20093
rect 27245 20088 27495 20090
rect 27245 20032 27250 20088
rect 27306 20032 27434 20088
rect 27490 20032 27495 20088
rect 27245 20030 27495 20032
rect 27245 20027 27311 20030
rect 27429 20027 27495 20030
rect 28257 20090 28323 20093
rect 28574 20090 28580 20092
rect 28257 20088 28580 20090
rect 28257 20032 28262 20088
rect 28318 20032 28580 20088
rect 28257 20030 28580 20032
rect 28257 20027 28323 20030
rect 28574 20028 28580 20030
rect 28644 20028 28650 20092
rect 28942 20028 28948 20092
rect 29012 20090 29018 20092
rect 30741 20090 30807 20093
rect 29012 20088 30807 20090
rect 29012 20032 30746 20088
rect 30802 20032 30807 20088
rect 29012 20030 30807 20032
rect 29012 20028 29018 20030
rect 30741 20027 30807 20030
rect 22737 19954 22803 19957
rect 23054 19954 23060 19956
rect 22737 19952 23060 19954
rect 22737 19896 22742 19952
rect 22798 19896 23060 19952
rect 22737 19894 23060 19896
rect 22737 19891 22803 19894
rect 23054 19892 23060 19894
rect 23124 19892 23130 19956
rect 23238 19892 23244 19956
rect 23308 19954 23314 19956
rect 30465 19954 30531 19957
rect 23308 19952 30531 19954
rect 23308 19896 30470 19952
rect 30526 19896 30531 19952
rect 23308 19894 30531 19896
rect 23308 19892 23314 19894
rect 30465 19891 30531 19894
rect 19149 19816 22202 19818
rect 19149 19760 19154 19816
rect 19210 19760 22202 19816
rect 19149 19758 22202 19760
rect 19149 19755 19215 19758
rect 24894 19756 24900 19820
rect 24964 19818 24970 19820
rect 25037 19818 25103 19821
rect 25681 19820 25747 19821
rect 25630 19818 25636 19820
rect 24964 19816 25103 19818
rect 24964 19760 25042 19816
rect 25098 19760 25103 19816
rect 24964 19758 25103 19760
rect 25590 19758 25636 19818
rect 25700 19816 25747 19820
rect 26877 19820 26943 19821
rect 26877 19818 26924 19820
rect 25742 19760 25747 19816
rect 24964 19756 24970 19758
rect 25037 19755 25103 19758
rect 25630 19756 25636 19758
rect 25700 19756 25747 19760
rect 26832 19816 26924 19818
rect 26832 19760 26882 19816
rect 26832 19758 26924 19760
rect 25681 19755 25747 19756
rect 26877 19756 26924 19758
rect 26988 19756 26994 19820
rect 27102 19756 27108 19820
rect 27172 19818 27178 19820
rect 30465 19818 30531 19821
rect 31385 19818 31451 19821
rect 27172 19816 31451 19818
rect 27172 19760 30470 19816
rect 30526 19760 31390 19816
rect 31446 19760 31451 19816
rect 27172 19758 31451 19760
rect 27172 19756 27178 19758
rect 26877 19755 26943 19756
rect 30465 19755 30531 19758
rect 31385 19755 31451 19758
rect 12065 19682 12131 19685
rect 13997 19682 14063 19685
rect 15837 19682 15903 19685
rect 12065 19680 13830 19682
rect 12065 19624 12070 19680
rect 12126 19624 13830 19680
rect 12065 19622 13830 19624
rect 12065 19619 12131 19622
rect 8628 19616 8944 19617
rect 0 19456 800 19576
rect 8628 19552 8634 19616
rect 8698 19552 8714 19616
rect 8778 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8944 19616
rect 8628 19551 8944 19552
rect 10777 19546 10843 19549
rect 11789 19546 11855 19549
rect 10777 19544 11855 19546
rect 10777 19488 10782 19544
rect 10838 19488 11794 19544
rect 11850 19488 11855 19544
rect 10777 19486 11855 19488
rect 10777 19483 10843 19486
rect 11789 19483 11855 19486
rect 12525 19546 12591 19549
rect 12985 19546 13051 19549
rect 12525 19544 13051 19546
rect 12525 19488 12530 19544
rect 12586 19488 12990 19544
rect 13046 19488 13051 19544
rect 12525 19486 13051 19488
rect 12525 19483 12591 19486
rect 12985 19483 13051 19486
rect 13445 19546 13511 19549
rect 13770 19546 13830 19622
rect 13997 19680 15903 19682
rect 13997 19624 14002 19680
rect 14058 19624 15842 19680
rect 15898 19624 15903 19680
rect 13997 19622 15903 19624
rect 13997 19619 14063 19622
rect 15837 19619 15903 19622
rect 16757 19682 16823 19685
rect 18781 19682 18847 19685
rect 16757 19680 18847 19682
rect 16757 19624 16762 19680
rect 16818 19624 18786 19680
rect 18842 19624 18847 19680
rect 16757 19622 18847 19624
rect 16757 19619 16823 19622
rect 18781 19619 18847 19622
rect 18965 19682 19031 19685
rect 20069 19682 20135 19685
rect 22093 19682 22159 19685
rect 18965 19680 19856 19682
rect 18965 19624 18970 19680
rect 19026 19624 19856 19680
rect 18965 19622 19856 19624
rect 18965 19619 19031 19622
rect 16310 19616 16626 19617
rect 16310 19552 16316 19616
rect 16380 19552 16396 19616
rect 16460 19552 16476 19616
rect 16540 19552 16556 19616
rect 16620 19552 16626 19616
rect 16310 19551 16626 19552
rect 19796 19549 19856 19622
rect 20069 19680 22159 19682
rect 20069 19624 20074 19680
rect 20130 19624 22098 19680
rect 22154 19624 22159 19680
rect 20069 19622 22159 19624
rect 20069 19619 20135 19622
rect 22093 19619 22159 19622
rect 27705 19682 27771 19685
rect 27705 19680 30114 19682
rect 27705 19624 27710 19680
rect 27766 19624 30114 19680
rect 27705 19622 30114 19624
rect 27705 19619 27771 19622
rect 23992 19616 24308 19617
rect 23992 19552 23998 19616
rect 24062 19552 24078 19616
rect 24142 19552 24158 19616
rect 24222 19552 24238 19616
rect 24302 19552 24308 19616
rect 23992 19551 24308 19552
rect 15510 19546 15516 19548
rect 13445 19544 13554 19546
rect 13445 19488 13450 19544
rect 13506 19488 13554 19544
rect 13445 19483 13554 19488
rect 13770 19486 15516 19546
rect 15510 19484 15516 19486
rect 15580 19484 15586 19548
rect 15878 19484 15884 19548
rect 15948 19546 15954 19548
rect 16113 19546 16179 19549
rect 15948 19544 16179 19546
rect 15948 19488 16118 19544
rect 16174 19488 16179 19544
rect 15948 19486 16179 19488
rect 15948 19484 15954 19486
rect 16113 19483 16179 19486
rect 16849 19546 16915 19549
rect 18638 19546 18644 19548
rect 16849 19544 18644 19546
rect 16849 19488 16854 19544
rect 16910 19488 18644 19544
rect 16849 19486 18644 19488
rect 16849 19483 16915 19486
rect 18638 19484 18644 19486
rect 18708 19484 18714 19548
rect 18781 19546 18847 19549
rect 19374 19546 19380 19548
rect 18781 19544 19380 19546
rect 18781 19488 18786 19544
rect 18842 19488 19380 19544
rect 18781 19486 19380 19488
rect 18781 19483 18847 19486
rect 19374 19484 19380 19486
rect 19444 19484 19450 19548
rect 19793 19544 19859 19549
rect 19793 19488 19798 19544
rect 19854 19488 19859 19544
rect 19793 19483 19859 19488
rect 19926 19484 19932 19548
rect 19996 19546 20002 19548
rect 23565 19546 23631 19549
rect 19996 19544 23631 19546
rect 19996 19488 23570 19544
rect 23626 19488 23631 19544
rect 19996 19486 23631 19488
rect 19996 19484 20002 19486
rect 23565 19483 23631 19486
rect 24577 19546 24643 19549
rect 25589 19546 25655 19549
rect 24577 19544 25655 19546
rect 24577 19488 24582 19544
rect 24638 19488 25594 19544
rect 25650 19488 25655 19544
rect 24577 19486 25655 19488
rect 24577 19483 24643 19486
rect 25589 19483 25655 19486
rect 25773 19546 25839 19549
rect 29494 19546 29500 19548
rect 25773 19544 29500 19546
rect 25773 19488 25778 19544
rect 25834 19488 29500 19544
rect 25773 19486 29500 19488
rect 25773 19483 25839 19486
rect 29494 19484 29500 19486
rect 29564 19546 29570 19548
rect 29913 19546 29979 19549
rect 29564 19544 29979 19546
rect 29564 19488 29918 19544
rect 29974 19488 29979 19544
rect 29564 19486 29979 19488
rect 30054 19546 30114 19622
rect 30414 19620 30420 19684
rect 30484 19682 30490 19684
rect 31109 19682 31175 19685
rect 30484 19680 31175 19682
rect 30484 19624 31114 19680
rect 31170 19624 31175 19680
rect 30484 19622 31175 19624
rect 30484 19620 30490 19622
rect 31109 19619 31175 19622
rect 31674 19616 31990 19617
rect 31674 19552 31680 19616
rect 31744 19552 31760 19616
rect 31824 19552 31840 19616
rect 31904 19552 31920 19616
rect 31984 19552 31990 19616
rect 31674 19551 31990 19552
rect 30782 19546 30788 19548
rect 30054 19486 30788 19546
rect 29564 19484 29570 19486
rect 29913 19483 29979 19486
rect 30782 19484 30788 19486
rect 30852 19484 30858 19548
rect 32206 19546 33006 19576
rect 32078 19486 33006 19546
rect 7649 19410 7715 19413
rect 12801 19410 12867 19413
rect 7649 19408 12867 19410
rect 7649 19352 7654 19408
rect 7710 19352 12806 19408
rect 12862 19352 12867 19408
rect 7649 19350 12867 19352
rect 7649 19347 7715 19350
rect 12801 19347 12867 19350
rect 13261 19412 13327 19413
rect 13261 19408 13308 19412
rect 13372 19410 13378 19412
rect 13494 19410 13554 19483
rect 16297 19410 16363 19413
rect 18689 19410 18755 19413
rect 19149 19410 19215 19413
rect 13261 19352 13266 19408
rect 13261 19348 13308 19352
rect 13372 19350 13418 19410
rect 13494 19408 19215 19410
rect 13494 19352 16302 19408
rect 16358 19352 18694 19408
rect 18750 19352 19154 19408
rect 19210 19352 19215 19408
rect 13494 19350 19215 19352
rect 13372 19348 13378 19350
rect 13261 19347 13327 19348
rect 16297 19347 16363 19350
rect 18689 19347 18755 19350
rect 19149 19347 19215 19350
rect 19374 19348 19380 19412
rect 19444 19410 19450 19412
rect 20524 19410 20530 19412
rect 19444 19350 20530 19410
rect 19444 19348 19450 19350
rect 20524 19348 20530 19350
rect 20594 19348 20600 19412
rect 24853 19410 24919 19413
rect 20670 19408 24919 19410
rect 20670 19352 24858 19408
rect 24914 19352 24919 19408
rect 20670 19350 24919 19352
rect 10961 19274 11027 19277
rect 13445 19274 13511 19277
rect 20670 19274 20730 19350
rect 24853 19347 24919 19350
rect 25037 19410 25103 19413
rect 27245 19410 27311 19413
rect 27705 19410 27771 19413
rect 25037 19408 27771 19410
rect 25037 19352 25042 19408
rect 25098 19352 27250 19408
rect 27306 19352 27710 19408
rect 27766 19352 27771 19408
rect 25037 19350 27771 19352
rect 25037 19347 25103 19350
rect 27245 19347 27311 19350
rect 27705 19347 27771 19350
rect 28206 19348 28212 19412
rect 28276 19410 28282 19412
rect 28625 19410 28691 19413
rect 28276 19408 28691 19410
rect 28276 19352 28630 19408
rect 28686 19352 28691 19408
rect 28276 19350 28691 19352
rect 28276 19348 28282 19350
rect 28625 19347 28691 19350
rect 28993 19410 29059 19413
rect 29310 19410 29316 19412
rect 28993 19408 29316 19410
rect 28993 19352 28998 19408
rect 29054 19352 29316 19408
rect 28993 19350 29316 19352
rect 28993 19347 29059 19350
rect 29310 19348 29316 19350
rect 29380 19348 29386 19412
rect 29862 19348 29868 19412
rect 29932 19410 29938 19412
rect 30005 19410 30071 19413
rect 30281 19412 30347 19413
rect 29932 19408 30071 19410
rect 29932 19352 30010 19408
rect 30066 19352 30071 19408
rect 29932 19350 30071 19352
rect 29932 19348 29938 19350
rect 30005 19347 30071 19350
rect 30230 19348 30236 19412
rect 30300 19410 30347 19412
rect 31385 19410 31451 19413
rect 32078 19410 32138 19486
rect 32206 19456 33006 19486
rect 30300 19408 30392 19410
rect 30342 19352 30392 19408
rect 30300 19350 30392 19352
rect 31385 19408 32138 19410
rect 31385 19352 31390 19408
rect 31446 19352 32138 19408
rect 31385 19350 32138 19352
rect 30300 19348 30347 19350
rect 30281 19347 30347 19348
rect 31385 19347 31451 19350
rect 31017 19274 31083 19277
rect 10961 19272 13370 19274
rect 10961 19216 10966 19272
rect 11022 19216 13370 19272
rect 10961 19214 13370 19216
rect 10961 19211 11027 19214
rect 9673 19138 9739 19141
rect 12341 19138 12407 19141
rect 9673 19136 12407 19138
rect 9673 19080 9678 19136
rect 9734 19080 12346 19136
rect 12402 19080 12407 19136
rect 9673 19078 12407 19080
rect 9673 19075 9739 19078
rect 12341 19075 12407 19078
rect 4787 19072 5103 19073
rect 4787 19008 4793 19072
rect 4857 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5103 19072
rect 4787 19007 5103 19008
rect 12469 19072 12785 19073
rect 12469 19008 12475 19072
rect 12539 19008 12555 19072
rect 12619 19008 12635 19072
rect 12699 19008 12715 19072
rect 12779 19008 12785 19072
rect 12469 19007 12785 19008
rect 11789 18866 11855 18869
rect 12934 18866 12940 18868
rect 11789 18864 12940 18866
rect 11789 18808 11794 18864
rect 11850 18808 12940 18864
rect 11789 18806 12940 18808
rect 11789 18803 11855 18806
rect 12934 18804 12940 18806
rect 13004 18804 13010 18868
rect 0 18730 800 18760
rect 1577 18730 1643 18733
rect 0 18728 1643 18730
rect 0 18672 1582 18728
rect 1638 18672 1643 18728
rect 0 18670 1643 18672
rect 0 18640 800 18670
rect 1577 18667 1643 18670
rect 13310 18594 13370 19214
rect 13445 19272 20730 19274
rect 13445 19216 13450 19272
rect 13506 19216 20730 19272
rect 13445 19214 20730 19216
rect 21728 19272 31083 19274
rect 21728 19216 31022 19272
rect 31078 19216 31083 19272
rect 21728 19214 31083 19216
rect 13445 19211 13511 19214
rect 13721 19138 13787 19141
rect 14917 19138 14983 19141
rect 16941 19138 17007 19141
rect 13721 19136 17007 19138
rect 13721 19080 13726 19136
rect 13782 19080 14922 19136
rect 14978 19080 16946 19136
rect 17002 19080 17007 19136
rect 13721 19078 17007 19080
rect 13721 19075 13787 19078
rect 14917 19075 14983 19078
rect 16941 19075 17007 19078
rect 17585 19138 17651 19141
rect 18045 19138 18111 19141
rect 17585 19136 18111 19138
rect 17585 19080 17590 19136
rect 17646 19080 18050 19136
rect 18106 19080 18111 19136
rect 17585 19078 18111 19080
rect 17585 19075 17651 19078
rect 18045 19075 18111 19078
rect 18229 19138 18295 19141
rect 18822 19138 18828 19140
rect 18229 19136 18828 19138
rect 18229 19080 18234 19136
rect 18290 19080 18828 19136
rect 18229 19078 18828 19080
rect 18229 19075 18295 19078
rect 18822 19076 18828 19078
rect 18892 19138 18898 19140
rect 19149 19138 19215 19141
rect 18892 19136 19215 19138
rect 18892 19080 19154 19136
rect 19210 19080 19215 19136
rect 18892 19078 19215 19080
rect 18892 19076 18898 19078
rect 19149 19075 19215 19078
rect 19333 19138 19399 19141
rect 19885 19138 19951 19141
rect 19333 19136 19951 19138
rect 19333 19080 19338 19136
rect 19394 19080 19890 19136
rect 19946 19080 19951 19136
rect 19333 19078 19951 19080
rect 19333 19075 19399 19078
rect 19885 19075 19951 19078
rect 20529 19138 20595 19141
rect 21582 19138 21588 19140
rect 20529 19136 21588 19138
rect 20529 19080 20534 19136
rect 20590 19080 21588 19136
rect 20529 19078 21588 19080
rect 20529 19075 20595 19078
rect 21582 19076 21588 19078
rect 21652 19076 21658 19140
rect 20151 19072 20467 19073
rect 20151 19008 20157 19072
rect 20221 19008 20237 19072
rect 20301 19008 20317 19072
rect 20381 19008 20397 19072
rect 20461 19008 20467 19072
rect 20151 19007 20467 19008
rect 14457 19002 14523 19005
rect 16573 19002 16639 19005
rect 14457 19000 16639 19002
rect 14457 18944 14462 19000
rect 14518 18944 16578 19000
rect 16634 18944 16639 19000
rect 14457 18942 16639 18944
rect 14457 18939 14523 18942
rect 16573 18939 16639 18942
rect 16757 19002 16823 19005
rect 17677 19002 17743 19005
rect 16757 19000 17743 19002
rect 16757 18944 16762 19000
rect 16818 18944 17682 19000
rect 17738 18944 17743 19000
rect 16757 18942 17743 18944
rect 16757 18939 16823 18942
rect 17677 18939 17743 18942
rect 18137 19002 18203 19005
rect 19517 19002 19583 19005
rect 21728 19002 21788 19214
rect 31017 19211 31083 19214
rect 24025 19138 24091 19141
rect 26969 19140 27035 19141
rect 26182 19138 26188 19140
rect 24025 19136 26188 19138
rect 24025 19080 24030 19136
rect 24086 19080 26188 19136
rect 24025 19078 26188 19080
rect 24025 19075 24091 19078
rect 26182 19076 26188 19078
rect 26252 19076 26258 19140
rect 26550 19076 26556 19140
rect 26620 19138 26626 19140
rect 26620 19078 26848 19138
rect 26620 19076 26626 19078
rect 18137 19000 19583 19002
rect 18137 18944 18142 19000
rect 18198 18944 19522 19000
rect 19578 18944 19583 19000
rect 18137 18942 19583 18944
rect 18137 18939 18203 18942
rect 19517 18939 19583 18942
rect 20532 18942 21788 19002
rect 23105 19002 23171 19005
rect 24485 19002 24551 19005
rect 23105 19000 24551 19002
rect 23105 18944 23110 19000
rect 23166 18944 24490 19000
rect 24546 18944 24551 19000
rect 23105 18942 24551 18944
rect 13905 18866 13971 18869
rect 15377 18866 15443 18869
rect 15745 18868 15811 18869
rect 13905 18864 15443 18866
rect 13905 18808 13910 18864
rect 13966 18808 15382 18864
rect 15438 18808 15443 18864
rect 13905 18806 15443 18808
rect 13905 18803 13971 18806
rect 15377 18803 15443 18806
rect 15694 18804 15700 18868
rect 15764 18866 15811 18868
rect 15764 18864 15856 18866
rect 15806 18808 15856 18864
rect 15764 18806 15856 18808
rect 15764 18804 15811 18806
rect 16062 18804 16068 18868
rect 16132 18866 16138 18868
rect 17217 18866 17283 18869
rect 16132 18864 17283 18866
rect 16132 18808 17222 18864
rect 17278 18808 17283 18864
rect 16132 18806 17283 18808
rect 16132 18804 16138 18806
rect 15745 18803 15811 18804
rect 17217 18803 17283 18806
rect 17350 18804 17356 18868
rect 17420 18866 17426 18868
rect 20532 18866 20592 18942
rect 23105 18939 23171 18942
rect 24485 18939 24551 18942
rect 24894 18940 24900 19004
rect 24964 19002 24970 19004
rect 26509 19002 26575 19005
rect 24964 19000 26575 19002
rect 24964 18944 26514 19000
rect 26570 18944 26575 19000
rect 24964 18942 26575 18944
rect 26788 19002 26848 19078
rect 26918 19076 26924 19140
rect 26988 19138 27035 19140
rect 26988 19136 27080 19138
rect 27030 19080 27080 19136
rect 26988 19078 27080 19080
rect 28257 19136 28323 19141
rect 28257 19080 28262 19136
rect 28318 19080 28323 19136
rect 26988 19076 27035 19078
rect 26969 19075 27035 19076
rect 28257 19075 28323 19080
rect 28390 19076 28396 19140
rect 28460 19138 28466 19140
rect 28809 19138 28875 19141
rect 28460 19136 28875 19138
rect 28460 19080 28814 19136
rect 28870 19080 28875 19136
rect 28460 19078 28875 19080
rect 28460 19076 28466 19078
rect 28809 19075 28875 19078
rect 29177 19138 29243 19141
rect 29310 19138 29316 19140
rect 29177 19136 29316 19138
rect 29177 19080 29182 19136
rect 29238 19080 29316 19136
rect 29177 19078 29316 19080
rect 29177 19075 29243 19078
rect 29310 19076 29316 19078
rect 29380 19076 29386 19140
rect 27833 19072 28149 19073
rect 27833 19008 27839 19072
rect 27903 19008 27919 19072
rect 27983 19008 27999 19072
rect 28063 19008 28079 19072
rect 28143 19008 28149 19072
rect 27833 19007 28149 19008
rect 27429 19002 27495 19005
rect 26788 19000 27495 19002
rect 26788 18944 27434 19000
rect 27490 18944 27495 19000
rect 26788 18942 27495 18944
rect 28260 19002 28320 19075
rect 28441 19002 28507 19005
rect 28260 19000 28507 19002
rect 28260 18944 28446 19000
rect 28502 18944 28507 19000
rect 28260 18942 28507 18944
rect 24964 18940 24970 18942
rect 26509 18939 26575 18942
rect 27429 18939 27495 18942
rect 28441 18939 28507 18942
rect 29177 19002 29243 19005
rect 30465 19002 30531 19005
rect 29177 19000 30531 19002
rect 29177 18944 29182 19000
rect 29238 18944 30470 19000
rect 30526 18944 30531 19000
rect 29177 18942 30531 18944
rect 29177 18939 29243 18942
rect 30465 18939 30531 18942
rect 21950 18866 21956 18868
rect 17420 18806 20592 18866
rect 20670 18806 21956 18866
rect 17420 18804 17426 18806
rect 13445 18730 13511 18733
rect 14457 18730 14523 18733
rect 19517 18730 19583 18733
rect 13445 18728 19583 18730
rect 13445 18672 13450 18728
rect 13506 18672 14462 18728
rect 14518 18672 19522 18728
rect 19578 18672 19583 18728
rect 13445 18670 19583 18672
rect 13445 18667 13511 18670
rect 14457 18667 14523 18670
rect 19517 18667 19583 18670
rect 19742 18668 19748 18732
rect 19812 18730 19818 18732
rect 20670 18730 20730 18806
rect 21950 18804 21956 18806
rect 22020 18866 22026 18868
rect 30465 18866 30531 18869
rect 22020 18864 30531 18866
rect 22020 18808 30470 18864
rect 30526 18808 30531 18864
rect 22020 18806 30531 18808
rect 22020 18804 22026 18806
rect 30465 18803 30531 18806
rect 31017 18866 31083 18869
rect 32206 18866 33006 18896
rect 31017 18864 33006 18866
rect 31017 18808 31022 18864
rect 31078 18808 33006 18864
rect 31017 18806 33006 18808
rect 31017 18803 31083 18806
rect 32206 18776 33006 18806
rect 19812 18670 20730 18730
rect 19812 18668 19818 18670
rect 21398 18668 21404 18732
rect 21468 18730 21474 18732
rect 23105 18730 23171 18733
rect 21468 18728 23171 18730
rect 21468 18672 23110 18728
rect 23166 18672 23171 18728
rect 21468 18670 23171 18672
rect 21468 18668 21474 18670
rect 23105 18667 23171 18670
rect 23381 18730 23447 18733
rect 26693 18730 26759 18733
rect 23381 18728 26759 18730
rect 23381 18672 23386 18728
rect 23442 18672 26698 18728
rect 26754 18672 26759 18728
rect 23381 18670 26759 18672
rect 23381 18667 23447 18670
rect 26693 18667 26759 18670
rect 27245 18730 27311 18733
rect 27429 18730 27495 18733
rect 27245 18728 27495 18730
rect 27245 18672 27250 18728
rect 27306 18672 27434 18728
rect 27490 18672 27495 18728
rect 27245 18670 27495 18672
rect 27245 18667 27311 18670
rect 27429 18667 27495 18670
rect 27797 18730 27863 18733
rect 31334 18730 31340 18732
rect 27797 18728 31340 18730
rect 27797 18672 27802 18728
rect 27858 18672 31340 18728
rect 27797 18670 31340 18672
rect 27797 18667 27863 18670
rect 31334 18668 31340 18670
rect 31404 18730 31410 18732
rect 31661 18730 31727 18733
rect 31404 18728 31727 18730
rect 31404 18672 31666 18728
rect 31722 18672 31727 18728
rect 31404 18670 31727 18672
rect 31404 18668 31410 18670
rect 31661 18667 31727 18670
rect 16062 18594 16068 18596
rect 13310 18534 16068 18594
rect 16062 18532 16068 18534
rect 16132 18532 16138 18596
rect 17217 18594 17283 18597
rect 21081 18594 21147 18597
rect 17217 18592 21147 18594
rect 17217 18536 17222 18592
rect 17278 18536 21086 18592
rect 21142 18536 21147 18592
rect 17217 18534 21147 18536
rect 17217 18531 17283 18534
rect 21081 18531 21147 18534
rect 21582 18532 21588 18596
rect 21652 18594 21658 18596
rect 23013 18594 23079 18597
rect 21652 18592 23079 18594
rect 21652 18536 23018 18592
rect 23074 18536 23079 18592
rect 21652 18534 23079 18536
rect 21652 18532 21658 18534
rect 23013 18531 23079 18534
rect 24485 18594 24551 18597
rect 29085 18594 29151 18597
rect 24485 18592 29151 18594
rect 24485 18536 24490 18592
rect 24546 18536 29090 18592
rect 29146 18536 29151 18592
rect 24485 18534 29151 18536
rect 24485 18531 24551 18534
rect 29085 18531 29151 18534
rect 30097 18594 30163 18597
rect 30414 18594 30420 18596
rect 30097 18592 30420 18594
rect 30097 18536 30102 18592
rect 30158 18536 30420 18592
rect 30097 18534 30420 18536
rect 30097 18531 30163 18534
rect 30414 18532 30420 18534
rect 30484 18532 30490 18596
rect 30833 18594 30899 18597
rect 30833 18592 31034 18594
rect 30833 18536 30838 18592
rect 30894 18536 31034 18592
rect 30833 18534 31034 18536
rect 30833 18531 30899 18534
rect 8628 18528 8944 18529
rect 8628 18464 8634 18528
rect 8698 18464 8714 18528
rect 8778 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8944 18528
rect 8628 18463 8944 18464
rect 16310 18528 16626 18529
rect 16310 18464 16316 18528
rect 16380 18464 16396 18528
rect 16460 18464 16476 18528
rect 16540 18464 16556 18528
rect 16620 18464 16626 18528
rect 16310 18463 16626 18464
rect 23992 18528 24308 18529
rect 23992 18464 23998 18528
rect 24062 18464 24078 18528
rect 24142 18464 24158 18528
rect 24222 18464 24238 18528
rect 24302 18464 24308 18528
rect 23992 18463 24308 18464
rect 10041 18458 10107 18461
rect 10593 18458 10659 18461
rect 14917 18458 14983 18461
rect 16021 18458 16087 18461
rect 10041 18456 16087 18458
rect 10041 18400 10046 18456
rect 10102 18400 10598 18456
rect 10654 18400 14922 18456
rect 14978 18400 16026 18456
rect 16082 18400 16087 18456
rect 10041 18398 16087 18400
rect 10041 18395 10107 18398
rect 10593 18395 10659 18398
rect 14917 18395 14983 18398
rect 16021 18395 16087 18398
rect 16757 18460 16823 18461
rect 16757 18456 16804 18460
rect 16868 18458 16874 18460
rect 17033 18458 17099 18461
rect 24393 18458 24459 18461
rect 25773 18458 25839 18461
rect 16757 18400 16762 18456
rect 16757 18396 16804 18400
rect 16868 18398 16914 18458
rect 17033 18456 23352 18458
rect 17033 18400 17038 18456
rect 17094 18400 23352 18456
rect 17033 18398 23352 18400
rect 16868 18396 16874 18398
rect 16757 18395 16823 18396
rect 17033 18395 17099 18398
rect 13169 18322 13235 18325
rect 13813 18322 13879 18325
rect 13169 18320 13879 18322
rect 13169 18264 13174 18320
rect 13230 18264 13818 18320
rect 13874 18264 13879 18320
rect 13169 18262 13879 18264
rect 13169 18259 13235 18262
rect 13813 18259 13879 18262
rect 14089 18322 14155 18325
rect 22737 18322 22803 18325
rect 14089 18320 22803 18322
rect 14089 18264 14094 18320
rect 14150 18264 22742 18320
rect 22798 18264 22803 18320
rect 14089 18262 22803 18264
rect 23292 18322 23352 18398
rect 24393 18456 25839 18458
rect 24393 18400 24398 18456
rect 24454 18400 25778 18456
rect 25834 18400 25839 18456
rect 24393 18398 25839 18400
rect 24393 18395 24459 18398
rect 25773 18395 25839 18398
rect 25998 18396 26004 18460
rect 26068 18458 26074 18460
rect 30833 18458 30899 18461
rect 26068 18456 30899 18458
rect 26068 18400 30838 18456
rect 30894 18400 30899 18456
rect 26068 18398 30899 18400
rect 26068 18396 26074 18398
rect 30833 18395 30899 18398
rect 26509 18322 26575 18325
rect 23292 18320 26575 18322
rect 23292 18264 26514 18320
rect 26570 18264 26575 18320
rect 23292 18262 26575 18264
rect 14089 18259 14155 18262
rect 22737 18259 22803 18262
rect 26509 18259 26575 18262
rect 26877 18322 26943 18325
rect 28533 18322 28599 18325
rect 26877 18320 28599 18322
rect 26877 18264 26882 18320
rect 26938 18264 28538 18320
rect 28594 18264 28599 18320
rect 26877 18262 28599 18264
rect 26877 18259 26943 18262
rect 28533 18259 28599 18262
rect 29126 18260 29132 18324
rect 29196 18322 29202 18324
rect 29361 18322 29427 18325
rect 30974 18322 31034 18534
rect 31674 18528 31990 18529
rect 31674 18464 31680 18528
rect 31744 18464 31760 18528
rect 31824 18464 31840 18528
rect 31904 18464 31920 18528
rect 31984 18464 31990 18528
rect 31674 18463 31990 18464
rect 29196 18320 29427 18322
rect 29196 18264 29366 18320
rect 29422 18264 29427 18320
rect 29196 18262 29427 18264
rect 29196 18260 29202 18262
rect 29361 18259 29427 18262
rect 29502 18262 31034 18322
rect 11605 18186 11671 18189
rect 24485 18186 24551 18189
rect 11605 18184 24551 18186
rect 11605 18128 11610 18184
rect 11666 18128 24490 18184
rect 24546 18128 24551 18184
rect 11605 18126 24551 18128
rect 11605 18123 11671 18126
rect 24485 18123 24551 18126
rect 25446 18124 25452 18188
rect 25516 18186 25522 18188
rect 25957 18186 26023 18189
rect 25516 18184 26023 18186
rect 25516 18128 25962 18184
rect 26018 18128 26023 18184
rect 25516 18126 26023 18128
rect 25516 18124 25522 18126
rect 25957 18123 26023 18126
rect 26325 18188 26391 18189
rect 26325 18184 26372 18188
rect 26436 18186 26442 18188
rect 26969 18186 27035 18189
rect 27521 18186 27587 18189
rect 26325 18128 26330 18184
rect 26325 18124 26372 18128
rect 26436 18126 26482 18186
rect 26969 18184 27587 18186
rect 26969 18128 26974 18184
rect 27030 18128 27526 18184
rect 27582 18128 27587 18184
rect 26969 18126 27587 18128
rect 26436 18124 26442 18126
rect 26325 18123 26391 18124
rect 26969 18123 27035 18126
rect 27521 18123 27587 18126
rect 28073 18186 28139 18189
rect 28073 18184 28274 18186
rect 28073 18128 28078 18184
rect 28134 18128 28274 18184
rect 28073 18126 28274 18128
rect 28073 18123 28139 18126
rect 14825 18050 14891 18053
rect 19793 18050 19859 18053
rect 14825 18048 19859 18050
rect 14825 17992 14830 18048
rect 14886 17992 19798 18048
rect 19854 17992 19859 18048
rect 14825 17990 19859 17992
rect 14825 17987 14891 17990
rect 19793 17987 19859 17990
rect 21725 18050 21791 18053
rect 23657 18050 23723 18053
rect 24761 18052 24827 18053
rect 24710 18050 24716 18052
rect 21725 18048 23723 18050
rect 21725 17992 21730 18048
rect 21786 17992 23662 18048
rect 23718 17992 23723 18048
rect 21725 17990 23723 17992
rect 24670 17990 24716 18050
rect 24780 18048 24827 18052
rect 24822 17992 24827 18048
rect 21725 17987 21791 17990
rect 23657 17987 23723 17990
rect 24710 17988 24716 17990
rect 24780 17988 24827 17992
rect 24761 17987 24827 17988
rect 25221 18050 25287 18053
rect 27286 18050 27292 18052
rect 25221 18048 27292 18050
rect 25221 17992 25226 18048
rect 25282 17992 27292 18048
rect 25221 17990 27292 17992
rect 25221 17987 25287 17990
rect 27286 17988 27292 17990
rect 27356 18050 27362 18052
rect 27429 18050 27495 18053
rect 27356 18048 27495 18050
rect 27356 17992 27434 18048
rect 27490 17992 27495 18048
rect 27356 17990 27495 17992
rect 28214 18050 28274 18126
rect 28390 18124 28396 18188
rect 28460 18186 28466 18188
rect 28625 18186 28691 18189
rect 28460 18184 28691 18186
rect 28460 18128 28630 18184
rect 28686 18128 28691 18184
rect 28460 18126 28691 18128
rect 28460 18124 28466 18126
rect 28625 18123 28691 18126
rect 29126 18124 29132 18188
rect 29196 18186 29202 18188
rect 29502 18186 29562 18262
rect 29196 18126 29562 18186
rect 29729 18186 29795 18189
rect 30189 18186 30255 18189
rect 29729 18184 30255 18186
rect 29729 18128 29734 18184
rect 29790 18128 30194 18184
rect 30250 18128 30255 18184
rect 29729 18126 30255 18128
rect 29196 18124 29202 18126
rect 29729 18123 29795 18126
rect 30189 18123 30255 18126
rect 30833 18186 30899 18189
rect 32206 18186 33006 18216
rect 30833 18184 33006 18186
rect 30833 18128 30838 18184
rect 30894 18128 33006 18184
rect 30833 18126 33006 18128
rect 30833 18123 30899 18126
rect 32206 18096 33006 18126
rect 30741 18050 30807 18053
rect 28214 18048 30807 18050
rect 28214 17992 30746 18048
rect 30802 17992 30807 18048
rect 28214 17990 30807 17992
rect 27356 17988 27362 17990
rect 27429 17987 27495 17990
rect 30741 17987 30807 17990
rect 4787 17984 5103 17985
rect 0 17914 800 17944
rect 4787 17920 4793 17984
rect 4857 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5103 17984
rect 4787 17919 5103 17920
rect 12469 17984 12785 17985
rect 12469 17920 12475 17984
rect 12539 17920 12555 17984
rect 12619 17920 12635 17984
rect 12699 17920 12715 17984
rect 12779 17920 12785 17984
rect 12469 17919 12785 17920
rect 20151 17984 20467 17985
rect 20151 17920 20157 17984
rect 20221 17920 20237 17984
rect 20301 17920 20317 17984
rect 20381 17920 20397 17984
rect 20461 17920 20467 17984
rect 20151 17919 20467 17920
rect 27833 17984 28149 17985
rect 27833 17920 27839 17984
rect 27903 17920 27919 17984
rect 27983 17920 27999 17984
rect 28063 17920 28079 17984
rect 28143 17920 28149 17984
rect 27833 17919 28149 17920
rect 1577 17914 1643 17917
rect 0 17912 1643 17914
rect 0 17856 1582 17912
rect 1638 17856 1643 17912
rect 0 17854 1643 17856
rect 0 17824 800 17854
rect 1577 17851 1643 17854
rect 13261 17914 13327 17917
rect 14549 17914 14615 17917
rect 15745 17914 15811 17917
rect 13261 17912 14244 17914
rect 13261 17856 13266 17912
rect 13322 17856 14244 17912
rect 13261 17854 14244 17856
rect 13261 17851 13327 17854
rect 3877 17778 3943 17781
rect 14038 17778 14044 17780
rect 3877 17776 14044 17778
rect 3877 17720 3882 17776
rect 3938 17720 14044 17776
rect 3877 17718 14044 17720
rect 3877 17715 3943 17718
rect 14038 17716 14044 17718
rect 14108 17716 14114 17780
rect 14184 17778 14244 17854
rect 14549 17912 15811 17914
rect 14549 17856 14554 17912
rect 14610 17856 15750 17912
rect 15806 17856 15811 17912
rect 14549 17854 15811 17856
rect 14549 17851 14615 17854
rect 15745 17851 15811 17854
rect 16389 17914 16455 17917
rect 16798 17914 16804 17916
rect 16389 17912 16804 17914
rect 16389 17856 16394 17912
rect 16450 17856 16804 17912
rect 16389 17854 16804 17856
rect 16389 17851 16455 17854
rect 16798 17852 16804 17854
rect 16868 17852 16874 17916
rect 16982 17852 16988 17916
rect 17052 17914 17058 17916
rect 17401 17914 17467 17917
rect 17052 17912 17467 17914
rect 17052 17856 17406 17912
rect 17462 17856 17467 17912
rect 17052 17854 17467 17856
rect 17052 17852 17058 17854
rect 17401 17851 17467 17854
rect 17585 17914 17651 17917
rect 19885 17914 19951 17917
rect 17585 17912 19951 17914
rect 17585 17856 17590 17912
rect 17646 17856 19890 17912
rect 19946 17856 19951 17912
rect 17585 17854 19951 17856
rect 17585 17851 17651 17854
rect 19885 17851 19951 17854
rect 21214 17852 21220 17916
rect 21284 17914 21290 17916
rect 26693 17914 26759 17917
rect 21284 17912 26759 17914
rect 21284 17856 26698 17912
rect 26754 17856 26759 17912
rect 21284 17854 26759 17856
rect 21284 17852 21290 17854
rect 26693 17851 26759 17854
rect 26969 17914 27035 17917
rect 27705 17914 27771 17917
rect 26969 17912 27771 17914
rect 26969 17856 26974 17912
rect 27030 17856 27710 17912
rect 27766 17856 27771 17912
rect 26969 17854 27771 17856
rect 26969 17851 27035 17854
rect 27705 17851 27771 17854
rect 28257 17914 28323 17917
rect 29821 17914 29887 17917
rect 30281 17916 30347 17917
rect 30230 17914 30236 17916
rect 28257 17912 29887 17914
rect 28257 17856 28262 17912
rect 28318 17856 29826 17912
rect 29882 17856 29887 17912
rect 28257 17854 29887 17856
rect 30190 17854 30236 17914
rect 30300 17912 30347 17916
rect 30342 17856 30347 17912
rect 28257 17851 28323 17854
rect 29821 17851 29887 17854
rect 30230 17852 30236 17854
rect 30300 17852 30347 17856
rect 30281 17851 30347 17852
rect 14917 17778 14983 17781
rect 14184 17776 14983 17778
rect 14184 17720 14922 17776
rect 14978 17720 14983 17776
rect 14184 17718 14983 17720
rect 14917 17715 14983 17718
rect 15101 17778 15167 17781
rect 16481 17778 16547 17781
rect 15101 17776 17096 17778
rect 15101 17720 15106 17776
rect 15162 17720 16486 17776
rect 16542 17720 17096 17776
rect 15101 17718 17096 17720
rect 15101 17715 15167 17718
rect 16481 17715 16547 17718
rect 13445 17642 13511 17645
rect 17036 17642 17096 17718
rect 17166 17716 17172 17780
rect 17236 17778 17242 17780
rect 21449 17778 21515 17781
rect 17236 17776 21515 17778
rect 17236 17720 21454 17776
rect 21510 17720 21515 17776
rect 17236 17718 21515 17720
rect 17236 17716 17242 17718
rect 21449 17715 21515 17718
rect 23197 17778 23263 17781
rect 26233 17780 26299 17781
rect 24894 17778 24900 17780
rect 23197 17776 24900 17778
rect 23197 17720 23202 17776
rect 23258 17720 24900 17776
rect 23197 17718 24900 17720
rect 23197 17715 23263 17718
rect 24894 17716 24900 17718
rect 24964 17716 24970 17780
rect 26182 17778 26188 17780
rect 26142 17718 26188 17778
rect 26252 17776 26299 17780
rect 27470 17778 27476 17780
rect 26294 17720 26299 17776
rect 26182 17716 26188 17718
rect 26252 17716 26299 17720
rect 26233 17715 26299 17716
rect 26374 17718 27476 17778
rect 18321 17642 18387 17645
rect 13445 17640 16820 17642
rect 13445 17584 13450 17640
rect 13506 17584 16820 17640
rect 13445 17582 16820 17584
rect 17036 17640 18387 17642
rect 17036 17584 18326 17640
rect 18382 17584 18387 17640
rect 17036 17582 18387 17584
rect 13445 17579 13511 17582
rect 12893 17506 12959 17509
rect 16760 17506 16820 17582
rect 18321 17579 18387 17582
rect 18505 17642 18571 17645
rect 20621 17642 20687 17645
rect 18505 17640 20687 17642
rect 18505 17584 18510 17640
rect 18566 17584 20626 17640
rect 20682 17584 20687 17640
rect 18505 17582 20687 17584
rect 18505 17579 18571 17582
rect 20621 17579 20687 17582
rect 24761 17642 24827 17645
rect 26374 17642 26434 17718
rect 27470 17716 27476 17718
rect 27540 17716 27546 17780
rect 27705 17778 27771 17781
rect 28625 17778 28691 17781
rect 28758 17778 28764 17780
rect 27705 17776 28764 17778
rect 27705 17720 27710 17776
rect 27766 17720 28630 17776
rect 28686 17720 28764 17776
rect 27705 17718 28764 17720
rect 27705 17715 27771 17718
rect 28625 17715 28691 17718
rect 28758 17716 28764 17718
rect 28828 17716 28834 17780
rect 29361 17778 29427 17781
rect 30097 17778 30163 17781
rect 29361 17776 30163 17778
rect 29361 17720 29366 17776
rect 29422 17720 30102 17776
rect 30158 17720 30163 17776
rect 29361 17718 30163 17720
rect 29361 17715 29427 17718
rect 30097 17715 30163 17718
rect 24761 17640 26434 17642
rect 24761 17584 24766 17640
rect 24822 17584 26434 17640
rect 24761 17582 26434 17584
rect 26969 17642 27035 17645
rect 29678 17642 29684 17644
rect 26969 17640 29684 17642
rect 26969 17584 26974 17640
rect 27030 17584 29684 17640
rect 26969 17582 29684 17584
rect 24761 17579 24827 17582
rect 26969 17579 27035 17582
rect 29678 17580 29684 17582
rect 29748 17580 29754 17644
rect 32029 17642 32095 17645
rect 29824 17640 32095 17642
rect 29824 17584 32034 17640
rect 32090 17584 32095 17640
rect 29824 17582 32095 17584
rect 16941 17506 17007 17509
rect 12893 17504 16084 17506
rect 12893 17448 12898 17504
rect 12954 17448 16084 17504
rect 12893 17446 16084 17448
rect 16760 17504 17007 17506
rect 16760 17448 16946 17504
rect 17002 17448 17007 17504
rect 16760 17446 17007 17448
rect 12893 17443 12959 17446
rect 8628 17440 8944 17441
rect 8628 17376 8634 17440
rect 8698 17376 8714 17440
rect 8778 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8944 17440
rect 8628 17375 8944 17376
rect 16024 17373 16084 17446
rect 16941 17443 17007 17446
rect 17125 17506 17191 17509
rect 24853 17506 24919 17509
rect 26785 17506 26851 17509
rect 17125 17504 23812 17506
rect 17125 17448 17130 17504
rect 17186 17448 23812 17504
rect 17125 17446 23812 17448
rect 17125 17443 17191 17446
rect 16310 17440 16626 17441
rect 16310 17376 16316 17440
rect 16380 17376 16396 17440
rect 16460 17376 16476 17440
rect 16540 17376 16556 17440
rect 16620 17376 16626 17440
rect 16310 17375 16626 17376
rect 12617 17370 12683 17373
rect 13077 17370 13143 17373
rect 15837 17370 15903 17373
rect 12617 17368 15903 17370
rect 12617 17312 12622 17368
rect 12678 17312 13082 17368
rect 13138 17312 15842 17368
rect 15898 17312 15903 17368
rect 12617 17310 15903 17312
rect 12617 17307 12683 17310
rect 13077 17307 13143 17310
rect 15837 17307 15903 17310
rect 16021 17368 16087 17373
rect 16021 17312 16026 17368
rect 16082 17312 16087 17368
rect 16021 17307 16087 17312
rect 16941 17370 17007 17373
rect 17166 17370 17172 17372
rect 16941 17368 17172 17370
rect 16941 17312 16946 17368
rect 17002 17312 17172 17368
rect 16941 17310 17172 17312
rect 16941 17307 17007 17310
rect 17166 17308 17172 17310
rect 17236 17308 17242 17372
rect 17309 17370 17375 17373
rect 23565 17370 23631 17373
rect 17309 17368 23631 17370
rect 17309 17312 17314 17368
rect 17370 17312 23570 17368
rect 23626 17312 23631 17368
rect 17309 17310 23631 17312
rect 17309 17307 17375 17310
rect 23565 17307 23631 17310
rect 10910 17172 10916 17236
rect 10980 17234 10986 17236
rect 23381 17234 23447 17237
rect 10980 17232 23447 17234
rect 10980 17176 23386 17232
rect 23442 17176 23447 17232
rect 10980 17174 23447 17176
rect 10980 17172 10986 17174
rect 23381 17171 23447 17174
rect 0 17008 800 17128
rect 10409 17098 10475 17101
rect 14549 17098 14615 17101
rect 15745 17098 15811 17101
rect 16573 17098 16639 17101
rect 23197 17098 23263 17101
rect 10409 17096 15578 17098
rect 10409 17040 10414 17096
rect 10470 17040 14554 17096
rect 14610 17040 15578 17096
rect 10409 17038 15578 17040
rect 10409 17035 10475 17038
rect 14549 17035 14615 17038
rect 10501 16964 10567 16965
rect 10501 16962 10548 16964
rect 10456 16960 10548 16962
rect 10456 16904 10506 16960
rect 10456 16902 10548 16904
rect 10501 16900 10548 16902
rect 10612 16900 10618 16964
rect 15518 16962 15578 17038
rect 15745 17096 16639 17098
rect 15745 17040 15750 17096
rect 15806 17040 16578 17096
rect 16634 17040 16639 17096
rect 15745 17038 16639 17040
rect 15745 17035 15811 17038
rect 16573 17035 16639 17038
rect 17174 17096 23263 17098
rect 17174 17040 23202 17096
rect 23258 17040 23263 17096
rect 17174 17038 23263 17040
rect 23752 17098 23812 17446
rect 24853 17504 26851 17506
rect 24853 17448 24858 17504
rect 24914 17448 26790 17504
rect 26846 17448 26851 17504
rect 24853 17446 26851 17448
rect 24853 17443 24919 17446
rect 26785 17443 26851 17446
rect 27102 17444 27108 17508
rect 27172 17506 27178 17508
rect 27429 17506 27495 17509
rect 27172 17504 27495 17506
rect 27172 17448 27434 17504
rect 27490 17448 27495 17504
rect 27172 17446 27495 17448
rect 27172 17444 27178 17446
rect 27429 17443 27495 17446
rect 27654 17444 27660 17508
rect 27724 17506 27730 17508
rect 28073 17506 28139 17509
rect 27724 17504 28139 17506
rect 27724 17448 28078 17504
rect 28134 17448 28139 17504
rect 27724 17446 28139 17448
rect 27724 17444 27730 17446
rect 28073 17443 28139 17446
rect 28257 17506 28323 17509
rect 28574 17506 28580 17508
rect 28257 17504 28580 17506
rect 28257 17448 28262 17504
rect 28318 17448 28580 17504
rect 28257 17446 28580 17448
rect 28257 17443 28323 17446
rect 28574 17444 28580 17446
rect 28644 17506 28650 17508
rect 29824 17506 29884 17582
rect 32029 17579 32095 17582
rect 32206 17506 33006 17536
rect 28644 17446 29884 17506
rect 32078 17446 33006 17506
rect 28644 17444 28650 17446
rect 23992 17440 24308 17441
rect 23992 17376 23998 17440
rect 24062 17376 24078 17440
rect 24142 17376 24158 17440
rect 24222 17376 24238 17440
rect 24302 17376 24308 17440
rect 23992 17375 24308 17376
rect 31674 17440 31990 17441
rect 31674 17376 31680 17440
rect 31744 17376 31760 17440
rect 31824 17376 31840 17440
rect 31904 17376 31920 17440
rect 31984 17376 31990 17440
rect 31674 17375 31990 17376
rect 24669 17370 24735 17373
rect 30230 17370 30236 17372
rect 24669 17368 30236 17370
rect 24669 17312 24674 17368
rect 24730 17312 30236 17368
rect 24669 17310 30236 17312
rect 24669 17307 24735 17310
rect 30230 17308 30236 17310
rect 30300 17308 30306 17372
rect 30465 17370 30531 17373
rect 30649 17370 30715 17373
rect 30465 17368 30715 17370
rect 30465 17312 30470 17368
rect 30526 17312 30654 17368
rect 30710 17312 30715 17368
rect 30465 17310 30715 17312
rect 30465 17307 30531 17310
rect 30649 17307 30715 17310
rect 24853 17234 24919 17237
rect 26233 17234 26299 17237
rect 24853 17232 26299 17234
rect 24853 17176 24858 17232
rect 24914 17176 26238 17232
rect 26294 17176 26299 17232
rect 24853 17174 26299 17176
rect 24853 17171 24919 17174
rect 26233 17171 26299 17174
rect 26366 17172 26372 17236
rect 26436 17234 26442 17236
rect 26877 17234 26943 17237
rect 28533 17234 28599 17237
rect 26436 17232 28599 17234
rect 26436 17176 26882 17232
rect 26938 17176 28538 17232
rect 28594 17176 28599 17232
rect 26436 17174 28599 17176
rect 26436 17172 26442 17174
rect 26877 17171 26943 17174
rect 28533 17171 28599 17174
rect 28901 17234 28967 17237
rect 32078 17234 32138 17446
rect 32206 17416 33006 17446
rect 28901 17232 32138 17234
rect 28901 17176 28906 17232
rect 28962 17176 32138 17232
rect 28901 17174 32138 17176
rect 28901 17171 28967 17174
rect 29177 17098 29243 17101
rect 23752 17096 29243 17098
rect 23752 17040 29182 17096
rect 29238 17040 29243 17096
rect 23752 17038 29243 17040
rect 15929 16962 15995 16965
rect 15518 16960 15995 16962
rect 15518 16904 15934 16960
rect 15990 16904 15995 16960
rect 15518 16902 15995 16904
rect 10501 16899 10567 16900
rect 15929 16899 15995 16902
rect 16062 16900 16068 16964
rect 16132 16962 16138 16964
rect 17174 16962 17234 17038
rect 23197 17035 23263 17038
rect 29177 17035 29243 17038
rect 30465 17098 30531 17101
rect 30741 17098 30807 17101
rect 30465 17096 30807 17098
rect 30465 17040 30470 17096
rect 30526 17040 30746 17096
rect 30802 17040 30807 17096
rect 30465 17038 30807 17040
rect 30465 17035 30531 17038
rect 30741 17035 30807 17038
rect 31518 17036 31524 17100
rect 31588 17098 31594 17100
rect 31661 17098 31727 17101
rect 31588 17096 31727 17098
rect 31588 17040 31666 17096
rect 31722 17040 31727 17096
rect 31588 17038 31727 17040
rect 31588 17036 31594 17038
rect 31661 17035 31727 17038
rect 16132 16902 17234 16962
rect 16132 16900 16138 16902
rect 17350 16900 17356 16964
rect 17420 16962 17426 16964
rect 17493 16962 17559 16965
rect 17420 16960 17559 16962
rect 17420 16904 17498 16960
rect 17554 16904 17559 16960
rect 17420 16902 17559 16904
rect 17420 16900 17426 16902
rect 17493 16899 17559 16902
rect 17861 16962 17927 16965
rect 18413 16962 18479 16965
rect 19793 16962 19859 16965
rect 17861 16960 17970 16962
rect 17861 16904 17866 16960
rect 17922 16904 17970 16960
rect 17861 16899 17970 16904
rect 18413 16960 19859 16962
rect 18413 16904 18418 16960
rect 18474 16904 19798 16960
rect 19854 16904 19859 16960
rect 18413 16902 19859 16904
rect 18413 16899 18479 16902
rect 19793 16899 19859 16902
rect 22461 16962 22527 16965
rect 25497 16962 25563 16965
rect 25998 16962 26004 16964
rect 22461 16960 26004 16962
rect 22461 16904 22466 16960
rect 22522 16904 25502 16960
rect 25558 16904 26004 16960
rect 22461 16902 26004 16904
rect 22461 16899 22527 16902
rect 25497 16899 25563 16902
rect 25998 16900 26004 16902
rect 26068 16900 26074 16964
rect 26693 16962 26759 16965
rect 26918 16962 26924 16964
rect 26693 16960 26924 16962
rect 26693 16904 26698 16960
rect 26754 16904 26924 16960
rect 26693 16902 26924 16904
rect 26693 16899 26759 16902
rect 26918 16900 26924 16902
rect 26988 16900 26994 16964
rect 29126 16962 29132 16964
rect 28996 16902 29132 16962
rect 4787 16896 5103 16897
rect 4787 16832 4793 16896
rect 4857 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5103 16896
rect 4787 16831 5103 16832
rect 12469 16896 12785 16897
rect 12469 16832 12475 16896
rect 12539 16832 12555 16896
rect 12619 16832 12635 16896
rect 12699 16832 12715 16896
rect 12779 16832 12785 16896
rect 12469 16831 12785 16832
rect 14089 16826 14155 16829
rect 14457 16826 14523 16829
rect 17769 16826 17835 16829
rect 14089 16824 17835 16826
rect 14089 16768 14094 16824
rect 14150 16768 14462 16824
rect 14518 16768 17774 16824
rect 17830 16768 17835 16824
rect 14089 16766 17835 16768
rect 17910 16826 17970 16899
rect 20151 16896 20467 16897
rect 20151 16832 20157 16896
rect 20221 16832 20237 16896
rect 20301 16832 20317 16896
rect 20381 16832 20397 16896
rect 20461 16832 20467 16896
rect 20151 16831 20467 16832
rect 27833 16896 28149 16897
rect 27833 16832 27839 16896
rect 27903 16832 27919 16896
rect 27983 16832 27999 16896
rect 28063 16832 28079 16896
rect 28143 16832 28149 16896
rect 27833 16831 28149 16832
rect 19977 16826 20043 16829
rect 17910 16824 20043 16826
rect 17910 16768 19982 16824
rect 20038 16768 20043 16824
rect 17910 16766 20043 16768
rect 14089 16763 14155 16766
rect 14457 16763 14523 16766
rect 17769 16763 17835 16766
rect 19977 16763 20043 16766
rect 22277 16826 22343 16829
rect 23749 16828 23815 16829
rect 22277 16824 23260 16826
rect 22277 16768 22282 16824
rect 22338 16768 23260 16824
rect 22277 16766 23260 16768
rect 22277 16763 22343 16766
rect 12709 16690 12775 16693
rect 14181 16690 14247 16693
rect 12709 16688 14247 16690
rect 12709 16632 12714 16688
rect 12770 16632 14186 16688
rect 14242 16632 14247 16688
rect 12709 16630 14247 16632
rect 12709 16627 12775 16630
rect 14181 16627 14247 16630
rect 14365 16690 14431 16693
rect 20529 16690 20595 16693
rect 22369 16690 22435 16693
rect 14365 16688 22435 16690
rect 14365 16632 14370 16688
rect 14426 16632 20534 16688
rect 20590 16632 22374 16688
rect 22430 16632 22435 16688
rect 14365 16630 22435 16632
rect 14365 16627 14431 16630
rect 20529 16627 20595 16630
rect 22369 16627 22435 16630
rect 22737 16690 22803 16693
rect 23013 16690 23079 16693
rect 22737 16688 23079 16690
rect 22737 16632 22742 16688
rect 22798 16632 23018 16688
rect 23074 16632 23079 16688
rect 22737 16630 23079 16632
rect 23200 16690 23260 16766
rect 23749 16824 23796 16828
rect 23860 16826 23866 16828
rect 24669 16826 24735 16829
rect 25313 16826 25379 16829
rect 26969 16828 27035 16829
rect 23749 16768 23754 16824
rect 23749 16764 23796 16768
rect 23860 16766 23906 16826
rect 24669 16824 25379 16826
rect 24669 16768 24674 16824
rect 24730 16768 25318 16824
rect 25374 16768 25379 16824
rect 24669 16766 25379 16768
rect 23860 16764 23866 16766
rect 23749 16763 23815 16764
rect 24669 16763 24735 16766
rect 25313 16763 25379 16766
rect 26918 16764 26924 16828
rect 26988 16826 27035 16828
rect 27429 16826 27495 16829
rect 26988 16824 27080 16826
rect 27030 16768 27080 16824
rect 26988 16766 27080 16768
rect 27429 16824 27768 16826
rect 27429 16768 27434 16824
rect 27490 16768 27768 16824
rect 27429 16766 27768 16768
rect 26988 16764 27035 16766
rect 26969 16763 27035 16764
rect 27429 16763 27495 16766
rect 23606 16690 23612 16692
rect 23200 16630 23612 16690
rect 22737 16627 22803 16630
rect 23013 16627 23079 16630
rect 23606 16628 23612 16630
rect 23676 16690 23682 16692
rect 26509 16690 26575 16693
rect 27429 16690 27495 16693
rect 23676 16688 27495 16690
rect 23676 16632 26514 16688
rect 26570 16632 27434 16688
rect 27490 16632 27495 16688
rect 23676 16630 27495 16632
rect 23676 16628 23682 16630
rect 26509 16627 26575 16630
rect 27429 16627 27495 16630
rect 10726 16492 10732 16556
rect 10796 16554 10802 16556
rect 11145 16554 11211 16557
rect 12157 16556 12223 16557
rect 12157 16554 12204 16556
rect 10796 16552 11211 16554
rect 10796 16496 11150 16552
rect 11206 16496 11211 16552
rect 10796 16494 11211 16496
rect 12112 16552 12204 16554
rect 12112 16496 12162 16552
rect 12112 16494 12204 16496
rect 10796 16492 10802 16494
rect 11145 16491 11211 16494
rect 12157 16492 12204 16494
rect 12268 16492 12274 16556
rect 12985 16554 13051 16557
rect 21173 16554 21239 16557
rect 12985 16552 21239 16554
rect 12985 16496 12990 16552
rect 13046 16496 21178 16552
rect 21234 16496 21239 16552
rect 12985 16494 21239 16496
rect 12157 16491 12223 16492
rect 12985 16491 13051 16494
rect 21173 16491 21239 16494
rect 23013 16554 23079 16557
rect 24025 16554 24091 16557
rect 23013 16552 24091 16554
rect 23013 16496 23018 16552
rect 23074 16496 24030 16552
rect 24086 16496 24091 16552
rect 23013 16494 24091 16496
rect 23013 16491 23079 16494
rect 24025 16491 24091 16494
rect 25405 16552 25471 16557
rect 25405 16496 25410 16552
rect 25466 16496 25471 16552
rect 25405 16491 25471 16496
rect 25681 16554 25747 16557
rect 25814 16554 25820 16556
rect 25681 16552 25820 16554
rect 25681 16496 25686 16552
rect 25742 16496 25820 16552
rect 25681 16494 25820 16496
rect 25681 16491 25747 16494
rect 25814 16492 25820 16494
rect 25884 16492 25890 16556
rect 27708 16554 27768 16766
rect 28390 16764 28396 16828
rect 28460 16826 28466 16828
rect 28533 16826 28599 16829
rect 28996 16826 29056 16902
rect 29126 16900 29132 16902
rect 29196 16900 29202 16964
rect 29269 16962 29335 16965
rect 30468 16962 30528 17035
rect 29269 16960 30528 16962
rect 29269 16904 29274 16960
rect 29330 16904 30528 16960
rect 29269 16902 30528 16904
rect 29269 16899 29335 16902
rect 30598 16900 30604 16964
rect 30668 16962 30674 16964
rect 32029 16962 32095 16965
rect 30668 16960 32095 16962
rect 30668 16904 32034 16960
rect 32090 16904 32095 16960
rect 30668 16902 32095 16904
rect 30668 16900 30674 16902
rect 32029 16899 32095 16902
rect 28460 16824 28599 16826
rect 28460 16768 28538 16824
rect 28594 16768 28599 16824
rect 28460 16766 28599 16768
rect 28460 16764 28466 16766
rect 28533 16763 28599 16766
rect 28812 16766 29056 16826
rect 28165 16690 28231 16693
rect 28390 16690 28396 16692
rect 28165 16688 28396 16690
rect 28165 16632 28170 16688
rect 28226 16632 28396 16688
rect 28165 16630 28396 16632
rect 28165 16627 28231 16630
rect 28390 16628 28396 16630
rect 28460 16628 28466 16692
rect 28812 16554 28872 16766
rect 29126 16764 29132 16828
rect 29196 16826 29202 16828
rect 29545 16826 29611 16829
rect 29196 16824 29611 16826
rect 29196 16768 29550 16824
rect 29606 16768 29611 16824
rect 29196 16766 29611 16768
rect 29196 16764 29202 16766
rect 29545 16763 29611 16766
rect 32206 16736 33006 16856
rect 28993 16690 29059 16693
rect 29494 16690 29500 16692
rect 28993 16688 29500 16690
rect 28993 16632 28998 16688
rect 29054 16632 29500 16688
rect 28993 16630 29500 16632
rect 28993 16627 29059 16630
rect 29494 16628 29500 16630
rect 29564 16628 29570 16692
rect 30046 16690 30052 16692
rect 29640 16630 30052 16690
rect 27708 16494 28872 16554
rect 28942 16492 28948 16556
rect 29012 16554 29018 16556
rect 29361 16554 29427 16557
rect 29012 16552 29427 16554
rect 29012 16496 29366 16552
rect 29422 16496 29427 16552
rect 29012 16494 29427 16496
rect 29012 16492 29018 16494
rect 29361 16491 29427 16494
rect 29494 16492 29500 16556
rect 29564 16554 29570 16556
rect 29640 16554 29700 16630
rect 30046 16628 30052 16630
rect 30116 16628 30122 16692
rect 30966 16628 30972 16692
rect 31036 16690 31042 16692
rect 31293 16690 31359 16693
rect 31036 16688 31359 16690
rect 31036 16632 31298 16688
rect 31354 16632 31359 16688
rect 31036 16630 31359 16632
rect 31036 16628 31042 16630
rect 31293 16627 31359 16630
rect 29564 16494 29700 16554
rect 29564 16492 29570 16494
rect 30046 16492 30052 16556
rect 30116 16554 30122 16556
rect 30373 16554 30439 16557
rect 30116 16552 30439 16554
rect 30116 16496 30378 16552
rect 30434 16496 30439 16552
rect 30116 16494 30439 16496
rect 30116 16492 30122 16494
rect 30373 16491 30439 16494
rect 25408 16421 25468 16491
rect 12617 16418 12683 16421
rect 14457 16418 14523 16421
rect 12617 16416 14523 16418
rect 12617 16360 12622 16416
rect 12678 16360 14462 16416
rect 14518 16360 14523 16416
rect 12617 16358 14523 16360
rect 12617 16355 12683 16358
rect 14457 16355 14523 16358
rect 14733 16418 14799 16421
rect 15837 16418 15903 16421
rect 14733 16416 15903 16418
rect 14733 16360 14738 16416
rect 14794 16360 15842 16416
rect 15898 16360 15903 16416
rect 14733 16358 15903 16360
rect 14733 16355 14799 16358
rect 15837 16355 15903 16358
rect 16021 16416 16087 16421
rect 16021 16360 16026 16416
rect 16082 16360 16087 16416
rect 16021 16355 16087 16360
rect 16757 16416 16823 16421
rect 16757 16360 16762 16416
rect 16818 16360 16823 16416
rect 16757 16355 16823 16360
rect 16941 16418 17007 16421
rect 24853 16418 24919 16421
rect 25037 16418 25103 16421
rect 16941 16416 23858 16418
rect 16941 16360 16946 16416
rect 17002 16360 23858 16416
rect 16941 16358 23858 16360
rect 16941 16355 17007 16358
rect 8628 16352 8944 16353
rect 0 16282 800 16312
rect 8628 16288 8634 16352
rect 8698 16288 8714 16352
rect 8778 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8944 16352
rect 8628 16287 8944 16288
rect 1577 16282 1643 16285
rect 15193 16284 15259 16285
rect 0 16280 1643 16282
rect 0 16224 1582 16280
rect 1638 16224 1643 16280
rect 0 16222 1643 16224
rect 0 16192 800 16222
rect 1577 16219 1643 16222
rect 15142 16220 15148 16284
rect 15212 16282 15259 16284
rect 15377 16282 15443 16285
rect 16024 16282 16084 16355
rect 16310 16352 16626 16353
rect 16310 16288 16316 16352
rect 16380 16288 16396 16352
rect 16460 16288 16476 16352
rect 16540 16288 16556 16352
rect 16620 16288 16626 16352
rect 16310 16287 16626 16288
rect 15212 16280 15304 16282
rect 15254 16224 15304 16280
rect 15212 16222 15304 16224
rect 15377 16280 16084 16282
rect 15377 16224 15382 16280
rect 15438 16224 16084 16280
rect 15377 16222 16084 16224
rect 16760 16282 16820 16355
rect 18413 16282 18479 16285
rect 19057 16284 19123 16285
rect 19006 16282 19012 16284
rect 16760 16280 18479 16282
rect 16760 16224 18418 16280
rect 18474 16224 18479 16280
rect 16760 16222 18479 16224
rect 18966 16222 19012 16282
rect 19076 16280 19123 16284
rect 19118 16224 19123 16280
rect 15212 16220 15259 16222
rect 15193 16219 15259 16220
rect 15377 16219 15443 16222
rect 18413 16219 18479 16222
rect 19006 16220 19012 16222
rect 19076 16220 19123 16224
rect 19057 16219 19123 16220
rect 19609 16282 19675 16285
rect 19609 16280 22524 16282
rect 19609 16224 19614 16280
rect 19670 16224 22524 16280
rect 19609 16222 22524 16224
rect 19609 16219 19675 16222
rect 11605 16146 11671 16149
rect 22277 16146 22343 16149
rect 11605 16144 22343 16146
rect 11605 16088 11610 16144
rect 11666 16088 22282 16144
rect 22338 16088 22343 16144
rect 11605 16086 22343 16088
rect 22464 16146 22524 16222
rect 23657 16146 23723 16149
rect 22464 16144 23723 16146
rect 22464 16088 23662 16144
rect 23718 16088 23723 16144
rect 22464 16086 23723 16088
rect 23798 16146 23858 16358
rect 24853 16416 25103 16418
rect 24853 16360 24858 16416
rect 24914 16360 25042 16416
rect 25098 16360 25103 16416
rect 24853 16358 25103 16360
rect 24853 16355 24919 16358
rect 25037 16355 25103 16358
rect 25405 16416 25471 16421
rect 25405 16360 25410 16416
rect 25466 16360 25471 16416
rect 25405 16355 25471 16360
rect 26877 16418 26943 16421
rect 29269 16418 29335 16421
rect 29545 16418 29611 16421
rect 26877 16416 29611 16418
rect 26877 16360 26882 16416
rect 26938 16360 29274 16416
rect 29330 16360 29550 16416
rect 29606 16360 29611 16416
rect 26877 16358 29611 16360
rect 26877 16355 26943 16358
rect 29269 16355 29335 16358
rect 29545 16355 29611 16358
rect 23992 16352 24308 16353
rect 23992 16288 23998 16352
rect 24062 16288 24078 16352
rect 24142 16288 24158 16352
rect 24222 16288 24238 16352
rect 24302 16288 24308 16352
rect 23992 16287 24308 16288
rect 31674 16352 31990 16353
rect 31674 16288 31680 16352
rect 31744 16288 31760 16352
rect 31824 16288 31840 16352
rect 31904 16288 31920 16352
rect 31984 16288 31990 16352
rect 31674 16287 31990 16288
rect 28073 16282 28139 16285
rect 24810 16280 28139 16282
rect 24810 16224 28078 16280
rect 28134 16224 28139 16280
rect 24810 16222 28139 16224
rect 24810 16146 24870 16222
rect 28073 16219 28139 16222
rect 28441 16282 28507 16285
rect 28993 16282 29059 16285
rect 28441 16280 29059 16282
rect 28441 16224 28446 16280
rect 28502 16224 28998 16280
rect 29054 16224 29059 16280
rect 28441 16222 29059 16224
rect 28441 16219 28507 16222
rect 28993 16219 29059 16222
rect 23798 16086 24870 16146
rect 26693 16146 26759 16149
rect 30649 16146 30715 16149
rect 26693 16144 30715 16146
rect 26693 16088 26698 16144
rect 26754 16088 30654 16144
rect 30710 16088 30715 16144
rect 26693 16086 30715 16088
rect 11605 16083 11671 16086
rect 22277 16083 22343 16086
rect 23657 16083 23723 16086
rect 26693 16083 26759 16086
rect 30649 16083 30715 16086
rect 31293 16146 31359 16149
rect 32206 16146 33006 16176
rect 31293 16144 33006 16146
rect 31293 16088 31298 16144
rect 31354 16088 33006 16144
rect 31293 16086 33006 16088
rect 31293 16083 31359 16086
rect 32206 16056 33006 16086
rect 14181 16010 14247 16013
rect 23289 16010 23355 16013
rect 14181 16008 23355 16010
rect 14181 15952 14186 16008
rect 14242 15952 23294 16008
rect 23350 15952 23355 16008
rect 14181 15950 23355 15952
rect 14181 15947 14247 15950
rect 23289 15947 23355 15950
rect 24853 16010 24919 16013
rect 25589 16010 25655 16013
rect 24853 16008 25655 16010
rect 24853 15952 24858 16008
rect 24914 15952 25594 16008
rect 25650 15952 25655 16008
rect 24853 15950 25655 15952
rect 24853 15947 24919 15950
rect 25589 15947 25655 15950
rect 26785 16010 26851 16013
rect 29085 16010 29151 16013
rect 29913 16010 29979 16013
rect 30741 16012 30807 16013
rect 30414 16010 30420 16012
rect 26785 16008 30420 16010
rect 26785 15952 26790 16008
rect 26846 15952 29090 16008
rect 29146 15952 29918 16008
rect 29974 15952 30420 16008
rect 26785 15950 30420 15952
rect 26785 15947 26851 15950
rect 29085 15947 29151 15950
rect 29913 15947 29979 15950
rect 30414 15948 30420 15950
rect 30484 15948 30490 16012
rect 30741 16010 30788 16012
rect 30696 16008 30788 16010
rect 30696 15952 30746 16008
rect 30696 15950 30788 15952
rect 30741 15948 30788 15950
rect 30852 15948 30858 16012
rect 30741 15947 30807 15948
rect 13353 15874 13419 15877
rect 18229 15874 18295 15877
rect 13353 15872 18295 15874
rect 13353 15816 13358 15872
rect 13414 15816 18234 15872
rect 18290 15816 18295 15872
rect 13353 15814 18295 15816
rect 13353 15811 13419 15814
rect 18229 15811 18295 15814
rect 18597 15874 18663 15877
rect 19609 15874 19675 15877
rect 18597 15872 19675 15874
rect 18597 15816 18602 15872
rect 18658 15816 19614 15872
rect 19670 15816 19675 15872
rect 18597 15814 19675 15816
rect 18597 15811 18663 15814
rect 19609 15811 19675 15814
rect 29177 15874 29243 15877
rect 32673 15874 32739 15877
rect 29177 15872 32739 15874
rect 29177 15816 29182 15872
rect 29238 15816 32678 15872
rect 32734 15816 32739 15872
rect 29177 15814 32739 15816
rect 29177 15811 29243 15814
rect 32673 15811 32739 15814
rect 4787 15808 5103 15809
rect 4787 15744 4793 15808
rect 4857 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5103 15808
rect 4787 15743 5103 15744
rect 12469 15808 12785 15809
rect 12469 15744 12475 15808
rect 12539 15744 12555 15808
rect 12619 15744 12635 15808
rect 12699 15744 12715 15808
rect 12779 15744 12785 15808
rect 12469 15743 12785 15744
rect 20151 15808 20467 15809
rect 20151 15744 20157 15808
rect 20221 15744 20237 15808
rect 20301 15744 20317 15808
rect 20381 15744 20397 15808
rect 20461 15744 20467 15808
rect 20151 15743 20467 15744
rect 27833 15808 28149 15809
rect 27833 15744 27839 15808
rect 27903 15744 27919 15808
rect 27983 15744 27999 15808
rect 28063 15744 28079 15808
rect 28143 15744 28149 15808
rect 27833 15743 28149 15744
rect 15285 15738 15351 15741
rect 16389 15738 16455 15741
rect 18229 15738 18295 15741
rect 15285 15736 16455 15738
rect 15285 15680 15290 15736
rect 15346 15680 16394 15736
rect 16450 15680 16455 15736
rect 15285 15678 16455 15680
rect 15285 15675 15351 15678
rect 16389 15675 16455 15678
rect 16530 15736 18295 15738
rect 16530 15680 18234 15736
rect 18290 15680 18295 15736
rect 16530 15678 18295 15680
rect 15193 15602 15259 15605
rect 16530 15602 16590 15678
rect 18229 15675 18295 15678
rect 18873 15738 18939 15741
rect 19885 15738 19951 15741
rect 18873 15736 19951 15738
rect 18873 15680 18878 15736
rect 18934 15680 19890 15736
rect 19946 15680 19951 15736
rect 18873 15678 19951 15680
rect 18873 15675 18939 15678
rect 19885 15675 19951 15678
rect 21081 15738 21147 15741
rect 24485 15738 24551 15741
rect 32121 15738 32187 15741
rect 21081 15736 24551 15738
rect 21081 15680 21086 15736
rect 21142 15680 24490 15736
rect 24546 15680 24551 15736
rect 21081 15678 24551 15680
rect 21081 15675 21147 15678
rect 24485 15675 24551 15678
rect 28214 15736 32187 15738
rect 28214 15680 32126 15736
rect 32182 15680 32187 15736
rect 28214 15678 32187 15680
rect 15193 15600 16590 15602
rect 15193 15544 15198 15600
rect 15254 15544 16590 15600
rect 15193 15542 16590 15544
rect 15193 15539 15259 15542
rect 16798 15540 16804 15604
rect 16868 15602 16874 15604
rect 17493 15602 17559 15605
rect 16868 15600 17559 15602
rect 16868 15544 17498 15600
rect 17554 15544 17559 15600
rect 16868 15542 17559 15544
rect 16868 15540 16874 15542
rect 17493 15539 17559 15542
rect 17769 15602 17835 15605
rect 23933 15602 23999 15605
rect 28214 15602 28274 15678
rect 32121 15675 32187 15678
rect 17769 15600 28274 15602
rect 17769 15544 17774 15600
rect 17830 15544 23938 15600
rect 23994 15544 28274 15600
rect 17769 15542 28274 15544
rect 28625 15602 28691 15605
rect 29126 15602 29132 15604
rect 28625 15600 29132 15602
rect 28625 15544 28630 15600
rect 28686 15544 29132 15600
rect 28625 15542 29132 15544
rect 17769 15539 17835 15542
rect 23933 15539 23999 15542
rect 28625 15539 28691 15542
rect 29126 15540 29132 15542
rect 29196 15540 29202 15604
rect 0 15466 800 15496
rect 1577 15466 1643 15469
rect 0 15464 1643 15466
rect 0 15408 1582 15464
rect 1638 15408 1643 15464
rect 0 15406 1643 15408
rect 0 15376 800 15406
rect 1577 15403 1643 15406
rect 12249 15466 12315 15469
rect 24025 15466 24091 15469
rect 12249 15464 24091 15466
rect 12249 15408 12254 15464
rect 12310 15408 24030 15464
rect 24086 15408 24091 15464
rect 12249 15406 24091 15408
rect 12249 15403 12315 15406
rect 24025 15403 24091 15406
rect 24526 15404 24532 15468
rect 24596 15466 24602 15468
rect 26049 15466 26115 15469
rect 24596 15464 26115 15466
rect 24596 15408 26054 15464
rect 26110 15408 26115 15464
rect 24596 15406 26115 15408
rect 24596 15404 24602 15406
rect 26049 15403 26115 15406
rect 26734 15404 26740 15468
rect 26804 15466 26810 15468
rect 26877 15466 26943 15469
rect 29269 15466 29335 15469
rect 26804 15464 29335 15466
rect 26804 15408 26882 15464
rect 26938 15408 29274 15464
rect 29330 15408 29335 15464
rect 26804 15406 29335 15408
rect 26804 15404 26810 15406
rect 26877 15403 26943 15406
rect 29269 15403 29335 15406
rect 30741 15466 30807 15469
rect 32206 15466 33006 15496
rect 30741 15464 33006 15466
rect 30741 15408 30746 15464
rect 30802 15408 33006 15464
rect 30741 15406 33006 15408
rect 30741 15403 30807 15406
rect 32206 15376 33006 15406
rect 11646 15268 11652 15332
rect 11716 15330 11722 15332
rect 16062 15330 16068 15332
rect 11716 15270 16068 15330
rect 11716 15268 11722 15270
rect 16062 15268 16068 15270
rect 16132 15268 16138 15332
rect 17902 15268 17908 15332
rect 17972 15330 17978 15332
rect 21398 15330 21404 15332
rect 17972 15270 21404 15330
rect 17972 15268 17978 15270
rect 21398 15268 21404 15270
rect 21468 15268 21474 15332
rect 24894 15268 24900 15332
rect 24964 15330 24970 15332
rect 25037 15330 25103 15333
rect 24964 15328 25103 15330
rect 24964 15272 25042 15328
rect 25098 15272 25103 15328
rect 24964 15270 25103 15272
rect 24964 15268 24970 15270
rect 25037 15267 25103 15270
rect 25814 15268 25820 15332
rect 25884 15330 25890 15332
rect 25957 15330 26023 15333
rect 25884 15328 26023 15330
rect 25884 15272 25962 15328
rect 26018 15272 26023 15328
rect 25884 15270 26023 15272
rect 25884 15268 25890 15270
rect 25957 15267 26023 15270
rect 27889 15330 27955 15333
rect 29637 15330 29703 15333
rect 27889 15328 29703 15330
rect 27889 15272 27894 15328
rect 27950 15272 29642 15328
rect 29698 15272 29703 15328
rect 27889 15270 29703 15272
rect 27889 15267 27955 15270
rect 29637 15267 29703 15270
rect 30230 15268 30236 15332
rect 30300 15330 30306 15332
rect 30465 15330 30531 15333
rect 30300 15328 30531 15330
rect 30300 15272 30470 15328
rect 30526 15272 30531 15328
rect 30300 15270 30531 15272
rect 30300 15268 30306 15270
rect 30465 15267 30531 15270
rect 8628 15264 8944 15265
rect 8628 15200 8634 15264
rect 8698 15200 8714 15264
rect 8778 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8944 15264
rect 8628 15199 8944 15200
rect 16310 15264 16626 15265
rect 16310 15200 16316 15264
rect 16380 15200 16396 15264
rect 16460 15200 16476 15264
rect 16540 15200 16556 15264
rect 16620 15200 16626 15264
rect 16310 15199 16626 15200
rect 23992 15264 24308 15265
rect 23992 15200 23998 15264
rect 24062 15200 24078 15264
rect 24142 15200 24158 15264
rect 24222 15200 24238 15264
rect 24302 15200 24308 15264
rect 23992 15199 24308 15200
rect 31674 15264 31990 15265
rect 31674 15200 31680 15264
rect 31744 15200 31760 15264
rect 31824 15200 31840 15264
rect 31904 15200 31920 15264
rect 31984 15200 31990 15264
rect 31674 15199 31990 15200
rect 16757 15194 16823 15197
rect 20713 15194 20779 15197
rect 16757 15192 20779 15194
rect 16757 15136 16762 15192
rect 16818 15136 20718 15192
rect 20774 15136 20779 15192
rect 16757 15134 20779 15136
rect 16757 15131 16823 15134
rect 20713 15131 20779 15134
rect 21398 15132 21404 15196
rect 21468 15194 21474 15196
rect 21541 15194 21607 15197
rect 21468 15192 21607 15194
rect 21468 15136 21546 15192
rect 21602 15136 21607 15192
rect 21468 15134 21607 15136
rect 21468 15132 21474 15134
rect 21541 15131 21607 15134
rect 25630 15132 25636 15196
rect 25700 15194 25706 15196
rect 29177 15194 29243 15197
rect 31518 15194 31524 15196
rect 25700 15134 28826 15194
rect 25700 15132 25706 15134
rect 13905 15058 13971 15061
rect 17769 15058 17835 15061
rect 13905 15056 17835 15058
rect 13905 15000 13910 15056
rect 13966 15000 17774 15056
rect 17830 15000 17835 15056
rect 13905 14998 17835 15000
rect 13905 14995 13971 14998
rect 17769 14995 17835 14998
rect 18045 15058 18111 15061
rect 20805 15058 20871 15061
rect 18045 15056 20871 15058
rect 18045 15000 18050 15056
rect 18106 15000 20810 15056
rect 20866 15000 20871 15056
rect 18045 14998 20871 15000
rect 18045 14995 18111 14998
rect 20805 14995 20871 14998
rect 22461 15058 22527 15061
rect 28625 15058 28691 15061
rect 22461 15056 28691 15058
rect 22461 15000 22466 15056
rect 22522 15000 28630 15056
rect 28686 15000 28691 15056
rect 22461 14998 28691 15000
rect 28766 15058 28826 15134
rect 29177 15192 31524 15194
rect 29177 15136 29182 15192
rect 29238 15136 31524 15192
rect 29177 15134 31524 15136
rect 29177 15131 29243 15134
rect 31518 15132 31524 15134
rect 31588 15132 31594 15196
rect 30005 15058 30071 15061
rect 28766 15056 30071 15058
rect 28766 15000 30010 15056
rect 30066 15000 30071 15056
rect 28766 14998 30071 15000
rect 22461 14995 22527 14998
rect 28625 14995 28691 14998
rect 30005 14995 30071 14998
rect 12065 14922 12131 14925
rect 20989 14922 21055 14925
rect 12065 14920 21055 14922
rect 12065 14864 12070 14920
rect 12126 14864 20994 14920
rect 21050 14864 21055 14920
rect 12065 14862 21055 14864
rect 12065 14859 12131 14862
rect 20989 14859 21055 14862
rect 26049 14922 26115 14925
rect 30465 14922 30531 14925
rect 26049 14920 30531 14922
rect 26049 14864 26054 14920
rect 26110 14864 30470 14920
rect 30526 14864 30531 14920
rect 26049 14862 30531 14864
rect 26049 14859 26115 14862
rect 30465 14859 30531 14862
rect 18045 14786 18111 14789
rect 14598 14784 18111 14786
rect 14598 14728 18050 14784
rect 18106 14728 18111 14784
rect 14598 14726 18111 14728
rect 4787 14720 5103 14721
rect 0 14560 800 14680
rect 4787 14656 4793 14720
rect 4857 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5103 14720
rect 4787 14655 5103 14656
rect 12469 14720 12785 14721
rect 12469 14656 12475 14720
rect 12539 14656 12555 14720
rect 12619 14656 12635 14720
rect 12699 14656 12715 14720
rect 12779 14656 12785 14720
rect 12469 14655 12785 14656
rect 11973 14514 12039 14517
rect 14598 14514 14658 14726
rect 18045 14723 18111 14726
rect 20846 14724 20852 14788
rect 20916 14786 20922 14788
rect 21541 14786 21607 14789
rect 20916 14784 21607 14786
rect 20916 14728 21546 14784
rect 21602 14728 21607 14784
rect 20916 14726 21607 14728
rect 20916 14724 20922 14726
rect 21541 14723 21607 14726
rect 28625 14786 28691 14789
rect 29310 14786 29316 14788
rect 28625 14784 29316 14786
rect 28625 14728 28630 14784
rect 28686 14728 29316 14784
rect 28625 14726 29316 14728
rect 28625 14723 28691 14726
rect 29310 14724 29316 14726
rect 29380 14724 29386 14788
rect 20151 14720 20467 14721
rect 20151 14656 20157 14720
rect 20221 14656 20237 14720
rect 20301 14656 20317 14720
rect 20381 14656 20397 14720
rect 20461 14656 20467 14720
rect 20151 14655 20467 14656
rect 27833 14720 28149 14721
rect 27833 14656 27839 14720
rect 27903 14656 27919 14720
rect 27983 14656 27999 14720
rect 28063 14656 28079 14720
rect 28143 14656 28149 14720
rect 32206 14696 33006 14816
rect 27833 14655 28149 14656
rect 15469 14650 15535 14653
rect 19425 14650 19491 14653
rect 15469 14648 19491 14650
rect 15469 14592 15474 14648
rect 15530 14592 19430 14648
rect 19486 14592 19491 14648
rect 15469 14590 19491 14592
rect 15469 14587 15535 14590
rect 19425 14587 19491 14590
rect 19558 14588 19564 14652
rect 19628 14650 19634 14652
rect 19701 14650 19767 14653
rect 19628 14648 19767 14650
rect 19628 14592 19706 14648
rect 19762 14592 19767 14648
rect 19628 14590 19767 14592
rect 19628 14588 19634 14590
rect 19701 14587 19767 14590
rect 23841 14650 23907 14653
rect 24485 14650 24551 14653
rect 23841 14648 24551 14650
rect 23841 14592 23846 14648
rect 23902 14592 24490 14648
rect 24546 14592 24551 14648
rect 23841 14590 24551 14592
rect 23841 14587 23907 14590
rect 24485 14587 24551 14590
rect 25497 14650 25563 14653
rect 26325 14650 26391 14653
rect 25497 14648 26391 14650
rect 25497 14592 25502 14648
rect 25558 14592 26330 14648
rect 26386 14592 26391 14648
rect 25497 14590 26391 14592
rect 25497 14587 25563 14590
rect 26325 14587 26391 14590
rect 28625 14650 28691 14653
rect 29678 14650 29684 14652
rect 28625 14648 29684 14650
rect 28625 14592 28630 14648
rect 28686 14592 29684 14648
rect 28625 14590 29684 14592
rect 28625 14587 28691 14590
rect 29678 14588 29684 14590
rect 29748 14650 29754 14652
rect 30281 14650 30347 14653
rect 29748 14648 30347 14650
rect 29748 14592 30286 14648
rect 30342 14592 30347 14648
rect 29748 14590 30347 14592
rect 29748 14588 29754 14590
rect 30281 14587 30347 14590
rect 16757 14514 16823 14517
rect 11973 14512 14658 14514
rect 11973 14456 11978 14512
rect 12034 14456 14658 14512
rect 11973 14454 14658 14456
rect 14782 14512 16823 14514
rect 14782 14456 16762 14512
rect 16818 14456 16823 14512
rect 14782 14454 16823 14456
rect 11973 14451 12039 14454
rect 8628 14176 8944 14177
rect 8628 14112 8634 14176
rect 8698 14112 8714 14176
rect 8778 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8944 14176
rect 8628 14111 8944 14112
rect 12014 14044 12020 14108
rect 12084 14106 12090 14108
rect 14782 14106 14842 14454
rect 16757 14451 16823 14454
rect 17493 14514 17559 14517
rect 17861 14514 17927 14517
rect 17493 14512 17927 14514
rect 17493 14456 17498 14512
rect 17554 14456 17866 14512
rect 17922 14456 17927 14512
rect 17493 14454 17927 14456
rect 17493 14451 17559 14454
rect 17861 14451 17927 14454
rect 18413 14514 18479 14517
rect 20345 14514 20411 14517
rect 18413 14512 20411 14514
rect 18413 14456 18418 14512
rect 18474 14456 20350 14512
rect 20406 14456 20411 14512
rect 18413 14454 20411 14456
rect 18413 14451 18479 14454
rect 20345 14451 20411 14454
rect 25262 14452 25268 14516
rect 25332 14514 25338 14516
rect 26049 14514 26115 14517
rect 25332 14512 26115 14514
rect 25332 14456 26054 14512
rect 26110 14456 26115 14512
rect 25332 14454 26115 14456
rect 25332 14452 25338 14454
rect 26049 14451 26115 14454
rect 28073 14514 28139 14517
rect 28993 14514 29059 14517
rect 28073 14512 29059 14514
rect 28073 14456 28078 14512
rect 28134 14456 28998 14512
rect 29054 14456 29059 14512
rect 28073 14454 29059 14456
rect 28073 14451 28139 14454
rect 28993 14451 29059 14454
rect 15009 14378 15075 14381
rect 20529 14378 20595 14381
rect 15009 14376 16590 14378
rect 15009 14320 15014 14376
rect 15070 14344 16590 14376
rect 16806 14376 20595 14378
rect 16806 14344 20534 14376
rect 15070 14320 20534 14344
rect 20590 14320 20595 14376
rect 15009 14318 20595 14320
rect 15009 14315 15075 14318
rect 16530 14284 16866 14318
rect 20529 14315 20595 14318
rect 23054 14316 23060 14380
rect 23124 14378 23130 14380
rect 23473 14378 23539 14381
rect 28441 14378 28507 14381
rect 30373 14378 30439 14381
rect 32213 14378 32279 14381
rect 23124 14376 25514 14378
rect 23124 14320 23478 14376
rect 23534 14320 25514 14376
rect 23124 14318 25514 14320
rect 23124 14316 23130 14318
rect 23473 14315 23539 14318
rect 15142 14180 15148 14244
rect 15212 14242 15218 14244
rect 15929 14242 15995 14245
rect 15212 14240 15995 14242
rect 15212 14184 15934 14240
rect 15990 14184 15995 14240
rect 15212 14182 15995 14184
rect 15212 14180 15218 14182
rect 15929 14179 15995 14182
rect 16941 14242 17007 14245
rect 21582 14242 21588 14244
rect 16941 14240 21588 14242
rect 16941 14184 16946 14240
rect 17002 14184 21588 14240
rect 16941 14182 21588 14184
rect 16941 14179 17007 14182
rect 21582 14180 21588 14182
rect 21652 14180 21658 14244
rect 16310 14176 16626 14177
rect 16310 14112 16316 14176
rect 16380 14112 16396 14176
rect 16460 14112 16476 14176
rect 16540 14112 16556 14176
rect 16620 14112 16626 14176
rect 16310 14111 16626 14112
rect 23992 14176 24308 14177
rect 23992 14112 23998 14176
rect 24062 14112 24078 14176
rect 24142 14112 24158 14176
rect 24222 14112 24238 14176
rect 24302 14112 24308 14176
rect 23992 14111 24308 14112
rect 12084 14046 14842 14106
rect 12084 14044 12090 14046
rect 15510 14044 15516 14108
rect 15580 14106 15586 14108
rect 15837 14106 15903 14109
rect 15580 14104 15903 14106
rect 15580 14048 15842 14104
rect 15898 14048 15903 14104
rect 15580 14046 15903 14048
rect 15580 14044 15586 14046
rect 15837 14043 15903 14046
rect 16941 14106 17007 14109
rect 19609 14106 19675 14109
rect 16941 14104 19675 14106
rect 16941 14048 16946 14104
rect 17002 14048 19614 14104
rect 19670 14048 19675 14104
rect 16941 14046 19675 14048
rect 16941 14043 17007 14046
rect 19609 14043 19675 14046
rect 19885 14106 19951 14109
rect 24853 14106 24919 14109
rect 19885 14104 23904 14106
rect 19885 14048 19890 14104
rect 19946 14048 23904 14104
rect 19885 14046 23904 14048
rect 19885 14043 19951 14046
rect 14549 13970 14615 13973
rect 17493 13970 17559 13973
rect 18321 13970 18387 13973
rect 14549 13968 18387 13970
rect 14549 13912 14554 13968
rect 14610 13912 17498 13968
rect 17554 13912 18326 13968
rect 18382 13912 18387 13968
rect 14549 13910 18387 13912
rect 14549 13907 14615 13910
rect 17493 13907 17559 13910
rect 18321 13907 18387 13910
rect 18873 13970 18939 13973
rect 19006 13970 19012 13972
rect 18873 13968 19012 13970
rect 18873 13912 18878 13968
rect 18934 13912 19012 13968
rect 18873 13910 19012 13912
rect 18873 13907 18939 13910
rect 19006 13908 19012 13910
rect 19076 13908 19082 13972
rect 23844 13970 23904 14046
rect 24718 14104 24919 14106
rect 24718 14048 24858 14104
rect 24914 14048 24919 14104
rect 24718 14046 24919 14048
rect 25454 14106 25514 14318
rect 28441 14376 32279 14378
rect 28441 14320 28446 14376
rect 28502 14320 30378 14376
rect 30434 14320 32218 14376
rect 32274 14320 32279 14376
rect 28441 14318 32279 14320
rect 28441 14315 28507 14318
rect 30373 14315 30439 14318
rect 32213 14315 32279 14318
rect 26785 14242 26851 14245
rect 29361 14242 29427 14245
rect 26785 14240 29427 14242
rect 26785 14184 26790 14240
rect 26846 14184 29366 14240
rect 29422 14184 29427 14240
rect 26785 14182 29427 14184
rect 26785 14179 26851 14182
rect 29361 14179 29427 14182
rect 31674 14176 31990 14177
rect 31674 14112 31680 14176
rect 31744 14112 31760 14176
rect 31824 14112 31840 14176
rect 31904 14112 31920 14176
rect 31984 14112 31990 14176
rect 31674 14111 31990 14112
rect 29085 14106 29151 14109
rect 32206 14106 33006 14136
rect 25454 14104 29151 14106
rect 25454 14048 29090 14104
rect 29146 14048 29151 14104
rect 25454 14046 29151 14048
rect 24718 13970 24778 14046
rect 24853 14043 24919 14046
rect 29085 14043 29151 14046
rect 32078 14046 33006 14106
rect 23844 13910 24778 13970
rect 24853 13970 24919 13973
rect 25681 13970 25747 13973
rect 24853 13968 25747 13970
rect 24853 13912 24858 13968
rect 24914 13912 25686 13968
rect 25742 13912 25747 13968
rect 24853 13910 25747 13912
rect 24853 13907 24919 13910
rect 25681 13907 25747 13910
rect 25998 13908 26004 13972
rect 26068 13970 26074 13972
rect 26233 13970 26299 13973
rect 26068 13968 26299 13970
rect 26068 13912 26238 13968
rect 26294 13912 26299 13968
rect 26068 13910 26299 13912
rect 26068 13908 26074 13910
rect 26233 13907 26299 13910
rect 26601 13970 26667 13973
rect 29637 13970 29703 13973
rect 26601 13968 29703 13970
rect 26601 13912 26606 13968
rect 26662 13912 29642 13968
rect 29698 13912 29703 13968
rect 26601 13910 29703 13912
rect 26601 13907 26667 13910
rect 29637 13907 29703 13910
rect 30005 13970 30071 13973
rect 32078 13970 32138 14046
rect 32206 14016 33006 14046
rect 30005 13968 32138 13970
rect 30005 13912 30010 13968
rect 30066 13912 32138 13968
rect 30005 13910 32138 13912
rect 30005 13907 30071 13910
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 14733 13834 14799 13837
rect 17217 13834 17283 13837
rect 20846 13834 20852 13836
rect 14733 13832 20852 13834
rect 14733 13776 14738 13832
rect 14794 13776 17222 13832
rect 17278 13776 20852 13832
rect 14733 13774 20852 13776
rect 14733 13771 14799 13774
rect 17217 13771 17283 13774
rect 20846 13772 20852 13774
rect 20916 13772 20922 13836
rect 22461 13834 22527 13837
rect 24025 13834 24091 13837
rect 22461 13832 24091 13834
rect 22461 13776 22466 13832
rect 22522 13776 24030 13832
rect 24086 13776 24091 13832
rect 22461 13774 24091 13776
rect 22461 13771 22527 13774
rect 24025 13771 24091 13774
rect 24761 13834 24827 13837
rect 25262 13834 25268 13836
rect 24761 13832 25268 13834
rect 24761 13776 24766 13832
rect 24822 13776 25268 13832
rect 24761 13774 25268 13776
rect 24761 13771 24827 13774
rect 25262 13772 25268 13774
rect 25332 13772 25338 13836
rect 25814 13772 25820 13836
rect 25884 13834 25890 13836
rect 25957 13834 26023 13837
rect 25884 13832 26023 13834
rect 25884 13776 25962 13832
rect 26018 13776 26023 13832
rect 25884 13774 26023 13776
rect 25884 13772 25890 13774
rect 25957 13771 26023 13774
rect 26550 13772 26556 13836
rect 26620 13834 26626 13836
rect 26877 13834 26943 13837
rect 28165 13836 28231 13837
rect 28165 13834 28212 13836
rect 26620 13832 26943 13834
rect 26620 13776 26882 13832
rect 26938 13776 26943 13832
rect 26620 13774 26943 13776
rect 28120 13832 28212 13834
rect 28120 13776 28170 13832
rect 28120 13774 28212 13776
rect 26620 13772 26626 13774
rect 26877 13771 26943 13774
rect 28165 13772 28212 13774
rect 28276 13772 28282 13836
rect 29729 13834 29795 13837
rect 29862 13834 29868 13836
rect 29729 13832 29868 13834
rect 29729 13776 29734 13832
rect 29790 13776 29868 13832
rect 29729 13774 29868 13776
rect 28165 13771 28231 13772
rect 29729 13771 29795 13774
rect 29862 13772 29868 13774
rect 29932 13772 29938 13836
rect 13445 13698 13511 13701
rect 19977 13698 20043 13701
rect 13445 13696 20043 13698
rect 13445 13640 13450 13696
rect 13506 13640 19982 13696
rect 20038 13640 20043 13696
rect 13445 13638 20043 13640
rect 13445 13635 13511 13638
rect 19977 13635 20043 13638
rect 21541 13698 21607 13701
rect 23565 13698 23631 13701
rect 21541 13696 23631 13698
rect 21541 13640 21546 13696
rect 21602 13640 23570 13696
rect 23626 13640 23631 13696
rect 21541 13638 23631 13640
rect 21541 13635 21607 13638
rect 23565 13635 23631 13638
rect 4787 13632 5103 13633
rect 4787 13568 4793 13632
rect 4857 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5103 13632
rect 4787 13567 5103 13568
rect 12469 13632 12785 13633
rect 12469 13568 12475 13632
rect 12539 13568 12555 13632
rect 12619 13568 12635 13632
rect 12699 13568 12715 13632
rect 12779 13568 12785 13632
rect 12469 13567 12785 13568
rect 20151 13632 20467 13633
rect 20151 13568 20157 13632
rect 20221 13568 20237 13632
rect 20301 13568 20317 13632
rect 20381 13568 20397 13632
rect 20461 13568 20467 13632
rect 20151 13567 20467 13568
rect 27833 13632 28149 13633
rect 27833 13568 27839 13632
rect 27903 13568 27919 13632
rect 27983 13568 27999 13632
rect 28063 13568 28079 13632
rect 28143 13568 28149 13632
rect 27833 13567 28149 13568
rect 19149 13562 19215 13565
rect 19149 13560 19580 13562
rect 19149 13504 19154 13560
rect 19210 13504 19580 13560
rect 19149 13502 19580 13504
rect 19149 13499 19215 13502
rect 6862 13364 6868 13428
rect 6932 13426 6938 13428
rect 19333 13426 19399 13429
rect 6932 13424 19399 13426
rect 6932 13368 19338 13424
rect 19394 13368 19399 13424
rect 6932 13366 19399 13368
rect 19520 13426 19580 13502
rect 21030 13500 21036 13564
rect 21100 13562 21106 13564
rect 25405 13562 25471 13565
rect 21100 13560 25471 13562
rect 21100 13504 25410 13560
rect 25466 13504 25471 13560
rect 21100 13502 25471 13504
rect 21100 13500 21106 13502
rect 25405 13499 25471 13502
rect 31109 13564 31175 13565
rect 31109 13560 31156 13564
rect 31220 13562 31226 13564
rect 31109 13504 31114 13560
rect 31109 13500 31156 13504
rect 31220 13502 31266 13562
rect 31220 13500 31226 13502
rect 31109 13499 31175 13500
rect 22093 13426 22159 13429
rect 24577 13426 24643 13429
rect 19520 13366 22018 13426
rect 6932 13364 6938 13366
rect 19333 13363 19399 13366
rect 16297 13290 16363 13293
rect 18505 13290 18571 13293
rect 19057 13290 19123 13293
rect 20805 13290 20871 13293
rect 21725 13290 21791 13293
rect 16297 13288 21791 13290
rect 16297 13232 16302 13288
rect 16358 13232 18510 13288
rect 18566 13232 19062 13288
rect 19118 13232 20810 13288
rect 20866 13232 21730 13288
rect 21786 13232 21791 13288
rect 16297 13230 21791 13232
rect 21958 13290 22018 13366
rect 22093 13424 24643 13426
rect 22093 13368 22098 13424
rect 22154 13368 24582 13424
rect 24638 13368 24643 13424
rect 22093 13366 24643 13368
rect 22093 13363 22159 13366
rect 24577 13363 24643 13366
rect 26325 13426 26391 13429
rect 29177 13426 29243 13429
rect 26325 13424 29243 13426
rect 26325 13368 26330 13424
rect 26386 13368 29182 13424
rect 29238 13368 29243 13424
rect 26325 13366 29243 13368
rect 26325 13363 26391 13366
rect 29177 13363 29243 13366
rect 31385 13426 31451 13429
rect 32206 13426 33006 13456
rect 31385 13424 33006 13426
rect 31385 13368 31390 13424
rect 31446 13368 33006 13424
rect 31385 13366 33006 13368
rect 31385 13363 31451 13366
rect 32206 13336 33006 13366
rect 22369 13290 22435 13293
rect 21958 13288 22435 13290
rect 21958 13232 22374 13288
rect 22430 13232 22435 13288
rect 21958 13230 22435 13232
rect 16297 13227 16363 13230
rect 18505 13227 18571 13230
rect 19057 13227 19123 13230
rect 20805 13227 20871 13230
rect 21725 13227 21791 13230
rect 22369 13227 22435 13230
rect 25681 13290 25747 13293
rect 28717 13290 28783 13293
rect 25681 13288 28783 13290
rect 25681 13232 25686 13288
rect 25742 13232 28722 13288
rect 28778 13232 28783 13288
rect 25681 13230 28783 13232
rect 25681 13227 25747 13230
rect 28717 13227 28783 13230
rect 16757 13154 16823 13157
rect 17953 13154 18019 13157
rect 16757 13152 18019 13154
rect 16757 13096 16762 13152
rect 16818 13096 17958 13152
rect 18014 13096 18019 13152
rect 16757 13094 18019 13096
rect 16757 13091 16823 13094
rect 17953 13091 18019 13094
rect 18781 13154 18847 13157
rect 19793 13154 19859 13157
rect 18781 13152 19859 13154
rect 18781 13096 18786 13152
rect 18842 13096 19798 13152
rect 19854 13096 19859 13152
rect 18781 13094 19859 13096
rect 18781 13091 18847 13094
rect 19793 13091 19859 13094
rect 20529 13154 20595 13157
rect 21357 13154 21423 13157
rect 20529 13152 21423 13154
rect 20529 13096 20534 13152
rect 20590 13096 21362 13152
rect 21418 13096 21423 13152
rect 20529 13094 21423 13096
rect 20529 13091 20595 13094
rect 21357 13091 21423 13094
rect 21950 13092 21956 13156
rect 22020 13154 22026 13156
rect 23841 13154 23907 13157
rect 25497 13156 25563 13157
rect 25446 13154 25452 13156
rect 22020 13152 23907 13154
rect 22020 13096 23846 13152
rect 23902 13096 23907 13152
rect 22020 13094 23907 13096
rect 25406 13094 25452 13154
rect 25516 13152 25563 13156
rect 25558 13096 25563 13152
rect 22020 13092 22026 13094
rect 23841 13091 23907 13094
rect 25446 13092 25452 13094
rect 25516 13092 25563 13096
rect 27654 13092 27660 13156
rect 27724 13154 27730 13156
rect 28901 13154 28967 13157
rect 27724 13152 28967 13154
rect 27724 13096 28906 13152
rect 28962 13096 28967 13152
rect 27724 13094 28967 13096
rect 27724 13092 27730 13094
rect 25497 13091 25563 13092
rect 28901 13091 28967 13094
rect 8628 13088 8944 13089
rect 0 13018 800 13048
rect 8628 13024 8634 13088
rect 8698 13024 8714 13088
rect 8778 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8944 13088
rect 8628 13023 8944 13024
rect 16310 13088 16626 13089
rect 16310 13024 16316 13088
rect 16380 13024 16396 13088
rect 16460 13024 16476 13088
rect 16540 13024 16556 13088
rect 16620 13024 16626 13088
rect 16310 13023 16626 13024
rect 23992 13088 24308 13089
rect 23992 13024 23998 13088
rect 24062 13024 24078 13088
rect 24142 13024 24158 13088
rect 24222 13024 24238 13088
rect 24302 13024 24308 13088
rect 23992 13023 24308 13024
rect 31674 13088 31990 13089
rect 31674 13024 31680 13088
rect 31744 13024 31760 13088
rect 31824 13024 31840 13088
rect 31904 13024 31920 13088
rect 31984 13024 31990 13088
rect 31674 13023 31990 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 800 12958
rect 1577 12955 1643 12958
rect 16849 13018 16915 13021
rect 25037 13018 25103 13021
rect 26366 13018 26372 13020
rect 16849 13016 23858 13018
rect 16849 12960 16854 13016
rect 16910 12960 23858 13016
rect 16849 12958 23858 12960
rect 16849 12955 16915 12958
rect 12893 12882 12959 12885
rect 21541 12882 21607 12885
rect 23798 12884 23858 12958
rect 25037 13016 26372 13018
rect 25037 12960 25042 13016
rect 25098 12960 26372 13016
rect 25037 12958 26372 12960
rect 25037 12955 25103 12958
rect 26366 12956 26372 12958
rect 26436 12956 26442 13020
rect 27337 13018 27403 13021
rect 29494 13018 29500 13020
rect 27337 13016 29500 13018
rect 27337 12960 27342 13016
rect 27398 12960 29500 13016
rect 27337 12958 29500 12960
rect 27337 12955 27403 12958
rect 29494 12956 29500 12958
rect 29564 12956 29570 13020
rect 12893 12880 21607 12882
rect 12893 12824 12898 12880
rect 12954 12824 21546 12880
rect 21602 12824 21607 12880
rect 12893 12822 21607 12824
rect 12893 12819 12959 12822
rect 21541 12819 21607 12822
rect 23790 12820 23796 12884
rect 23860 12882 23866 12884
rect 24209 12882 24275 12885
rect 23860 12880 24275 12882
rect 23860 12824 24214 12880
rect 24270 12824 24275 12880
rect 23860 12822 24275 12824
rect 23860 12820 23866 12822
rect 24209 12819 24275 12822
rect 27286 12820 27292 12884
rect 27356 12882 27362 12884
rect 27705 12882 27771 12885
rect 27356 12880 27771 12882
rect 27356 12824 27710 12880
rect 27766 12824 27771 12880
rect 27356 12822 27771 12824
rect 27356 12820 27362 12822
rect 27705 12819 27771 12822
rect 28390 12820 28396 12884
rect 28460 12882 28466 12884
rect 28533 12882 28599 12885
rect 28460 12880 28599 12882
rect 28460 12824 28538 12880
rect 28594 12824 28599 12880
rect 28460 12822 28599 12824
rect 28460 12820 28466 12822
rect 28533 12819 28599 12822
rect 4061 12746 4127 12749
rect 25405 12746 25471 12749
rect 28942 12746 28948 12748
rect 4061 12744 25471 12746
rect 4061 12688 4066 12744
rect 4122 12688 25410 12744
rect 25466 12688 25471 12744
rect 4061 12686 25471 12688
rect 4061 12683 4127 12686
rect 25405 12683 25471 12686
rect 25592 12686 28948 12746
rect 15653 12610 15719 12613
rect 19885 12610 19951 12613
rect 15653 12608 19951 12610
rect 15653 12552 15658 12608
rect 15714 12552 19890 12608
rect 19946 12552 19951 12608
rect 15653 12550 19951 12552
rect 15653 12547 15719 12550
rect 19885 12547 19951 12550
rect 21398 12548 21404 12612
rect 21468 12610 21474 12612
rect 21541 12610 21607 12613
rect 21468 12608 21607 12610
rect 21468 12552 21546 12608
rect 21602 12552 21607 12608
rect 21468 12550 21607 12552
rect 21468 12548 21474 12550
rect 21541 12547 21607 12550
rect 21725 12610 21791 12613
rect 25592 12610 25652 12686
rect 28942 12684 28948 12686
rect 29012 12684 29018 12748
rect 32206 12656 33006 12776
rect 21725 12608 25652 12610
rect 21725 12552 21730 12608
rect 21786 12552 25652 12608
rect 21725 12550 25652 12552
rect 21725 12547 21791 12550
rect 4787 12544 5103 12545
rect 4787 12480 4793 12544
rect 4857 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5103 12544
rect 4787 12479 5103 12480
rect 12469 12544 12785 12545
rect 12469 12480 12475 12544
rect 12539 12480 12555 12544
rect 12619 12480 12635 12544
rect 12699 12480 12715 12544
rect 12779 12480 12785 12544
rect 12469 12479 12785 12480
rect 20151 12544 20467 12545
rect 20151 12480 20157 12544
rect 20221 12480 20237 12544
rect 20301 12480 20317 12544
rect 20381 12480 20397 12544
rect 20461 12480 20467 12544
rect 20151 12479 20467 12480
rect 27833 12544 28149 12545
rect 27833 12480 27839 12544
rect 27903 12480 27919 12544
rect 27983 12480 27999 12544
rect 28063 12480 28079 12544
rect 28143 12480 28149 12544
rect 27833 12479 28149 12480
rect 16021 12474 16087 12477
rect 18873 12474 18939 12477
rect 16021 12472 18939 12474
rect 16021 12416 16026 12472
rect 16082 12416 18878 12472
rect 18934 12416 18939 12472
rect 16021 12414 18939 12416
rect 16021 12411 16087 12414
rect 18873 12411 18939 12414
rect 21449 12474 21515 12477
rect 23841 12474 23907 12477
rect 27613 12474 27679 12477
rect 21449 12472 23907 12474
rect 21449 12416 21454 12472
rect 21510 12416 23846 12472
rect 23902 12416 23907 12472
rect 21449 12414 23907 12416
rect 21449 12411 21515 12414
rect 23841 12411 23907 12414
rect 24948 12472 27679 12474
rect 24948 12416 27618 12472
rect 27674 12416 27679 12472
rect 24948 12414 27679 12416
rect 10685 12338 10751 12341
rect 17902 12338 17908 12340
rect 10685 12336 17908 12338
rect 10685 12280 10690 12336
rect 10746 12280 17908 12336
rect 10685 12278 17908 12280
rect 10685 12275 10751 12278
rect 17902 12276 17908 12278
rect 17972 12276 17978 12340
rect 24948 12338 25008 12414
rect 27613 12411 27679 12414
rect 20670 12278 25008 12338
rect 0 12112 800 12232
rect 18822 12140 18828 12204
rect 18892 12202 18898 12204
rect 20670 12202 20730 12278
rect 25078 12276 25084 12340
rect 25148 12338 25154 12340
rect 25865 12338 25931 12341
rect 25148 12336 25931 12338
rect 25148 12280 25870 12336
rect 25926 12280 25931 12336
rect 25148 12278 25931 12280
rect 25148 12276 25154 12278
rect 25865 12275 25931 12278
rect 24894 12202 24900 12204
rect 18892 12142 20730 12202
rect 23430 12142 24900 12202
rect 18892 12140 18898 12142
rect 19517 12068 19583 12069
rect 19517 12066 19564 12068
rect 19472 12064 19564 12066
rect 19472 12008 19522 12064
rect 19472 12006 19564 12008
rect 19517 12004 19564 12006
rect 19628 12004 19634 12068
rect 19977 12066 20043 12069
rect 23430 12066 23490 12142
rect 24894 12140 24900 12142
rect 24964 12140 24970 12204
rect 25129 12202 25195 12205
rect 31569 12202 31635 12205
rect 25129 12200 31635 12202
rect 25129 12144 25134 12200
rect 25190 12144 31574 12200
rect 31630 12144 31635 12200
rect 25129 12142 31635 12144
rect 25129 12139 25195 12142
rect 31569 12139 31635 12142
rect 32206 12066 33006 12096
rect 19977 12064 23490 12066
rect 19977 12008 19982 12064
rect 20038 12008 23490 12064
rect 19977 12006 23490 12008
rect 32078 12006 33006 12066
rect 19517 12003 19583 12004
rect 19977 12003 20043 12006
rect 8628 12000 8944 12001
rect 8628 11936 8634 12000
rect 8698 11936 8714 12000
rect 8778 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8944 12000
rect 8628 11935 8944 11936
rect 16310 12000 16626 12001
rect 16310 11936 16316 12000
rect 16380 11936 16396 12000
rect 16460 11936 16476 12000
rect 16540 11936 16556 12000
rect 16620 11936 16626 12000
rect 16310 11935 16626 11936
rect 23992 12000 24308 12001
rect 23992 11936 23998 12000
rect 24062 11936 24078 12000
rect 24142 11936 24158 12000
rect 24222 11936 24238 12000
rect 24302 11936 24308 12000
rect 23992 11935 24308 11936
rect 31674 12000 31990 12001
rect 31674 11936 31680 12000
rect 31744 11936 31760 12000
rect 31824 11936 31840 12000
rect 31904 11936 31920 12000
rect 31984 11936 31990 12000
rect 31674 11935 31990 11936
rect 17769 11930 17835 11933
rect 23565 11930 23631 11933
rect 17769 11928 23631 11930
rect 17769 11872 17774 11928
rect 17830 11872 23570 11928
rect 23626 11872 23631 11928
rect 17769 11870 23631 11872
rect 17769 11867 17835 11870
rect 23565 11867 23631 11870
rect 24710 11868 24716 11932
rect 24780 11930 24786 11932
rect 26141 11930 26207 11933
rect 26969 11932 27035 11933
rect 26918 11930 26924 11932
rect 24780 11928 26207 11930
rect 24780 11872 26146 11928
rect 26202 11872 26207 11928
rect 24780 11870 26207 11872
rect 26878 11870 26924 11930
rect 26988 11928 27035 11932
rect 27030 11872 27035 11928
rect 24780 11868 24786 11870
rect 26141 11867 26207 11870
rect 26918 11868 26924 11870
rect 26988 11868 27035 11872
rect 26969 11867 27035 11868
rect 10317 11794 10383 11797
rect 20662 11794 20668 11796
rect 10317 11792 20668 11794
rect 10317 11736 10322 11792
rect 10378 11736 20668 11792
rect 10317 11734 20668 11736
rect 10317 11731 10383 11734
rect 20662 11732 20668 11734
rect 20732 11732 20738 11796
rect 31293 11794 31359 11797
rect 32078 11794 32138 12006
rect 32206 11976 33006 12006
rect 31293 11792 32138 11794
rect 31293 11736 31298 11792
rect 31354 11736 32138 11792
rect 31293 11734 32138 11736
rect 31293 11731 31359 11734
rect 13169 11658 13235 11661
rect 21449 11658 21515 11661
rect 13169 11656 21515 11658
rect 13169 11600 13174 11656
rect 13230 11600 21454 11656
rect 21510 11600 21515 11656
rect 13169 11598 21515 11600
rect 13169 11595 13235 11598
rect 21449 11595 21515 11598
rect 12985 11522 13051 11525
rect 19977 11522 20043 11525
rect 12985 11520 20043 11522
rect 12985 11464 12990 11520
rect 13046 11464 19982 11520
rect 20038 11464 20043 11520
rect 12985 11462 20043 11464
rect 12985 11459 13051 11462
rect 19977 11459 20043 11462
rect 4787 11456 5103 11457
rect 0 11386 800 11416
rect 4787 11392 4793 11456
rect 4857 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5103 11456
rect 4787 11391 5103 11392
rect 12469 11456 12785 11457
rect 12469 11392 12475 11456
rect 12539 11392 12555 11456
rect 12619 11392 12635 11456
rect 12699 11392 12715 11456
rect 12779 11392 12785 11456
rect 12469 11391 12785 11392
rect 20151 11456 20467 11457
rect 20151 11392 20157 11456
rect 20221 11392 20237 11456
rect 20301 11392 20317 11456
rect 20381 11392 20397 11456
rect 20461 11392 20467 11456
rect 20151 11391 20467 11392
rect 27833 11456 28149 11457
rect 27833 11392 27839 11456
rect 27903 11392 27919 11456
rect 27983 11392 27999 11456
rect 28063 11392 28079 11456
rect 28143 11392 28149 11456
rect 27833 11391 28149 11392
rect 1577 11386 1643 11389
rect 0 11384 1643 11386
rect 0 11328 1582 11384
rect 1638 11328 1643 11384
rect 0 11326 1643 11328
rect 0 11296 800 11326
rect 1577 11323 1643 11326
rect 26182 11324 26188 11388
rect 26252 11386 26258 11388
rect 26601 11386 26667 11389
rect 26252 11384 26667 11386
rect 26252 11328 26606 11384
rect 26662 11328 26667 11384
rect 26252 11326 26667 11328
rect 26252 11324 26258 11326
rect 26601 11323 26667 11326
rect 31293 11386 31359 11389
rect 32206 11386 33006 11416
rect 31293 11384 33006 11386
rect 31293 11328 31298 11384
rect 31354 11328 33006 11384
rect 31293 11326 33006 11328
rect 31293 11323 31359 11326
rect 32206 11296 33006 11326
rect 7281 11250 7347 11253
rect 28809 11250 28875 11253
rect 7281 11248 28875 11250
rect 7281 11192 7286 11248
rect 7342 11192 28814 11248
rect 28870 11192 28875 11248
rect 7281 11190 28875 11192
rect 7281 11187 7347 11190
rect 28809 11187 28875 11190
rect 7373 11114 7439 11117
rect 28533 11116 28599 11117
rect 28533 11114 28580 11116
rect 7373 11112 28580 11114
rect 28644 11114 28650 11116
rect 7373 11056 7378 11112
rect 7434 11056 28538 11112
rect 7373 11054 28580 11056
rect 7373 11051 7439 11054
rect 28533 11052 28580 11054
rect 28644 11054 28726 11114
rect 28644 11052 28650 11054
rect 28533 11051 28599 11052
rect 27102 10916 27108 10980
rect 27172 10978 27178 10980
rect 27613 10978 27679 10981
rect 31385 10980 31451 10981
rect 27172 10976 27679 10978
rect 27172 10920 27618 10976
rect 27674 10920 27679 10976
rect 27172 10918 27679 10920
rect 27172 10916 27178 10918
rect 27613 10915 27679 10918
rect 31334 10916 31340 10980
rect 31404 10978 31451 10980
rect 31404 10976 31496 10978
rect 31446 10920 31496 10976
rect 31404 10918 31496 10920
rect 31404 10916 31451 10918
rect 31385 10915 31451 10916
rect 8628 10912 8944 10913
rect 8628 10848 8634 10912
rect 8698 10848 8714 10912
rect 8778 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8944 10912
rect 8628 10847 8944 10848
rect 16310 10912 16626 10913
rect 16310 10848 16316 10912
rect 16380 10848 16396 10912
rect 16460 10848 16476 10912
rect 16540 10848 16556 10912
rect 16620 10848 16626 10912
rect 16310 10847 16626 10848
rect 23992 10912 24308 10913
rect 23992 10848 23998 10912
rect 24062 10848 24078 10912
rect 24142 10848 24158 10912
rect 24222 10848 24238 10912
rect 24302 10848 24308 10912
rect 23992 10847 24308 10848
rect 31674 10912 31990 10913
rect 31674 10848 31680 10912
rect 31744 10848 31760 10912
rect 31824 10848 31840 10912
rect 31904 10848 31920 10912
rect 31984 10848 31990 10912
rect 31674 10847 31990 10848
rect 20897 10842 20963 10845
rect 22277 10842 22343 10845
rect 20897 10840 22343 10842
rect 20897 10784 20902 10840
rect 20958 10784 22282 10840
rect 22338 10784 22343 10840
rect 20897 10782 22343 10784
rect 20897 10779 20963 10782
rect 22277 10779 22343 10782
rect 29637 10842 29703 10845
rect 30414 10842 30420 10844
rect 29637 10840 30420 10842
rect 29637 10784 29642 10840
rect 29698 10784 30420 10840
rect 29637 10782 30420 10784
rect 29637 10779 29703 10782
rect 30414 10780 30420 10782
rect 30484 10842 30490 10844
rect 31017 10842 31083 10845
rect 30484 10840 31083 10842
rect 30484 10784 31022 10840
rect 31078 10784 31083 10840
rect 30484 10782 31083 10784
rect 30484 10780 30490 10782
rect 31017 10779 31083 10782
rect 20897 10708 20963 10709
rect 20846 10644 20852 10708
rect 20916 10706 20963 10708
rect 20916 10704 21008 10706
rect 20958 10648 21008 10704
rect 20916 10646 21008 10648
rect 20916 10644 20963 10646
rect 23606 10644 23612 10708
rect 23676 10706 23682 10708
rect 24301 10706 24367 10709
rect 23676 10704 24367 10706
rect 23676 10648 24306 10704
rect 24362 10648 24367 10704
rect 23676 10646 24367 10648
rect 23676 10644 23682 10646
rect 20897 10643 20963 10644
rect 24301 10643 24367 10646
rect 32206 10616 33006 10736
rect 0 10570 800 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 800 10510
rect 1577 10507 1643 10510
rect 10542 10508 10548 10572
rect 10612 10570 10618 10572
rect 29913 10570 29979 10573
rect 10612 10568 29979 10570
rect 10612 10512 29918 10568
rect 29974 10512 29979 10568
rect 10612 10510 29979 10512
rect 10612 10508 10618 10510
rect 29913 10507 29979 10510
rect 15745 10434 15811 10437
rect 19701 10434 19767 10437
rect 15745 10432 19767 10434
rect 15745 10376 15750 10432
rect 15806 10376 19706 10432
rect 19762 10376 19767 10432
rect 15745 10374 19767 10376
rect 15745 10371 15811 10374
rect 19701 10371 19767 10374
rect 22185 10434 22251 10437
rect 23197 10434 23263 10437
rect 22185 10432 23263 10434
rect 22185 10376 22190 10432
rect 22246 10376 23202 10432
rect 23258 10376 23263 10432
rect 22185 10374 23263 10376
rect 22185 10371 22251 10374
rect 23197 10371 23263 10374
rect 23841 10434 23907 10437
rect 26601 10434 26667 10437
rect 23841 10432 26667 10434
rect 23841 10376 23846 10432
rect 23902 10376 26606 10432
rect 26662 10376 26667 10432
rect 23841 10374 26667 10376
rect 23841 10371 23907 10374
rect 26601 10371 26667 10374
rect 4787 10368 5103 10369
rect 4787 10304 4793 10368
rect 4857 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5103 10368
rect 4787 10303 5103 10304
rect 12469 10368 12785 10369
rect 12469 10304 12475 10368
rect 12539 10304 12555 10368
rect 12619 10304 12635 10368
rect 12699 10304 12715 10368
rect 12779 10304 12785 10368
rect 12469 10303 12785 10304
rect 20151 10368 20467 10369
rect 20151 10304 20157 10368
rect 20221 10304 20237 10368
rect 20301 10304 20317 10368
rect 20381 10304 20397 10368
rect 20461 10304 20467 10368
rect 20151 10303 20467 10304
rect 27833 10368 28149 10369
rect 27833 10304 27839 10368
rect 27903 10304 27919 10368
rect 27983 10304 27999 10368
rect 28063 10304 28079 10368
rect 28143 10304 28149 10368
rect 27833 10303 28149 10304
rect 20897 10298 20963 10301
rect 25129 10298 25195 10301
rect 20897 10296 25195 10298
rect 20897 10240 20902 10296
rect 20958 10240 25134 10296
rect 25190 10240 25195 10296
rect 20897 10238 25195 10240
rect 20897 10235 20963 10238
rect 25129 10235 25195 10238
rect 6494 10100 6500 10164
rect 6564 10162 6570 10164
rect 30925 10162 30991 10165
rect 6564 10160 30991 10162
rect 6564 10104 30930 10160
rect 30986 10104 30991 10160
rect 6564 10102 30991 10104
rect 6564 10100 6570 10102
rect 30925 10099 30991 10102
rect 15878 9964 15884 10028
rect 15948 10026 15954 10028
rect 29729 10026 29795 10029
rect 15948 10024 29795 10026
rect 15948 9968 29734 10024
rect 29790 9968 29795 10024
rect 15948 9966 29795 9968
rect 15948 9964 15954 9966
rect 29729 9963 29795 9966
rect 31293 10026 31359 10029
rect 32206 10026 33006 10056
rect 31293 10024 33006 10026
rect 31293 9968 31298 10024
rect 31354 9968 33006 10024
rect 31293 9966 33006 9968
rect 31293 9963 31359 9966
rect 32206 9936 33006 9966
rect 8628 9824 8944 9825
rect 0 9664 800 9784
rect 8628 9760 8634 9824
rect 8698 9760 8714 9824
rect 8778 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8944 9824
rect 8628 9759 8944 9760
rect 16310 9824 16626 9825
rect 16310 9760 16316 9824
rect 16380 9760 16396 9824
rect 16460 9760 16476 9824
rect 16540 9760 16556 9824
rect 16620 9760 16626 9824
rect 16310 9759 16626 9760
rect 23992 9824 24308 9825
rect 23992 9760 23998 9824
rect 24062 9760 24078 9824
rect 24142 9760 24158 9824
rect 24222 9760 24238 9824
rect 24302 9760 24308 9824
rect 23992 9759 24308 9760
rect 31674 9824 31990 9825
rect 31674 9760 31680 9824
rect 31744 9760 31760 9824
rect 31824 9760 31840 9824
rect 31904 9760 31920 9824
rect 31984 9760 31990 9824
rect 31674 9759 31990 9760
rect 26417 9754 26483 9757
rect 27102 9754 27108 9756
rect 26374 9752 27108 9754
rect 26374 9696 26422 9752
rect 26478 9696 27108 9752
rect 26374 9694 27108 9696
rect 26374 9691 26483 9694
rect 27102 9692 27108 9694
rect 27172 9692 27178 9756
rect 5441 9620 5507 9621
rect 5390 9618 5396 9620
rect 5350 9558 5396 9618
rect 5460 9616 5507 9620
rect 5502 9560 5507 9616
rect 5390 9556 5396 9558
rect 5460 9556 5507 9560
rect 5441 9555 5507 9556
rect 6545 9618 6611 9621
rect 25405 9618 25471 9621
rect 25814 9618 25820 9620
rect 6545 9616 25330 9618
rect 6545 9560 6550 9616
rect 6606 9560 25330 9616
rect 6545 9558 25330 9560
rect 6545 9555 6611 9558
rect 8385 9482 8451 9485
rect 25037 9482 25103 9485
rect 8385 9480 25103 9482
rect 8385 9424 8390 9480
rect 8446 9424 25042 9480
rect 25098 9424 25103 9480
rect 8385 9422 25103 9424
rect 25270 9482 25330 9558
rect 25405 9616 25820 9618
rect 25405 9560 25410 9616
rect 25466 9560 25820 9616
rect 25405 9558 25820 9560
rect 25405 9555 25471 9558
rect 25814 9556 25820 9558
rect 25884 9556 25890 9620
rect 26374 9482 26434 9691
rect 25270 9422 26434 9482
rect 8385 9419 8451 9422
rect 25037 9419 25103 9422
rect 26417 9346 26483 9349
rect 26734 9346 26740 9348
rect 26417 9344 26740 9346
rect 26417 9288 26422 9344
rect 26478 9288 26740 9344
rect 26417 9286 26740 9288
rect 26417 9283 26483 9286
rect 26734 9284 26740 9286
rect 26804 9284 26810 9348
rect 31293 9346 31359 9349
rect 32206 9346 33006 9376
rect 31293 9344 33006 9346
rect 31293 9288 31298 9344
rect 31354 9288 33006 9344
rect 31293 9286 33006 9288
rect 31293 9283 31359 9286
rect 4787 9280 5103 9281
rect 4787 9216 4793 9280
rect 4857 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5103 9280
rect 4787 9215 5103 9216
rect 12469 9280 12785 9281
rect 12469 9216 12475 9280
rect 12539 9216 12555 9280
rect 12619 9216 12635 9280
rect 12699 9216 12715 9280
rect 12779 9216 12785 9280
rect 12469 9215 12785 9216
rect 20151 9280 20467 9281
rect 20151 9216 20157 9280
rect 20221 9216 20237 9280
rect 20301 9216 20317 9280
rect 20381 9216 20397 9280
rect 20461 9216 20467 9280
rect 20151 9215 20467 9216
rect 27833 9280 28149 9281
rect 27833 9216 27839 9280
rect 27903 9216 27919 9280
rect 27983 9216 27999 9280
rect 28063 9216 28079 9280
rect 28143 9216 28149 9280
rect 32206 9256 33006 9286
rect 27833 9215 28149 9216
rect 13302 9012 13308 9076
rect 13372 9074 13378 9076
rect 25405 9074 25471 9077
rect 13372 9072 25471 9074
rect 13372 9016 25410 9072
rect 25466 9016 25471 9072
rect 13372 9014 25471 9016
rect 13372 9012 13378 9014
rect 25405 9011 25471 9014
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 15326 8876 15332 8940
rect 15396 8938 15402 8940
rect 25221 8938 25287 8941
rect 15396 8936 25287 8938
rect 15396 8880 25226 8936
rect 25282 8880 25287 8936
rect 15396 8878 25287 8880
rect 15396 8876 15402 8878
rect 25221 8875 25287 8878
rect 28942 8740 28948 8804
rect 29012 8802 29018 8804
rect 29085 8802 29151 8805
rect 29012 8800 29151 8802
rect 29012 8744 29090 8800
rect 29146 8744 29151 8800
rect 29012 8742 29151 8744
rect 29012 8740 29018 8742
rect 29085 8739 29151 8742
rect 8628 8736 8944 8737
rect 8628 8672 8634 8736
rect 8698 8672 8714 8736
rect 8778 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8944 8736
rect 8628 8671 8944 8672
rect 16310 8736 16626 8737
rect 16310 8672 16316 8736
rect 16380 8672 16396 8736
rect 16460 8672 16476 8736
rect 16540 8672 16556 8736
rect 16620 8672 16626 8736
rect 16310 8671 16626 8672
rect 23992 8736 24308 8737
rect 23992 8672 23998 8736
rect 24062 8672 24078 8736
rect 24142 8672 24158 8736
rect 24222 8672 24238 8736
rect 24302 8672 24308 8736
rect 23992 8671 24308 8672
rect 31674 8736 31990 8737
rect 31674 8672 31680 8736
rect 31744 8672 31760 8736
rect 31824 8672 31840 8736
rect 31904 8672 31920 8736
rect 31984 8672 31990 8736
rect 31674 8671 31990 8672
rect 17718 8604 17724 8668
rect 17788 8666 17794 8668
rect 19517 8666 19583 8669
rect 29729 8668 29795 8669
rect 17788 8664 19583 8666
rect 17788 8608 19522 8664
rect 19578 8608 19583 8664
rect 17788 8606 19583 8608
rect 17788 8604 17794 8606
rect 19517 8603 19583 8606
rect 29678 8604 29684 8668
rect 29748 8666 29795 8668
rect 30046 8666 30052 8668
rect 29748 8664 30052 8666
rect 29790 8608 30052 8664
rect 29748 8606 30052 8608
rect 29748 8604 29795 8606
rect 30046 8604 30052 8606
rect 30116 8604 30122 8668
rect 29729 8603 29795 8604
rect 32206 8576 33006 8696
rect 13118 8468 13124 8532
rect 13188 8530 13194 8532
rect 30097 8530 30163 8533
rect 13188 8528 30163 8530
rect 13188 8472 30102 8528
rect 30158 8472 30163 8528
rect 13188 8470 30163 8472
rect 13188 8468 13194 8470
rect 30097 8467 30163 8470
rect 5717 8394 5783 8397
rect 19374 8394 19380 8396
rect 5717 8392 19380 8394
rect 5717 8336 5722 8392
rect 5778 8336 19380 8392
rect 5717 8334 19380 8336
rect 5717 8331 5783 8334
rect 19374 8332 19380 8334
rect 19444 8332 19450 8396
rect 19517 8394 19583 8397
rect 30373 8394 30439 8397
rect 19517 8392 30439 8394
rect 19517 8336 19522 8392
rect 19578 8336 30378 8392
rect 30434 8336 30439 8392
rect 19517 8334 30439 8336
rect 19517 8331 19583 8334
rect 30373 8331 30439 8334
rect 4787 8192 5103 8193
rect 0 8122 800 8152
rect 4787 8128 4793 8192
rect 4857 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5103 8192
rect 4787 8127 5103 8128
rect 12469 8192 12785 8193
rect 12469 8128 12475 8192
rect 12539 8128 12555 8192
rect 12619 8128 12635 8192
rect 12699 8128 12715 8192
rect 12779 8128 12785 8192
rect 12469 8127 12785 8128
rect 20151 8192 20467 8193
rect 20151 8128 20157 8192
rect 20221 8128 20237 8192
rect 20301 8128 20317 8192
rect 20381 8128 20397 8192
rect 20461 8128 20467 8192
rect 20151 8127 20467 8128
rect 27833 8192 28149 8193
rect 27833 8128 27839 8192
rect 27903 8128 27919 8192
rect 27983 8128 27999 8192
rect 28063 8128 28079 8192
rect 28143 8128 28149 8192
rect 27833 8127 28149 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 800 8062
rect 1577 8059 1643 8062
rect 11145 7986 11211 7989
rect 21030 7986 21036 7988
rect 11145 7984 21036 7986
rect 11145 7928 11150 7984
rect 11206 7928 21036 7984
rect 11145 7926 21036 7928
rect 11145 7923 11211 7926
rect 21030 7924 21036 7926
rect 21100 7924 21106 7988
rect 31293 7986 31359 7989
rect 32206 7986 33006 8016
rect 31293 7984 33006 7986
rect 31293 7928 31298 7984
rect 31354 7928 33006 7984
rect 31293 7926 33006 7928
rect 31293 7923 31359 7926
rect 32206 7896 33006 7926
rect 9438 7788 9444 7852
rect 9508 7850 9514 7852
rect 27613 7850 27679 7853
rect 9508 7848 27679 7850
rect 9508 7792 27618 7848
rect 27674 7792 27679 7848
rect 9508 7790 27679 7792
rect 9508 7788 9514 7790
rect 27613 7787 27679 7790
rect 8628 7648 8944 7649
rect 8628 7584 8634 7648
rect 8698 7584 8714 7648
rect 8778 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8944 7648
rect 8628 7583 8944 7584
rect 16310 7648 16626 7649
rect 16310 7584 16316 7648
rect 16380 7584 16396 7648
rect 16460 7584 16476 7648
rect 16540 7584 16556 7648
rect 16620 7584 16626 7648
rect 16310 7583 16626 7584
rect 23992 7648 24308 7649
rect 23992 7584 23998 7648
rect 24062 7584 24078 7648
rect 24142 7584 24158 7648
rect 24222 7584 24238 7648
rect 24302 7584 24308 7648
rect 23992 7583 24308 7584
rect 31674 7648 31990 7649
rect 31674 7584 31680 7648
rect 31744 7584 31760 7648
rect 31824 7584 31840 7648
rect 31904 7584 31920 7648
rect 31984 7584 31990 7648
rect 31674 7583 31990 7584
rect 14406 7380 14412 7444
rect 14476 7442 14482 7444
rect 24945 7442 25011 7445
rect 14476 7440 25011 7442
rect 14476 7384 24950 7440
rect 25006 7384 25011 7440
rect 14476 7382 25011 7384
rect 14476 7380 14482 7382
rect 24945 7379 25011 7382
rect 0 7216 800 7336
rect 11830 7244 11836 7308
rect 11900 7306 11906 7308
rect 29913 7306 29979 7309
rect 11900 7304 29979 7306
rect 11900 7248 29918 7304
rect 29974 7248 29979 7304
rect 11900 7246 29979 7248
rect 11900 7244 11906 7246
rect 29913 7243 29979 7246
rect 31293 7306 31359 7309
rect 32206 7306 33006 7336
rect 31293 7304 33006 7306
rect 31293 7248 31298 7304
rect 31354 7248 33006 7304
rect 31293 7246 33006 7248
rect 31293 7243 31359 7246
rect 32206 7216 33006 7246
rect 4787 7104 5103 7105
rect 4787 7040 4793 7104
rect 4857 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5103 7104
rect 4787 7039 5103 7040
rect 12469 7104 12785 7105
rect 12469 7040 12475 7104
rect 12539 7040 12555 7104
rect 12619 7040 12635 7104
rect 12699 7040 12715 7104
rect 12779 7040 12785 7104
rect 12469 7039 12785 7040
rect 20151 7104 20467 7105
rect 20151 7040 20157 7104
rect 20221 7040 20237 7104
rect 20301 7040 20317 7104
rect 20381 7040 20397 7104
rect 20461 7040 20467 7104
rect 20151 7039 20467 7040
rect 27833 7104 28149 7105
rect 27833 7040 27839 7104
rect 27903 7040 27919 7104
rect 27983 7040 27999 7104
rect 28063 7040 28079 7104
rect 28143 7040 28149 7104
rect 27833 7039 28149 7040
rect 14038 6836 14044 6900
rect 14108 6898 14114 6900
rect 29361 6898 29427 6901
rect 14108 6896 29427 6898
rect 14108 6840 29366 6896
rect 29422 6840 29427 6896
rect 14108 6838 29427 6840
rect 14108 6836 14114 6838
rect 29361 6835 29427 6838
rect 18638 6700 18644 6764
rect 18708 6762 18714 6764
rect 30465 6762 30531 6765
rect 18708 6760 30531 6762
rect 18708 6704 30470 6760
rect 30526 6704 30531 6760
rect 18708 6702 30531 6704
rect 18708 6700 18714 6702
rect 30465 6699 30531 6702
rect 8628 6560 8944 6561
rect 0 6490 800 6520
rect 8628 6496 8634 6560
rect 8698 6496 8714 6560
rect 8778 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8944 6560
rect 8628 6495 8944 6496
rect 16310 6560 16626 6561
rect 16310 6496 16316 6560
rect 16380 6496 16396 6560
rect 16460 6496 16476 6560
rect 16540 6496 16556 6560
rect 16620 6496 16626 6560
rect 16310 6495 16626 6496
rect 23992 6560 24308 6561
rect 23992 6496 23998 6560
rect 24062 6496 24078 6560
rect 24142 6496 24158 6560
rect 24222 6496 24238 6560
rect 24302 6496 24308 6560
rect 23992 6495 24308 6496
rect 31674 6560 31990 6561
rect 31674 6496 31680 6560
rect 31744 6496 31760 6560
rect 31824 6496 31840 6560
rect 31904 6496 31920 6560
rect 31984 6496 31990 6560
rect 32206 6536 33006 6656
rect 31674 6495 31990 6496
rect 1577 6490 1643 6493
rect 0 6488 1643 6490
rect 0 6432 1582 6488
rect 1638 6432 1643 6488
rect 0 6430 1643 6432
rect 0 6400 800 6430
rect 1577 6427 1643 6430
rect 2681 6218 2747 6221
rect 28717 6220 28783 6221
rect 28717 6218 28764 6220
rect 2681 6216 28764 6218
rect 28828 6218 28834 6220
rect 2681 6160 2686 6216
rect 2742 6160 28722 6216
rect 2681 6158 28764 6160
rect 2681 6155 2747 6158
rect 28717 6156 28764 6158
rect 28828 6158 28910 6218
rect 28828 6156 28834 6158
rect 28717 6155 28783 6156
rect 4787 6016 5103 6017
rect 4787 5952 4793 6016
rect 4857 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5103 6016
rect 4787 5951 5103 5952
rect 12469 6016 12785 6017
rect 12469 5952 12475 6016
rect 12539 5952 12555 6016
rect 12619 5952 12635 6016
rect 12699 5952 12715 6016
rect 12779 5952 12785 6016
rect 12469 5951 12785 5952
rect 20151 6016 20467 6017
rect 20151 5952 20157 6016
rect 20221 5952 20237 6016
rect 20301 5952 20317 6016
rect 20381 5952 20397 6016
rect 20461 5952 20467 6016
rect 20151 5951 20467 5952
rect 27833 6016 28149 6017
rect 27833 5952 27839 6016
rect 27903 5952 27919 6016
rect 27983 5952 27999 6016
rect 28063 5952 28079 6016
rect 28143 5952 28149 6016
rect 27833 5951 28149 5952
rect 31293 5946 31359 5949
rect 32206 5946 33006 5976
rect 31293 5944 33006 5946
rect 31293 5888 31298 5944
rect 31354 5888 33006 5944
rect 31293 5886 33006 5888
rect 31293 5883 31359 5886
rect 32206 5856 33006 5886
rect 0 5674 800 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 800 5614
rect 1577 5611 1643 5614
rect 8628 5472 8944 5473
rect 8628 5408 8634 5472
rect 8698 5408 8714 5472
rect 8778 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8944 5472
rect 8628 5407 8944 5408
rect 16310 5472 16626 5473
rect 16310 5408 16316 5472
rect 16380 5408 16396 5472
rect 16460 5408 16476 5472
rect 16540 5408 16556 5472
rect 16620 5408 16626 5472
rect 16310 5407 16626 5408
rect 23992 5472 24308 5473
rect 23992 5408 23998 5472
rect 24062 5408 24078 5472
rect 24142 5408 24158 5472
rect 24222 5408 24238 5472
rect 24302 5408 24308 5472
rect 23992 5407 24308 5408
rect 31674 5472 31990 5473
rect 31674 5408 31680 5472
rect 31744 5408 31760 5472
rect 31824 5408 31840 5472
rect 31904 5408 31920 5472
rect 31984 5408 31990 5472
rect 31674 5407 31990 5408
rect 5165 5266 5231 5269
rect 28942 5266 28948 5268
rect 5165 5264 28948 5266
rect 5165 5208 5170 5264
rect 5226 5208 28948 5264
rect 5165 5206 28948 5208
rect 5165 5203 5231 5206
rect 28942 5204 28948 5206
rect 29012 5204 29018 5268
rect 31293 5266 31359 5269
rect 32206 5266 33006 5296
rect 31293 5264 33006 5266
rect 31293 5208 31298 5264
rect 31354 5208 33006 5264
rect 31293 5206 33006 5208
rect 31293 5203 31359 5206
rect 32206 5176 33006 5206
rect 13486 5068 13492 5132
rect 13556 5130 13562 5132
rect 28625 5130 28691 5133
rect 13556 5128 28691 5130
rect 13556 5072 28630 5128
rect 28686 5072 28691 5128
rect 13556 5070 28691 5072
rect 13556 5068 13562 5070
rect 28625 5067 28691 5070
rect 4787 4928 5103 4929
rect 0 4768 800 4888
rect 4787 4864 4793 4928
rect 4857 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5103 4928
rect 4787 4863 5103 4864
rect 12469 4928 12785 4929
rect 12469 4864 12475 4928
rect 12539 4864 12555 4928
rect 12619 4864 12635 4928
rect 12699 4864 12715 4928
rect 12779 4864 12785 4928
rect 12469 4863 12785 4864
rect 20151 4928 20467 4929
rect 20151 4864 20157 4928
rect 20221 4864 20237 4928
rect 20301 4864 20317 4928
rect 20381 4864 20397 4928
rect 20461 4864 20467 4928
rect 20151 4863 20467 4864
rect 27833 4928 28149 4929
rect 27833 4864 27839 4928
rect 27903 4864 27919 4928
rect 27983 4864 27999 4928
rect 28063 4864 28079 4928
rect 28143 4864 28149 4928
rect 27833 4863 28149 4864
rect 15694 4660 15700 4724
rect 15764 4722 15770 4724
rect 29678 4722 29684 4724
rect 15764 4662 29684 4722
rect 15764 4660 15770 4662
rect 29678 4660 29684 4662
rect 29748 4660 29754 4724
rect 32206 4496 33006 4616
rect 8628 4384 8944 4385
rect 8628 4320 8634 4384
rect 8698 4320 8714 4384
rect 8778 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8944 4384
rect 8628 4319 8944 4320
rect 16310 4384 16626 4385
rect 16310 4320 16316 4384
rect 16380 4320 16396 4384
rect 16460 4320 16476 4384
rect 16540 4320 16556 4384
rect 16620 4320 16626 4384
rect 16310 4319 16626 4320
rect 23992 4384 24308 4385
rect 23992 4320 23998 4384
rect 24062 4320 24078 4384
rect 24142 4320 24158 4384
rect 24222 4320 24238 4384
rect 24302 4320 24308 4384
rect 23992 4319 24308 4320
rect 31674 4384 31990 4385
rect 31674 4320 31680 4384
rect 31744 4320 31760 4384
rect 31824 4320 31840 4384
rect 31904 4320 31920 4384
rect 31984 4320 31990 4384
rect 31674 4319 31990 4320
rect 0 4042 800 4072
rect 1577 4042 1643 4045
rect 0 4040 1643 4042
rect 0 3984 1582 4040
rect 1638 3984 1643 4040
rect 0 3982 1643 3984
rect 0 3952 800 3982
rect 1577 3979 1643 3982
rect 31293 3906 31359 3909
rect 32206 3906 33006 3936
rect 31293 3904 33006 3906
rect 31293 3848 31298 3904
rect 31354 3848 33006 3904
rect 31293 3846 33006 3848
rect 31293 3843 31359 3846
rect 4787 3840 5103 3841
rect 4787 3776 4793 3840
rect 4857 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5103 3840
rect 4787 3775 5103 3776
rect 12469 3840 12785 3841
rect 12469 3776 12475 3840
rect 12539 3776 12555 3840
rect 12619 3776 12635 3840
rect 12699 3776 12715 3840
rect 12779 3776 12785 3840
rect 12469 3775 12785 3776
rect 20151 3840 20467 3841
rect 20151 3776 20157 3840
rect 20221 3776 20237 3840
rect 20301 3776 20317 3840
rect 20381 3776 20397 3840
rect 20461 3776 20467 3840
rect 20151 3775 20467 3776
rect 27833 3840 28149 3841
rect 27833 3776 27839 3840
rect 27903 3776 27919 3840
rect 27983 3776 27999 3840
rect 28063 3776 28079 3840
rect 28143 3776 28149 3840
rect 32206 3816 33006 3846
rect 27833 3775 28149 3776
rect 31293 3498 31359 3501
rect 31293 3496 32138 3498
rect 31293 3440 31298 3496
rect 31354 3440 32138 3496
rect 31293 3438 32138 3440
rect 31293 3435 31359 3438
rect 8628 3296 8944 3297
rect 0 3226 800 3256
rect 8628 3232 8634 3296
rect 8698 3232 8714 3296
rect 8778 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8944 3296
rect 8628 3231 8944 3232
rect 16310 3296 16626 3297
rect 16310 3232 16316 3296
rect 16380 3232 16396 3296
rect 16460 3232 16476 3296
rect 16540 3232 16556 3296
rect 16620 3232 16626 3296
rect 16310 3231 16626 3232
rect 23992 3296 24308 3297
rect 23992 3232 23998 3296
rect 24062 3232 24078 3296
rect 24142 3232 24158 3296
rect 24222 3232 24238 3296
rect 24302 3232 24308 3296
rect 23992 3231 24308 3232
rect 31674 3296 31990 3297
rect 31674 3232 31680 3296
rect 31744 3232 31760 3296
rect 31824 3232 31840 3296
rect 31904 3232 31920 3296
rect 31984 3232 31990 3296
rect 31674 3231 31990 3232
rect 1577 3226 1643 3229
rect 0 3224 1643 3226
rect 0 3168 1582 3224
rect 1638 3168 1643 3224
rect 0 3166 1643 3168
rect 32078 3226 32138 3438
rect 32206 3226 33006 3256
rect 32078 3166 33006 3226
rect 0 3136 800 3166
rect 1577 3163 1643 3166
rect 32206 3136 33006 3166
rect 4787 2752 5103 2753
rect 4787 2688 4793 2752
rect 4857 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5103 2752
rect 4787 2687 5103 2688
rect 12469 2752 12785 2753
rect 12469 2688 12475 2752
rect 12539 2688 12555 2752
rect 12619 2688 12635 2752
rect 12699 2688 12715 2752
rect 12779 2688 12785 2752
rect 12469 2687 12785 2688
rect 20151 2752 20467 2753
rect 20151 2688 20157 2752
rect 20221 2688 20237 2752
rect 20301 2688 20317 2752
rect 20381 2688 20397 2752
rect 20461 2688 20467 2752
rect 20151 2687 20467 2688
rect 27833 2752 28149 2753
rect 27833 2688 27839 2752
rect 27903 2688 27919 2752
rect 27983 2688 27999 2752
rect 28063 2688 28079 2752
rect 28143 2688 28149 2752
rect 27833 2687 28149 2688
rect 32206 2456 33006 2576
rect 0 2320 800 2440
rect 8628 2208 8944 2209
rect 8628 2144 8634 2208
rect 8698 2144 8714 2208
rect 8778 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8944 2208
rect 8628 2143 8944 2144
rect 16310 2208 16626 2209
rect 16310 2144 16316 2208
rect 16380 2144 16396 2208
rect 16460 2144 16476 2208
rect 16540 2144 16556 2208
rect 16620 2144 16626 2208
rect 16310 2143 16626 2144
rect 23992 2208 24308 2209
rect 23992 2144 23998 2208
rect 24062 2144 24078 2208
rect 24142 2144 24158 2208
rect 24222 2144 24238 2208
rect 24302 2144 24308 2208
rect 23992 2143 24308 2144
rect 31674 2208 31990 2209
rect 31674 2144 31680 2208
rect 31744 2144 31760 2208
rect 31824 2144 31840 2208
rect 31904 2144 31920 2208
rect 31984 2144 31990 2208
rect 31674 2143 31990 2144
rect 0 1594 800 1624
rect 1577 1594 1643 1597
rect 0 1592 1643 1594
rect 0 1536 1582 1592
rect 1638 1536 1643 1592
rect 0 1534 1643 1536
rect 0 1504 800 1534
rect 1577 1531 1643 1534
rect 0 778 800 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 800 718
rect 1393 715 1459 718
<< via3 >>
rect 22140 34852 22204 34916
rect 20852 34716 20916 34780
rect 10180 34580 10244 34644
rect 26556 34172 26620 34236
rect 9260 34036 9324 34100
rect 12204 33764 12268 33828
rect 23796 33764 23860 33828
rect 15148 33356 15212 33420
rect 30236 33356 30300 33420
rect 16068 33220 16132 33284
rect 6316 33084 6380 33148
rect 30052 32812 30116 32876
rect 19932 32676 19996 32740
rect 8634 32668 8698 32672
rect 8634 32612 8638 32668
rect 8638 32612 8694 32668
rect 8694 32612 8698 32668
rect 8634 32608 8698 32612
rect 8714 32668 8778 32672
rect 8714 32612 8718 32668
rect 8718 32612 8774 32668
rect 8774 32612 8778 32668
rect 8714 32608 8778 32612
rect 8794 32668 8858 32672
rect 8794 32612 8798 32668
rect 8798 32612 8854 32668
rect 8854 32612 8858 32668
rect 8794 32608 8858 32612
rect 8874 32668 8938 32672
rect 8874 32612 8878 32668
rect 8878 32612 8934 32668
rect 8934 32612 8938 32668
rect 8874 32608 8938 32612
rect 16316 32668 16380 32672
rect 16316 32612 16320 32668
rect 16320 32612 16376 32668
rect 16376 32612 16380 32668
rect 16316 32608 16380 32612
rect 16396 32668 16460 32672
rect 16396 32612 16400 32668
rect 16400 32612 16456 32668
rect 16456 32612 16460 32668
rect 16396 32608 16460 32612
rect 16476 32668 16540 32672
rect 16476 32612 16480 32668
rect 16480 32612 16536 32668
rect 16536 32612 16540 32668
rect 16476 32608 16540 32612
rect 16556 32668 16620 32672
rect 16556 32612 16560 32668
rect 16560 32612 16616 32668
rect 16616 32612 16620 32668
rect 16556 32608 16620 32612
rect 23998 32668 24062 32672
rect 23998 32612 24002 32668
rect 24002 32612 24058 32668
rect 24058 32612 24062 32668
rect 23998 32608 24062 32612
rect 24078 32668 24142 32672
rect 24078 32612 24082 32668
rect 24082 32612 24138 32668
rect 24138 32612 24142 32668
rect 24078 32608 24142 32612
rect 24158 32668 24222 32672
rect 24158 32612 24162 32668
rect 24162 32612 24218 32668
rect 24218 32612 24222 32668
rect 24158 32608 24222 32612
rect 24238 32668 24302 32672
rect 24238 32612 24242 32668
rect 24242 32612 24298 32668
rect 24298 32612 24302 32668
rect 24238 32608 24302 32612
rect 31680 32668 31744 32672
rect 31680 32612 31684 32668
rect 31684 32612 31740 32668
rect 31740 32612 31744 32668
rect 31680 32608 31744 32612
rect 31760 32668 31824 32672
rect 31760 32612 31764 32668
rect 31764 32612 31820 32668
rect 31820 32612 31824 32668
rect 31760 32608 31824 32612
rect 31840 32668 31904 32672
rect 31840 32612 31844 32668
rect 31844 32612 31900 32668
rect 31900 32612 31904 32668
rect 31840 32608 31904 32612
rect 31920 32668 31984 32672
rect 31920 32612 31924 32668
rect 31924 32612 31980 32668
rect 31980 32612 31984 32668
rect 31920 32608 31984 32612
rect 22324 32540 22388 32604
rect 20668 32404 20732 32468
rect 4793 32124 4857 32128
rect 4793 32068 4797 32124
rect 4797 32068 4853 32124
rect 4853 32068 4857 32124
rect 4793 32064 4857 32068
rect 4873 32124 4937 32128
rect 4873 32068 4877 32124
rect 4877 32068 4933 32124
rect 4933 32068 4937 32124
rect 4873 32064 4937 32068
rect 4953 32124 5017 32128
rect 4953 32068 4957 32124
rect 4957 32068 5013 32124
rect 5013 32068 5017 32124
rect 4953 32064 5017 32068
rect 5033 32124 5097 32128
rect 5033 32068 5037 32124
rect 5037 32068 5093 32124
rect 5093 32068 5097 32124
rect 5033 32064 5097 32068
rect 12475 32124 12539 32128
rect 12475 32068 12479 32124
rect 12479 32068 12535 32124
rect 12535 32068 12539 32124
rect 12475 32064 12539 32068
rect 12555 32124 12619 32128
rect 12555 32068 12559 32124
rect 12559 32068 12615 32124
rect 12615 32068 12619 32124
rect 12555 32064 12619 32068
rect 12635 32124 12699 32128
rect 12635 32068 12639 32124
rect 12639 32068 12695 32124
rect 12695 32068 12699 32124
rect 12635 32064 12699 32068
rect 12715 32124 12779 32128
rect 12715 32068 12719 32124
rect 12719 32068 12775 32124
rect 12775 32068 12779 32124
rect 12715 32064 12779 32068
rect 20157 32124 20221 32128
rect 20157 32068 20161 32124
rect 20161 32068 20217 32124
rect 20217 32068 20221 32124
rect 20157 32064 20221 32068
rect 20237 32124 20301 32128
rect 20237 32068 20241 32124
rect 20241 32068 20297 32124
rect 20297 32068 20301 32124
rect 20237 32064 20301 32068
rect 20317 32124 20381 32128
rect 20317 32068 20321 32124
rect 20321 32068 20377 32124
rect 20377 32068 20381 32124
rect 20317 32064 20381 32068
rect 20397 32124 20461 32128
rect 20397 32068 20401 32124
rect 20401 32068 20457 32124
rect 20457 32068 20461 32124
rect 20397 32064 20461 32068
rect 27839 32124 27903 32128
rect 27839 32068 27843 32124
rect 27843 32068 27899 32124
rect 27899 32068 27903 32124
rect 27839 32064 27903 32068
rect 27919 32124 27983 32128
rect 27919 32068 27923 32124
rect 27923 32068 27979 32124
rect 27979 32068 27983 32124
rect 27919 32064 27983 32068
rect 27999 32124 28063 32128
rect 27999 32068 28003 32124
rect 28003 32068 28059 32124
rect 28059 32068 28063 32124
rect 27999 32064 28063 32068
rect 28079 32124 28143 32128
rect 28079 32068 28083 32124
rect 28083 32068 28139 32124
rect 28139 32068 28143 32124
rect 28079 32064 28143 32068
rect 26188 31996 26252 32060
rect 8156 31860 8220 31924
rect 21956 31860 22020 31924
rect 25452 31724 25516 31788
rect 24532 31648 24596 31652
rect 24532 31592 24546 31648
rect 24546 31592 24596 31648
rect 24532 31588 24596 31592
rect 26004 31588 26068 31652
rect 27292 31588 27356 31652
rect 28764 31588 28828 31652
rect 8634 31580 8698 31584
rect 8634 31524 8638 31580
rect 8638 31524 8694 31580
rect 8694 31524 8698 31580
rect 8634 31520 8698 31524
rect 8714 31580 8778 31584
rect 8714 31524 8718 31580
rect 8718 31524 8774 31580
rect 8774 31524 8778 31580
rect 8714 31520 8778 31524
rect 8794 31580 8858 31584
rect 8794 31524 8798 31580
rect 8798 31524 8854 31580
rect 8854 31524 8858 31580
rect 8794 31520 8858 31524
rect 8874 31580 8938 31584
rect 8874 31524 8878 31580
rect 8878 31524 8934 31580
rect 8934 31524 8938 31580
rect 8874 31520 8938 31524
rect 16316 31580 16380 31584
rect 16316 31524 16320 31580
rect 16320 31524 16376 31580
rect 16376 31524 16380 31580
rect 16316 31520 16380 31524
rect 16396 31580 16460 31584
rect 16396 31524 16400 31580
rect 16400 31524 16456 31580
rect 16456 31524 16460 31580
rect 16396 31520 16460 31524
rect 16476 31580 16540 31584
rect 16476 31524 16480 31580
rect 16480 31524 16536 31580
rect 16536 31524 16540 31580
rect 16476 31520 16540 31524
rect 16556 31580 16620 31584
rect 16556 31524 16560 31580
rect 16560 31524 16616 31580
rect 16616 31524 16620 31580
rect 16556 31520 16620 31524
rect 23998 31580 24062 31584
rect 23998 31524 24002 31580
rect 24002 31524 24058 31580
rect 24058 31524 24062 31580
rect 23998 31520 24062 31524
rect 24078 31580 24142 31584
rect 24078 31524 24082 31580
rect 24082 31524 24138 31580
rect 24138 31524 24142 31580
rect 24078 31520 24142 31524
rect 24158 31580 24222 31584
rect 24158 31524 24162 31580
rect 24162 31524 24218 31580
rect 24218 31524 24222 31580
rect 24158 31520 24222 31524
rect 24238 31580 24302 31584
rect 24238 31524 24242 31580
rect 24242 31524 24298 31580
rect 24298 31524 24302 31580
rect 24238 31520 24302 31524
rect 31680 31580 31744 31584
rect 31680 31524 31684 31580
rect 31684 31524 31740 31580
rect 31740 31524 31744 31580
rect 31680 31520 31744 31524
rect 31760 31580 31824 31584
rect 31760 31524 31764 31580
rect 31764 31524 31820 31580
rect 31820 31524 31824 31580
rect 31760 31520 31824 31524
rect 31840 31580 31904 31584
rect 31840 31524 31844 31580
rect 31844 31524 31900 31580
rect 31900 31524 31904 31580
rect 31840 31520 31904 31524
rect 31920 31580 31984 31584
rect 31920 31524 31924 31580
rect 31924 31524 31980 31580
rect 31980 31524 31984 31580
rect 31920 31520 31984 31524
rect 22508 31452 22572 31516
rect 17724 31316 17788 31380
rect 10732 31180 10796 31244
rect 22692 31180 22756 31244
rect 32260 31316 32324 31380
rect 30788 31180 30852 31244
rect 18092 31044 18156 31108
rect 25268 31044 25332 31108
rect 29316 31044 29380 31108
rect 4793 31036 4857 31040
rect 4793 30980 4797 31036
rect 4797 30980 4853 31036
rect 4853 30980 4857 31036
rect 4793 30976 4857 30980
rect 4873 31036 4937 31040
rect 4873 30980 4877 31036
rect 4877 30980 4933 31036
rect 4933 30980 4937 31036
rect 4873 30976 4937 30980
rect 4953 31036 5017 31040
rect 4953 30980 4957 31036
rect 4957 30980 5013 31036
rect 5013 30980 5017 31036
rect 4953 30976 5017 30980
rect 5033 31036 5097 31040
rect 5033 30980 5037 31036
rect 5037 30980 5093 31036
rect 5093 30980 5097 31036
rect 5033 30976 5097 30980
rect 12475 31036 12539 31040
rect 12475 30980 12479 31036
rect 12479 30980 12535 31036
rect 12535 30980 12539 31036
rect 12475 30976 12539 30980
rect 12555 31036 12619 31040
rect 12555 30980 12559 31036
rect 12559 30980 12615 31036
rect 12615 30980 12619 31036
rect 12555 30976 12619 30980
rect 12635 31036 12699 31040
rect 12635 30980 12639 31036
rect 12639 30980 12695 31036
rect 12695 30980 12699 31036
rect 12635 30976 12699 30980
rect 12715 31036 12779 31040
rect 12715 30980 12719 31036
rect 12719 30980 12775 31036
rect 12775 30980 12779 31036
rect 12715 30976 12779 30980
rect 20157 31036 20221 31040
rect 20157 30980 20161 31036
rect 20161 30980 20217 31036
rect 20217 30980 20221 31036
rect 20157 30976 20221 30980
rect 20237 31036 20301 31040
rect 20237 30980 20241 31036
rect 20241 30980 20297 31036
rect 20297 30980 20301 31036
rect 20237 30976 20301 30980
rect 20317 31036 20381 31040
rect 20317 30980 20321 31036
rect 20321 30980 20377 31036
rect 20377 30980 20381 31036
rect 20317 30976 20381 30980
rect 20397 31036 20461 31040
rect 20397 30980 20401 31036
rect 20401 30980 20457 31036
rect 20457 30980 20461 31036
rect 20397 30976 20461 30980
rect 27839 31036 27903 31040
rect 27839 30980 27843 31036
rect 27843 30980 27899 31036
rect 27899 30980 27903 31036
rect 27839 30976 27903 30980
rect 27919 31036 27983 31040
rect 27919 30980 27923 31036
rect 27923 30980 27979 31036
rect 27979 30980 27983 31036
rect 27919 30976 27983 30980
rect 27999 31036 28063 31040
rect 27999 30980 28003 31036
rect 28003 30980 28059 31036
rect 28059 30980 28063 31036
rect 27999 30976 28063 30980
rect 28079 31036 28143 31040
rect 28079 30980 28083 31036
rect 28083 30980 28139 31036
rect 28139 30980 28143 31036
rect 28079 30976 28143 30980
rect 14228 30908 14292 30972
rect 15516 30908 15580 30972
rect 28396 30968 28460 30972
rect 28396 30912 28446 30968
rect 28446 30912 28460 30968
rect 28396 30908 28460 30912
rect 6684 30772 6748 30836
rect 6868 30636 6932 30700
rect 11468 30636 11532 30700
rect 19748 30772 19812 30836
rect 19196 30636 19260 30700
rect 25820 30772 25884 30836
rect 27476 30772 27540 30836
rect 23428 30500 23492 30564
rect 27108 30636 27172 30700
rect 30420 30772 30484 30836
rect 8634 30492 8698 30496
rect 8634 30436 8638 30492
rect 8638 30436 8694 30492
rect 8694 30436 8698 30492
rect 8634 30432 8698 30436
rect 8714 30492 8778 30496
rect 8714 30436 8718 30492
rect 8718 30436 8774 30492
rect 8774 30436 8778 30492
rect 8714 30432 8778 30436
rect 8794 30492 8858 30496
rect 8794 30436 8798 30492
rect 8798 30436 8854 30492
rect 8854 30436 8858 30492
rect 8794 30432 8858 30436
rect 8874 30492 8938 30496
rect 8874 30436 8878 30492
rect 8878 30436 8934 30492
rect 8934 30436 8938 30492
rect 8874 30432 8938 30436
rect 16316 30492 16380 30496
rect 16316 30436 16320 30492
rect 16320 30436 16376 30492
rect 16376 30436 16380 30492
rect 16316 30432 16380 30436
rect 16396 30492 16460 30496
rect 16396 30436 16400 30492
rect 16400 30436 16456 30492
rect 16456 30436 16460 30492
rect 16396 30432 16460 30436
rect 16476 30492 16540 30496
rect 16476 30436 16480 30492
rect 16480 30436 16536 30492
rect 16536 30436 16540 30492
rect 16476 30432 16540 30436
rect 16556 30492 16620 30496
rect 16556 30436 16560 30492
rect 16560 30436 16616 30492
rect 16616 30436 16620 30492
rect 16556 30432 16620 30436
rect 23998 30492 24062 30496
rect 23998 30436 24002 30492
rect 24002 30436 24058 30492
rect 24058 30436 24062 30492
rect 23998 30432 24062 30436
rect 24078 30492 24142 30496
rect 24078 30436 24082 30492
rect 24082 30436 24138 30492
rect 24138 30436 24142 30492
rect 24078 30432 24142 30436
rect 24158 30492 24222 30496
rect 24158 30436 24162 30492
rect 24162 30436 24218 30492
rect 24218 30436 24222 30492
rect 24158 30432 24222 30436
rect 24238 30492 24302 30496
rect 24238 30436 24242 30492
rect 24242 30436 24298 30492
rect 24298 30436 24302 30492
rect 24238 30432 24302 30436
rect 11836 30364 11900 30428
rect 14412 30364 14476 30428
rect 19012 30364 19076 30428
rect 19932 30364 19996 30428
rect 21036 30364 21100 30428
rect 26740 30500 26804 30564
rect 26924 30500 26988 30564
rect 31680 30492 31744 30496
rect 31680 30436 31684 30492
rect 31684 30436 31740 30492
rect 31740 30436 31744 30492
rect 31680 30432 31744 30436
rect 31760 30492 31824 30496
rect 31760 30436 31764 30492
rect 31764 30436 31820 30492
rect 31820 30436 31824 30492
rect 31760 30432 31824 30436
rect 31840 30492 31904 30496
rect 31840 30436 31844 30492
rect 31844 30436 31900 30492
rect 31900 30436 31904 30492
rect 31840 30432 31904 30436
rect 31920 30492 31984 30496
rect 31920 30436 31924 30492
rect 31924 30436 31980 30492
rect 31980 30436 31984 30492
rect 31920 30432 31984 30436
rect 27660 30364 27724 30428
rect 30604 30424 30668 30428
rect 30604 30368 30618 30424
rect 30618 30368 30668 30424
rect 30604 30364 30668 30368
rect 19380 30228 19444 30292
rect 22876 30228 22940 30292
rect 7052 30092 7116 30156
rect 15148 30092 15212 30156
rect 25084 30092 25148 30156
rect 25636 30092 25700 30156
rect 17908 29956 17972 30020
rect 26372 30016 26436 30020
rect 26372 29960 26386 30016
rect 26386 29960 26436 30016
rect 26372 29956 26436 29960
rect 27292 29956 27356 30020
rect 28258 29956 28322 30020
rect 32628 29956 32692 30020
rect 4793 29948 4857 29952
rect 4793 29892 4797 29948
rect 4797 29892 4853 29948
rect 4853 29892 4857 29948
rect 4793 29888 4857 29892
rect 4873 29948 4937 29952
rect 4873 29892 4877 29948
rect 4877 29892 4933 29948
rect 4933 29892 4937 29948
rect 4873 29888 4937 29892
rect 4953 29948 5017 29952
rect 4953 29892 4957 29948
rect 4957 29892 5013 29948
rect 5013 29892 5017 29948
rect 4953 29888 5017 29892
rect 5033 29948 5097 29952
rect 5033 29892 5037 29948
rect 5037 29892 5093 29948
rect 5093 29892 5097 29948
rect 5033 29888 5097 29892
rect 12475 29948 12539 29952
rect 12475 29892 12479 29948
rect 12479 29892 12535 29948
rect 12535 29892 12539 29948
rect 12475 29888 12539 29892
rect 12555 29948 12619 29952
rect 12555 29892 12559 29948
rect 12559 29892 12615 29948
rect 12615 29892 12619 29948
rect 12555 29888 12619 29892
rect 12635 29948 12699 29952
rect 12635 29892 12639 29948
rect 12639 29892 12695 29948
rect 12695 29892 12699 29948
rect 12635 29888 12699 29892
rect 12715 29948 12779 29952
rect 12715 29892 12719 29948
rect 12719 29892 12775 29948
rect 12775 29892 12779 29948
rect 12715 29888 12779 29892
rect 20157 29948 20221 29952
rect 20157 29892 20161 29948
rect 20161 29892 20217 29948
rect 20217 29892 20221 29948
rect 20157 29888 20221 29892
rect 20237 29948 20301 29952
rect 20237 29892 20241 29948
rect 20241 29892 20297 29948
rect 20297 29892 20301 29948
rect 20237 29888 20301 29892
rect 20317 29948 20381 29952
rect 20317 29892 20321 29948
rect 20321 29892 20377 29948
rect 20377 29892 20381 29948
rect 20317 29888 20381 29892
rect 20397 29948 20461 29952
rect 20397 29892 20401 29948
rect 20401 29892 20457 29948
rect 20457 29892 20461 29948
rect 20397 29888 20461 29892
rect 27839 29948 27903 29952
rect 27839 29892 27843 29948
rect 27843 29892 27899 29948
rect 27899 29892 27903 29948
rect 27839 29888 27903 29892
rect 27919 29948 27983 29952
rect 27919 29892 27923 29948
rect 27923 29892 27979 29948
rect 27979 29892 27983 29948
rect 27919 29888 27983 29892
rect 27999 29948 28063 29952
rect 27999 29892 28003 29948
rect 28003 29892 28059 29948
rect 28059 29892 28063 29948
rect 27999 29888 28063 29892
rect 28079 29948 28143 29952
rect 28079 29892 28083 29948
rect 28083 29892 28139 29948
rect 28139 29892 28143 29948
rect 28079 29888 28143 29892
rect 17172 29820 17236 29884
rect 27292 29880 27356 29884
rect 27292 29824 27342 29880
rect 27342 29824 27356 29880
rect 12940 29684 13004 29748
rect 18276 29684 18340 29748
rect 27292 29820 27356 29824
rect 29500 29820 29564 29884
rect 21772 29684 21836 29748
rect 25084 29684 25148 29748
rect 25452 29684 25516 29748
rect 28580 29684 28644 29748
rect 17540 29412 17604 29476
rect 21404 29472 21468 29476
rect 22508 29548 22572 29612
rect 21404 29416 21454 29472
rect 21454 29416 21468 29472
rect 21404 29412 21468 29416
rect 23060 29412 23124 29476
rect 25452 29412 25516 29476
rect 25636 29472 25700 29476
rect 25636 29416 25650 29472
rect 25650 29416 25700 29472
rect 25636 29412 25700 29416
rect 26004 29412 26068 29476
rect 26924 29412 26988 29476
rect 28948 29548 29012 29612
rect 31156 29548 31220 29612
rect 29132 29412 29196 29476
rect 8634 29404 8698 29408
rect 8634 29348 8638 29404
rect 8638 29348 8694 29404
rect 8694 29348 8698 29404
rect 8634 29344 8698 29348
rect 8714 29404 8778 29408
rect 8714 29348 8718 29404
rect 8718 29348 8774 29404
rect 8774 29348 8778 29404
rect 8714 29344 8778 29348
rect 8794 29404 8858 29408
rect 8794 29348 8798 29404
rect 8798 29348 8854 29404
rect 8854 29348 8858 29404
rect 8794 29344 8858 29348
rect 8874 29404 8938 29408
rect 8874 29348 8878 29404
rect 8878 29348 8934 29404
rect 8934 29348 8938 29404
rect 8874 29344 8938 29348
rect 16316 29404 16380 29408
rect 16316 29348 16320 29404
rect 16320 29348 16376 29404
rect 16376 29348 16380 29404
rect 16316 29344 16380 29348
rect 16396 29404 16460 29408
rect 16396 29348 16400 29404
rect 16400 29348 16456 29404
rect 16456 29348 16460 29404
rect 16396 29344 16460 29348
rect 16476 29404 16540 29408
rect 16476 29348 16480 29404
rect 16480 29348 16536 29404
rect 16536 29348 16540 29404
rect 16476 29344 16540 29348
rect 16556 29404 16620 29408
rect 16556 29348 16560 29404
rect 16560 29348 16616 29404
rect 16616 29348 16620 29404
rect 16556 29344 16620 29348
rect 23998 29404 24062 29408
rect 23998 29348 24002 29404
rect 24002 29348 24058 29404
rect 24058 29348 24062 29404
rect 23998 29344 24062 29348
rect 24078 29404 24142 29408
rect 24078 29348 24082 29404
rect 24082 29348 24138 29404
rect 24138 29348 24142 29404
rect 24078 29344 24142 29348
rect 24158 29404 24222 29408
rect 24158 29348 24162 29404
rect 24162 29348 24218 29404
rect 24218 29348 24222 29404
rect 24158 29344 24222 29348
rect 24238 29404 24302 29408
rect 24238 29348 24242 29404
rect 24242 29348 24298 29404
rect 24298 29348 24302 29404
rect 24238 29344 24302 29348
rect 31680 29404 31744 29408
rect 31680 29348 31684 29404
rect 31684 29348 31740 29404
rect 31740 29348 31744 29404
rect 31680 29344 31744 29348
rect 31760 29404 31824 29408
rect 31760 29348 31764 29404
rect 31764 29348 31820 29404
rect 31820 29348 31824 29404
rect 31760 29344 31824 29348
rect 31840 29404 31904 29408
rect 31840 29348 31844 29404
rect 31844 29348 31900 29404
rect 31900 29348 31904 29404
rect 31840 29344 31904 29348
rect 31920 29404 31984 29408
rect 31920 29348 31924 29404
rect 31924 29348 31980 29404
rect 31980 29348 31984 29404
rect 31920 29344 31984 29348
rect 13492 29276 13556 29340
rect 21220 29276 21284 29340
rect 21588 29276 21652 29340
rect 21956 29276 22020 29340
rect 23244 29336 23308 29340
rect 23244 29280 23258 29336
rect 23258 29280 23308 29336
rect 23244 29276 23308 29280
rect 23612 29336 23676 29340
rect 23612 29280 23662 29336
rect 23662 29280 23676 29336
rect 23612 29276 23676 29280
rect 28212 29276 28276 29340
rect 29684 29276 29748 29340
rect 9444 29004 9508 29068
rect 15700 29004 15764 29068
rect 19932 29140 19996 29204
rect 21956 29140 22020 29204
rect 26556 29140 26620 29204
rect 26924 29140 26988 29204
rect 24900 29004 24964 29068
rect 26924 29004 26988 29068
rect 27292 29004 27356 29068
rect 19564 28868 19628 28932
rect 22692 28868 22756 28932
rect 31524 29004 31588 29068
rect 4793 28860 4857 28864
rect 4793 28804 4797 28860
rect 4797 28804 4853 28860
rect 4853 28804 4857 28860
rect 4793 28800 4857 28804
rect 4873 28860 4937 28864
rect 4873 28804 4877 28860
rect 4877 28804 4933 28860
rect 4933 28804 4937 28860
rect 4873 28800 4937 28804
rect 4953 28860 5017 28864
rect 4953 28804 4957 28860
rect 4957 28804 5013 28860
rect 5013 28804 5017 28860
rect 4953 28800 5017 28804
rect 5033 28860 5097 28864
rect 5033 28804 5037 28860
rect 5037 28804 5093 28860
rect 5093 28804 5097 28860
rect 5033 28800 5097 28804
rect 12475 28860 12539 28864
rect 12475 28804 12479 28860
rect 12479 28804 12535 28860
rect 12535 28804 12539 28860
rect 12475 28800 12539 28804
rect 12555 28860 12619 28864
rect 12555 28804 12559 28860
rect 12559 28804 12615 28860
rect 12615 28804 12619 28860
rect 12555 28800 12619 28804
rect 12635 28860 12699 28864
rect 12635 28804 12639 28860
rect 12639 28804 12695 28860
rect 12695 28804 12699 28860
rect 12635 28800 12699 28804
rect 12715 28860 12779 28864
rect 12715 28804 12719 28860
rect 12719 28804 12775 28860
rect 12775 28804 12779 28860
rect 12715 28800 12779 28804
rect 20157 28860 20221 28864
rect 20157 28804 20161 28860
rect 20161 28804 20217 28860
rect 20217 28804 20221 28860
rect 20157 28800 20221 28804
rect 20237 28860 20301 28864
rect 20237 28804 20241 28860
rect 20241 28804 20297 28860
rect 20297 28804 20301 28860
rect 20237 28800 20301 28804
rect 20317 28860 20381 28864
rect 20317 28804 20321 28860
rect 20321 28804 20377 28860
rect 20377 28804 20381 28860
rect 20317 28800 20381 28804
rect 20397 28860 20461 28864
rect 20397 28804 20401 28860
rect 20401 28804 20457 28860
rect 20457 28804 20461 28860
rect 20397 28800 20461 28804
rect 27839 28860 27903 28864
rect 27839 28804 27843 28860
rect 27843 28804 27899 28860
rect 27899 28804 27903 28860
rect 27839 28800 27903 28804
rect 27919 28860 27983 28864
rect 27919 28804 27923 28860
rect 27923 28804 27979 28860
rect 27979 28804 27983 28860
rect 27919 28800 27983 28804
rect 27999 28860 28063 28864
rect 27999 28804 28003 28860
rect 28003 28804 28059 28860
rect 28059 28804 28063 28860
rect 27999 28800 28063 28804
rect 28079 28860 28143 28864
rect 28079 28804 28083 28860
rect 28083 28804 28139 28860
rect 28139 28804 28143 28860
rect 28079 28800 28143 28804
rect 20852 28732 20916 28796
rect 28764 28868 28828 28932
rect 32444 28732 32508 28796
rect 19012 28596 19076 28660
rect 19748 28596 19812 28660
rect 16988 28460 17052 28524
rect 26004 28596 26068 28660
rect 29316 28596 29380 28660
rect 29500 28656 29564 28660
rect 29500 28600 29514 28656
rect 29514 28600 29564 28656
rect 29500 28596 29564 28600
rect 21956 28460 22020 28524
rect 22876 28460 22940 28524
rect 24532 28324 24596 28388
rect 24900 28324 24964 28388
rect 25084 28324 25148 28388
rect 26004 28324 26068 28388
rect 26188 28384 26252 28388
rect 26188 28328 26238 28384
rect 26238 28328 26252 28384
rect 26188 28324 26252 28328
rect 28212 28324 28276 28388
rect 28580 28324 28644 28388
rect 29500 28324 29564 28388
rect 31340 28324 31404 28388
rect 8634 28316 8698 28320
rect 8634 28260 8638 28316
rect 8638 28260 8694 28316
rect 8694 28260 8698 28316
rect 8634 28256 8698 28260
rect 8714 28316 8778 28320
rect 8714 28260 8718 28316
rect 8718 28260 8774 28316
rect 8774 28260 8778 28316
rect 8714 28256 8778 28260
rect 8794 28316 8858 28320
rect 8794 28260 8798 28316
rect 8798 28260 8854 28316
rect 8854 28260 8858 28316
rect 8794 28256 8858 28260
rect 8874 28316 8938 28320
rect 8874 28260 8878 28316
rect 8878 28260 8934 28316
rect 8934 28260 8938 28316
rect 8874 28256 8938 28260
rect 16316 28316 16380 28320
rect 16316 28260 16320 28316
rect 16320 28260 16376 28316
rect 16376 28260 16380 28316
rect 16316 28256 16380 28260
rect 16396 28316 16460 28320
rect 16396 28260 16400 28316
rect 16400 28260 16456 28316
rect 16456 28260 16460 28316
rect 16396 28256 16460 28260
rect 16476 28316 16540 28320
rect 16476 28260 16480 28316
rect 16480 28260 16536 28316
rect 16536 28260 16540 28316
rect 16476 28256 16540 28260
rect 16556 28316 16620 28320
rect 16556 28260 16560 28316
rect 16560 28260 16616 28316
rect 16616 28260 16620 28316
rect 16556 28256 16620 28260
rect 23998 28316 24062 28320
rect 23998 28260 24002 28316
rect 24002 28260 24058 28316
rect 24058 28260 24062 28316
rect 23998 28256 24062 28260
rect 24078 28316 24142 28320
rect 24078 28260 24082 28316
rect 24082 28260 24138 28316
rect 24138 28260 24142 28316
rect 24078 28256 24142 28260
rect 24158 28316 24222 28320
rect 24158 28260 24162 28316
rect 24162 28260 24218 28316
rect 24218 28260 24222 28316
rect 24158 28256 24222 28260
rect 24238 28316 24302 28320
rect 24238 28260 24242 28316
rect 24242 28260 24298 28316
rect 24298 28260 24302 28316
rect 24238 28256 24302 28260
rect 31680 28316 31744 28320
rect 31680 28260 31684 28316
rect 31684 28260 31740 28316
rect 31740 28260 31744 28316
rect 31680 28256 31744 28260
rect 31760 28316 31824 28320
rect 31760 28260 31764 28316
rect 31764 28260 31820 28316
rect 31820 28260 31824 28316
rect 31760 28256 31824 28260
rect 31840 28316 31904 28320
rect 31840 28260 31844 28316
rect 31844 28260 31900 28316
rect 31900 28260 31904 28316
rect 31840 28256 31904 28260
rect 31920 28316 31984 28320
rect 31920 28260 31924 28316
rect 31924 28260 31980 28316
rect 31980 28260 31984 28316
rect 31920 28256 31984 28260
rect 14780 28188 14844 28252
rect 16804 28188 16868 28252
rect 18460 28188 18524 28252
rect 18644 28248 18708 28252
rect 18644 28192 18658 28248
rect 18658 28192 18708 28248
rect 18644 28188 18708 28192
rect 22324 28188 22388 28252
rect 22692 28188 22756 28252
rect 23612 28248 23676 28252
rect 23612 28192 23662 28248
rect 23662 28192 23676 28248
rect 14596 28112 14660 28116
rect 14596 28056 14610 28112
rect 14610 28056 14660 28112
rect 14596 28052 14660 28056
rect 15884 28052 15948 28116
rect 23612 28188 23676 28192
rect 25820 28188 25884 28252
rect 26004 28188 26068 28252
rect 29316 28188 29380 28252
rect 25636 28052 25700 28116
rect 13308 27916 13372 27980
rect 28580 27916 28644 27980
rect 32076 27916 32140 27980
rect 13676 27780 13740 27844
rect 20668 27780 20732 27844
rect 21588 27840 21652 27844
rect 21588 27784 21602 27840
rect 21602 27784 21652 27840
rect 21588 27780 21652 27784
rect 21772 27840 21836 27844
rect 21772 27784 21822 27840
rect 21822 27784 21836 27840
rect 21772 27780 21836 27784
rect 22140 27780 22204 27844
rect 22692 27780 22756 27844
rect 24900 27780 24964 27844
rect 25268 27840 25332 27844
rect 25268 27784 25282 27840
rect 25282 27784 25332 27840
rect 25268 27780 25332 27784
rect 26372 27780 26436 27844
rect 26924 27780 26988 27844
rect 27660 27840 27724 27844
rect 27660 27784 27710 27840
rect 27710 27784 27724 27840
rect 27660 27780 27724 27784
rect 29868 27780 29932 27844
rect 4793 27772 4857 27776
rect 4793 27716 4797 27772
rect 4797 27716 4853 27772
rect 4853 27716 4857 27772
rect 4793 27712 4857 27716
rect 4873 27772 4937 27776
rect 4873 27716 4877 27772
rect 4877 27716 4933 27772
rect 4933 27716 4937 27772
rect 4873 27712 4937 27716
rect 4953 27772 5017 27776
rect 4953 27716 4957 27772
rect 4957 27716 5013 27772
rect 5013 27716 5017 27772
rect 4953 27712 5017 27716
rect 5033 27772 5097 27776
rect 5033 27716 5037 27772
rect 5037 27716 5093 27772
rect 5093 27716 5097 27772
rect 5033 27712 5097 27716
rect 12475 27772 12539 27776
rect 12475 27716 12479 27772
rect 12479 27716 12535 27772
rect 12535 27716 12539 27772
rect 12475 27712 12539 27716
rect 12555 27772 12619 27776
rect 12555 27716 12559 27772
rect 12559 27716 12615 27772
rect 12615 27716 12619 27772
rect 12555 27712 12619 27716
rect 12635 27772 12699 27776
rect 12635 27716 12639 27772
rect 12639 27716 12695 27772
rect 12695 27716 12699 27772
rect 12635 27712 12699 27716
rect 12715 27772 12779 27776
rect 12715 27716 12719 27772
rect 12719 27716 12775 27772
rect 12775 27716 12779 27772
rect 12715 27712 12779 27716
rect 20157 27772 20221 27776
rect 20157 27716 20161 27772
rect 20161 27716 20217 27772
rect 20217 27716 20221 27772
rect 20157 27712 20221 27716
rect 20237 27772 20301 27776
rect 20237 27716 20241 27772
rect 20241 27716 20297 27772
rect 20297 27716 20301 27772
rect 20237 27712 20301 27716
rect 20317 27772 20381 27776
rect 20317 27716 20321 27772
rect 20321 27716 20377 27772
rect 20377 27716 20381 27772
rect 20317 27712 20381 27716
rect 20397 27772 20461 27776
rect 20397 27716 20401 27772
rect 20401 27716 20457 27772
rect 20457 27716 20461 27772
rect 20397 27712 20461 27716
rect 27839 27772 27903 27776
rect 27839 27716 27843 27772
rect 27843 27716 27899 27772
rect 27899 27716 27903 27772
rect 27839 27712 27903 27716
rect 27919 27772 27983 27776
rect 27919 27716 27923 27772
rect 27923 27716 27979 27772
rect 27979 27716 27983 27772
rect 27919 27712 27983 27716
rect 27999 27772 28063 27776
rect 27999 27716 28003 27772
rect 28003 27716 28059 27772
rect 28059 27716 28063 27772
rect 27999 27712 28063 27716
rect 28079 27772 28143 27776
rect 28079 27716 28083 27772
rect 28083 27716 28139 27772
rect 28139 27716 28143 27772
rect 28079 27712 28143 27716
rect 12020 27508 12084 27572
rect 19196 27644 19260 27708
rect 20852 27644 20916 27708
rect 22140 27644 22204 27708
rect 22508 27644 22572 27708
rect 16068 27508 16132 27572
rect 18460 27508 18524 27572
rect 19196 27508 19260 27572
rect 21220 27508 21284 27572
rect 22508 27568 22572 27572
rect 22508 27512 22522 27568
rect 22522 27512 22572 27568
rect 22508 27508 22572 27512
rect 21220 27372 21284 27436
rect 27660 27704 27724 27708
rect 27660 27648 27674 27704
rect 27674 27648 27724 27704
rect 27660 27644 27724 27648
rect 28258 27644 28322 27708
rect 29500 27644 29564 27708
rect 23244 27568 23308 27572
rect 23244 27512 23258 27568
rect 23258 27512 23308 27568
rect 23244 27508 23308 27512
rect 23428 27568 23492 27572
rect 23428 27512 23442 27568
rect 23442 27512 23492 27568
rect 23428 27508 23492 27512
rect 23612 27508 23676 27572
rect 24716 27508 24780 27572
rect 17356 27236 17420 27300
rect 8634 27228 8698 27232
rect 8634 27172 8638 27228
rect 8638 27172 8694 27228
rect 8694 27172 8698 27228
rect 8634 27168 8698 27172
rect 8714 27228 8778 27232
rect 8714 27172 8718 27228
rect 8718 27172 8774 27228
rect 8774 27172 8778 27228
rect 8714 27168 8778 27172
rect 8794 27228 8858 27232
rect 8794 27172 8798 27228
rect 8798 27172 8854 27228
rect 8854 27172 8858 27228
rect 8794 27168 8858 27172
rect 8874 27228 8938 27232
rect 8874 27172 8878 27228
rect 8878 27172 8934 27228
rect 8934 27172 8938 27228
rect 8874 27168 8938 27172
rect 16316 27228 16380 27232
rect 16316 27172 16320 27228
rect 16320 27172 16376 27228
rect 16376 27172 16380 27228
rect 16316 27168 16380 27172
rect 16396 27228 16460 27232
rect 16396 27172 16400 27228
rect 16400 27172 16456 27228
rect 16456 27172 16460 27228
rect 16396 27168 16460 27172
rect 16476 27228 16540 27232
rect 16476 27172 16480 27228
rect 16480 27172 16536 27228
rect 16536 27172 16540 27228
rect 16476 27168 16540 27172
rect 16556 27228 16620 27232
rect 16556 27172 16560 27228
rect 16560 27172 16616 27228
rect 16616 27172 16620 27228
rect 16556 27168 16620 27172
rect 16068 27100 16132 27164
rect 23612 27100 23676 27164
rect 25084 27372 25148 27436
rect 26924 27508 26988 27572
rect 31524 27508 31588 27572
rect 30972 27372 31036 27436
rect 26740 27236 26804 27300
rect 29684 27236 29748 27300
rect 30052 27236 30116 27300
rect 23998 27228 24062 27232
rect 23998 27172 24002 27228
rect 24002 27172 24058 27228
rect 24058 27172 24062 27228
rect 23998 27168 24062 27172
rect 24078 27228 24142 27232
rect 24078 27172 24082 27228
rect 24082 27172 24138 27228
rect 24138 27172 24142 27228
rect 24078 27168 24142 27172
rect 24158 27228 24222 27232
rect 24158 27172 24162 27228
rect 24162 27172 24218 27228
rect 24218 27172 24222 27228
rect 24158 27168 24222 27172
rect 24238 27228 24302 27232
rect 24238 27172 24242 27228
rect 24242 27172 24298 27228
rect 24298 27172 24302 27228
rect 24238 27168 24302 27172
rect 31680 27228 31744 27232
rect 31680 27172 31684 27228
rect 31684 27172 31740 27228
rect 31740 27172 31744 27228
rect 31680 27168 31744 27172
rect 31760 27228 31824 27232
rect 31760 27172 31764 27228
rect 31764 27172 31820 27228
rect 31820 27172 31824 27228
rect 31760 27168 31824 27172
rect 31840 27228 31904 27232
rect 31840 27172 31844 27228
rect 31844 27172 31900 27228
rect 31900 27172 31904 27228
rect 31840 27168 31904 27172
rect 31920 27228 31984 27232
rect 31920 27172 31924 27228
rect 31924 27172 31980 27228
rect 31980 27172 31984 27228
rect 31920 27168 31984 27172
rect 25084 27160 25148 27164
rect 25084 27104 25134 27160
rect 25134 27104 25148 27160
rect 25084 27100 25148 27104
rect 27660 27100 27724 27164
rect 30236 27100 30300 27164
rect 17172 26828 17236 26892
rect 18460 26964 18524 27028
rect 23244 26964 23308 27028
rect 14228 26752 14292 26756
rect 14228 26696 14242 26752
rect 14242 26696 14292 26752
rect 14228 26692 14292 26696
rect 15148 26692 15212 26756
rect 17908 26692 17972 26756
rect 4793 26684 4857 26688
rect 4793 26628 4797 26684
rect 4797 26628 4853 26684
rect 4853 26628 4857 26684
rect 4793 26624 4857 26628
rect 4873 26684 4937 26688
rect 4873 26628 4877 26684
rect 4877 26628 4933 26684
rect 4933 26628 4937 26684
rect 4873 26624 4937 26628
rect 4953 26684 5017 26688
rect 4953 26628 4957 26684
rect 4957 26628 5013 26684
rect 5013 26628 5017 26684
rect 4953 26624 5017 26628
rect 5033 26684 5097 26688
rect 5033 26628 5037 26684
rect 5037 26628 5093 26684
rect 5093 26628 5097 26684
rect 5033 26624 5097 26628
rect 12475 26684 12539 26688
rect 12475 26628 12479 26684
rect 12479 26628 12535 26684
rect 12535 26628 12539 26684
rect 12475 26624 12539 26628
rect 12555 26684 12619 26688
rect 12555 26628 12559 26684
rect 12559 26628 12615 26684
rect 12615 26628 12619 26684
rect 12555 26624 12619 26628
rect 12635 26684 12699 26688
rect 12635 26628 12639 26684
rect 12639 26628 12695 26684
rect 12695 26628 12699 26684
rect 12635 26624 12699 26628
rect 12715 26684 12779 26688
rect 12715 26628 12719 26684
rect 12719 26628 12775 26684
rect 12775 26628 12779 26684
rect 12715 26624 12779 26628
rect 20668 26692 20732 26756
rect 24900 26828 24964 26892
rect 26740 26888 26804 26892
rect 26740 26832 26754 26888
rect 26754 26832 26804 26888
rect 26740 26828 26804 26832
rect 29684 26828 29748 26892
rect 30420 26964 30484 27028
rect 20157 26684 20221 26688
rect 20157 26628 20161 26684
rect 20161 26628 20217 26684
rect 20217 26628 20221 26684
rect 20157 26624 20221 26628
rect 20237 26684 20301 26688
rect 20237 26628 20241 26684
rect 20241 26628 20297 26684
rect 20297 26628 20301 26684
rect 20237 26624 20301 26628
rect 20317 26684 20381 26688
rect 20317 26628 20321 26684
rect 20321 26628 20377 26684
rect 20377 26628 20381 26684
rect 20317 26624 20381 26628
rect 20397 26684 20461 26688
rect 20397 26628 20401 26684
rect 20401 26628 20457 26684
rect 20457 26628 20461 26684
rect 20397 26624 20461 26628
rect 14780 26420 14844 26484
rect 15332 26420 15396 26484
rect 16804 26420 16868 26484
rect 17908 26480 17972 26484
rect 17908 26424 17958 26480
rect 17958 26424 17972 26480
rect 14964 26284 15028 26348
rect 15700 26284 15764 26348
rect 16804 26284 16868 26348
rect 17908 26420 17972 26424
rect 18092 26480 18156 26484
rect 18092 26424 18142 26480
rect 18142 26424 18156 26480
rect 18092 26420 18156 26424
rect 19380 26616 19444 26620
rect 19380 26560 19430 26616
rect 19430 26560 19444 26616
rect 19380 26556 19444 26560
rect 19932 26556 19996 26620
rect 21772 26556 21836 26620
rect 18644 26420 18708 26484
rect 18092 26284 18156 26348
rect 20668 26420 20732 26484
rect 13676 26148 13740 26212
rect 20852 26284 20916 26348
rect 27839 26684 27903 26688
rect 27839 26628 27843 26684
rect 27843 26628 27899 26684
rect 27899 26628 27903 26684
rect 27839 26624 27903 26628
rect 27919 26684 27983 26688
rect 27919 26628 27923 26684
rect 27923 26628 27979 26684
rect 27979 26628 27983 26684
rect 27919 26624 27983 26628
rect 27999 26684 28063 26688
rect 27999 26628 28003 26684
rect 28003 26628 28059 26684
rect 28059 26628 28063 26684
rect 27999 26624 28063 26628
rect 28079 26684 28143 26688
rect 28079 26628 28083 26684
rect 28083 26628 28139 26684
rect 28139 26628 28143 26684
rect 28079 26624 28143 26628
rect 23796 26616 23860 26620
rect 23796 26560 23846 26616
rect 23846 26560 23860 26616
rect 23796 26556 23860 26560
rect 24716 26556 24780 26620
rect 26740 26556 26804 26620
rect 27660 26556 27724 26620
rect 8634 26140 8698 26144
rect 8634 26084 8638 26140
rect 8638 26084 8694 26140
rect 8694 26084 8698 26140
rect 8634 26080 8698 26084
rect 8714 26140 8778 26144
rect 8714 26084 8718 26140
rect 8718 26084 8774 26140
rect 8774 26084 8778 26140
rect 8714 26080 8778 26084
rect 8794 26140 8858 26144
rect 8794 26084 8798 26140
rect 8798 26084 8854 26140
rect 8854 26084 8858 26140
rect 8794 26080 8858 26084
rect 8874 26140 8938 26144
rect 8874 26084 8878 26140
rect 8878 26084 8934 26140
rect 8934 26084 8938 26140
rect 8874 26080 8938 26084
rect 16316 26140 16380 26144
rect 16316 26084 16320 26140
rect 16320 26084 16376 26140
rect 16376 26084 16380 26140
rect 16316 26080 16380 26084
rect 16396 26140 16460 26144
rect 16396 26084 16400 26140
rect 16400 26084 16456 26140
rect 16456 26084 16460 26140
rect 16396 26080 16460 26084
rect 16476 26140 16540 26144
rect 16476 26084 16480 26140
rect 16480 26084 16536 26140
rect 16536 26084 16540 26140
rect 16476 26080 16540 26084
rect 16556 26140 16620 26144
rect 16556 26084 16560 26140
rect 16560 26084 16616 26140
rect 16616 26084 16620 26140
rect 16556 26080 16620 26084
rect 13492 26012 13556 26076
rect 14044 26012 14108 26076
rect 17172 26012 17236 26076
rect 14596 25876 14660 25940
rect 18092 26012 18156 26076
rect 20852 26148 20916 26212
rect 19932 25876 19996 25940
rect 20668 26012 20732 26076
rect 28764 26556 28828 26620
rect 29500 26556 29564 26620
rect 30052 26556 30116 26620
rect 28396 26420 28460 26484
rect 29500 26420 29564 26484
rect 30604 26556 30668 26620
rect 30420 26420 30484 26484
rect 21220 26208 21284 26212
rect 21220 26152 21234 26208
rect 21234 26152 21284 26208
rect 21220 26148 21284 26152
rect 24716 26284 24780 26348
rect 24900 26284 24964 26348
rect 25452 26284 25516 26348
rect 27292 26284 27356 26348
rect 28212 26284 28276 26348
rect 28764 26344 28828 26348
rect 28764 26288 28778 26344
rect 28778 26288 28828 26344
rect 28764 26284 28828 26288
rect 29684 26284 29748 26348
rect 23060 26148 23124 26212
rect 23796 26148 23860 26212
rect 23998 26140 24062 26144
rect 23998 26084 24002 26140
rect 24002 26084 24058 26140
rect 24058 26084 24062 26140
rect 23998 26080 24062 26084
rect 24078 26140 24142 26144
rect 24078 26084 24082 26140
rect 24082 26084 24138 26140
rect 24138 26084 24142 26140
rect 24078 26080 24142 26084
rect 24158 26140 24222 26144
rect 24158 26084 24162 26140
rect 24162 26084 24218 26140
rect 24218 26084 24222 26140
rect 24158 26080 24222 26084
rect 24238 26140 24302 26144
rect 24238 26084 24242 26140
rect 24242 26084 24298 26140
rect 24298 26084 24302 26140
rect 24238 26080 24302 26084
rect 31680 26140 31744 26144
rect 31680 26084 31684 26140
rect 31684 26084 31740 26140
rect 31740 26084 31744 26140
rect 31680 26080 31744 26084
rect 31760 26140 31824 26144
rect 31760 26084 31764 26140
rect 31764 26084 31820 26140
rect 31820 26084 31824 26140
rect 31760 26080 31824 26084
rect 31840 26140 31904 26144
rect 31840 26084 31844 26140
rect 31844 26084 31900 26140
rect 31900 26084 31904 26140
rect 31840 26080 31904 26084
rect 31920 26140 31984 26144
rect 31920 26084 31924 26140
rect 31924 26084 31980 26140
rect 31980 26084 31984 26140
rect 31920 26080 31984 26084
rect 21220 25936 21284 25940
rect 21220 25880 21270 25936
rect 21270 25880 21284 25936
rect 21220 25876 21284 25880
rect 23060 26012 23124 26076
rect 24900 26012 24964 26076
rect 28396 26012 28460 26076
rect 24394 25876 24458 25940
rect 26004 25876 26068 25940
rect 30788 26012 30852 26076
rect 17540 25604 17604 25668
rect 19196 25604 19260 25668
rect 25084 25740 25148 25804
rect 27660 25740 27724 25804
rect 29868 25876 29932 25940
rect 27660 25604 27724 25668
rect 29132 25604 29196 25668
rect 4793 25596 4857 25600
rect 4793 25540 4797 25596
rect 4797 25540 4853 25596
rect 4853 25540 4857 25596
rect 4793 25536 4857 25540
rect 4873 25596 4937 25600
rect 4873 25540 4877 25596
rect 4877 25540 4933 25596
rect 4933 25540 4937 25596
rect 4873 25536 4937 25540
rect 4953 25596 5017 25600
rect 4953 25540 4957 25596
rect 4957 25540 5013 25596
rect 5013 25540 5017 25596
rect 4953 25536 5017 25540
rect 5033 25596 5097 25600
rect 5033 25540 5037 25596
rect 5037 25540 5093 25596
rect 5093 25540 5097 25596
rect 5033 25536 5097 25540
rect 12475 25596 12539 25600
rect 12475 25540 12479 25596
rect 12479 25540 12535 25596
rect 12535 25540 12539 25596
rect 12475 25536 12539 25540
rect 12555 25596 12619 25600
rect 12555 25540 12559 25596
rect 12559 25540 12615 25596
rect 12615 25540 12619 25596
rect 12555 25536 12619 25540
rect 12635 25596 12699 25600
rect 12635 25540 12639 25596
rect 12639 25540 12695 25596
rect 12695 25540 12699 25596
rect 12635 25536 12699 25540
rect 12715 25596 12779 25600
rect 12715 25540 12719 25596
rect 12719 25540 12775 25596
rect 12775 25540 12779 25596
rect 12715 25536 12779 25540
rect 20157 25596 20221 25600
rect 20157 25540 20161 25596
rect 20161 25540 20217 25596
rect 20217 25540 20221 25596
rect 20157 25536 20221 25540
rect 20237 25596 20301 25600
rect 20237 25540 20241 25596
rect 20241 25540 20297 25596
rect 20297 25540 20301 25596
rect 20237 25536 20301 25540
rect 20317 25596 20381 25600
rect 20317 25540 20321 25596
rect 20321 25540 20377 25596
rect 20377 25540 20381 25596
rect 20317 25536 20381 25540
rect 20397 25596 20461 25600
rect 20397 25540 20401 25596
rect 20401 25540 20457 25596
rect 20457 25540 20461 25596
rect 20397 25536 20461 25540
rect 30604 25604 30668 25668
rect 27839 25596 27903 25600
rect 27839 25540 27843 25596
rect 27843 25540 27899 25596
rect 27899 25540 27903 25596
rect 27839 25536 27903 25540
rect 27919 25596 27983 25600
rect 27919 25540 27923 25596
rect 27923 25540 27979 25596
rect 27979 25540 27983 25596
rect 27919 25536 27983 25540
rect 27999 25596 28063 25600
rect 27999 25540 28003 25596
rect 28003 25540 28059 25596
rect 28059 25540 28063 25596
rect 27999 25536 28063 25540
rect 28079 25596 28143 25600
rect 28079 25540 28083 25596
rect 28083 25540 28139 25596
rect 28139 25540 28143 25596
rect 28079 25536 28143 25540
rect 5396 25468 5460 25532
rect 12020 25468 12084 25532
rect 14228 25528 14292 25532
rect 14228 25472 14278 25528
rect 14278 25472 14292 25528
rect 14228 25468 14292 25472
rect 14596 25468 14660 25532
rect 17356 25468 17420 25532
rect 19564 25392 19628 25396
rect 20668 25468 20732 25532
rect 25268 25468 25332 25532
rect 29132 25468 29196 25532
rect 32076 25468 32140 25532
rect 19564 25336 19578 25392
rect 19578 25336 19628 25392
rect 19564 25332 19628 25336
rect 23612 25392 23676 25396
rect 23612 25336 23662 25392
rect 23662 25336 23676 25392
rect 23612 25332 23676 25336
rect 24532 25332 24596 25396
rect 31156 25332 31220 25396
rect 32444 25392 32508 25396
rect 32444 25336 32494 25392
rect 32494 25336 32508 25392
rect 32444 25332 32508 25336
rect 14596 25196 14660 25260
rect 14780 25196 14844 25260
rect 8634 25052 8698 25056
rect 8634 24996 8638 25052
rect 8638 24996 8694 25052
rect 8694 24996 8698 25052
rect 8634 24992 8698 24996
rect 8714 25052 8778 25056
rect 8714 24996 8718 25052
rect 8718 24996 8774 25052
rect 8774 24996 8778 25052
rect 8714 24992 8778 24996
rect 8794 25052 8858 25056
rect 8794 24996 8798 25052
rect 8798 24996 8854 25052
rect 8854 24996 8858 25052
rect 8794 24992 8858 24996
rect 8874 25052 8938 25056
rect 8874 24996 8878 25052
rect 8878 24996 8934 25052
rect 8934 24996 8938 25052
rect 8874 24992 8938 24996
rect 17540 25060 17604 25124
rect 20668 25060 20732 25124
rect 16316 25052 16380 25056
rect 16316 24996 16320 25052
rect 16320 24996 16376 25052
rect 16376 24996 16380 25052
rect 16316 24992 16380 24996
rect 16396 25052 16460 25056
rect 16396 24996 16400 25052
rect 16400 24996 16456 25052
rect 16456 24996 16460 25052
rect 16396 24992 16460 24996
rect 16476 25052 16540 25056
rect 16476 24996 16480 25052
rect 16480 24996 16536 25052
rect 16536 24996 16540 25052
rect 16476 24992 16540 24996
rect 16556 25052 16620 25056
rect 16556 24996 16560 25052
rect 16560 24996 16616 25052
rect 16616 24996 16620 25052
rect 16556 24992 16620 24996
rect 25268 25196 25332 25260
rect 30604 25196 30668 25260
rect 32628 25196 32692 25260
rect 15884 24924 15948 24988
rect 18644 24924 18708 24988
rect 20530 24924 20594 24988
rect 21404 24924 21468 24988
rect 21772 24924 21836 24988
rect 22692 24924 22756 24988
rect 15516 24788 15580 24852
rect 26556 25060 26620 25124
rect 23998 25052 24062 25056
rect 23998 24996 24002 25052
rect 24002 24996 24058 25052
rect 24058 24996 24062 25052
rect 23998 24992 24062 24996
rect 24078 25052 24142 25056
rect 24078 24996 24082 25052
rect 24082 24996 24138 25052
rect 24138 24996 24142 25052
rect 24078 24992 24142 24996
rect 24158 25052 24222 25056
rect 24158 24996 24162 25052
rect 24162 24996 24218 25052
rect 24218 24996 24222 25052
rect 24158 24992 24222 24996
rect 24238 25052 24302 25056
rect 24238 24996 24242 25052
rect 24242 24996 24298 25052
rect 24298 24996 24302 25052
rect 24238 24992 24302 24996
rect 31680 25052 31744 25056
rect 31680 24996 31684 25052
rect 31684 24996 31740 25052
rect 31740 24996 31744 25052
rect 31680 24992 31744 24996
rect 31760 25052 31824 25056
rect 31760 24996 31764 25052
rect 31764 24996 31820 25052
rect 31820 24996 31824 25052
rect 31760 24992 31824 24996
rect 31840 25052 31904 25056
rect 31840 24996 31844 25052
rect 31844 24996 31900 25052
rect 31900 24996 31904 25052
rect 31840 24992 31904 24996
rect 31920 25052 31984 25056
rect 31920 24996 31924 25052
rect 31924 24996 31980 25052
rect 31980 24996 31984 25052
rect 31920 24992 31984 24996
rect 23612 24984 23676 24988
rect 23612 24928 23626 24984
rect 23626 24928 23676 24984
rect 23612 24924 23676 24928
rect 25084 24924 25148 24988
rect 29868 24924 29932 24988
rect 31156 24984 31220 24988
rect 31156 24928 31170 24984
rect 31170 24928 31220 24984
rect 31156 24924 31220 24928
rect 6868 24652 6932 24716
rect 14780 24652 14844 24716
rect 15516 24652 15580 24716
rect 16068 24652 16132 24716
rect 17356 24652 17420 24716
rect 26372 24788 26436 24852
rect 26740 24788 26804 24852
rect 29132 24848 29196 24852
rect 29132 24792 29146 24848
rect 29146 24792 29196 24848
rect 29132 24788 29196 24792
rect 13860 24516 13924 24580
rect 15332 24576 15396 24580
rect 15332 24520 15382 24576
rect 15382 24520 15396 24576
rect 15332 24516 15396 24520
rect 4793 24508 4857 24512
rect 4793 24452 4797 24508
rect 4797 24452 4853 24508
rect 4853 24452 4857 24508
rect 4793 24448 4857 24452
rect 4873 24508 4937 24512
rect 4873 24452 4877 24508
rect 4877 24452 4933 24508
rect 4933 24452 4937 24508
rect 4873 24448 4937 24452
rect 4953 24508 5017 24512
rect 4953 24452 4957 24508
rect 4957 24452 5013 24508
rect 5013 24452 5017 24508
rect 4953 24448 5017 24452
rect 5033 24508 5097 24512
rect 5033 24452 5037 24508
rect 5037 24452 5093 24508
rect 5093 24452 5097 24508
rect 5033 24448 5097 24452
rect 12475 24508 12539 24512
rect 12475 24452 12479 24508
rect 12479 24452 12535 24508
rect 12535 24452 12539 24508
rect 12475 24448 12539 24452
rect 12555 24508 12619 24512
rect 12555 24452 12559 24508
rect 12559 24452 12615 24508
rect 12615 24452 12619 24508
rect 12555 24448 12619 24452
rect 12635 24508 12699 24512
rect 12635 24452 12639 24508
rect 12639 24452 12695 24508
rect 12695 24452 12699 24508
rect 12635 24448 12699 24452
rect 12715 24508 12779 24512
rect 12715 24452 12719 24508
rect 12719 24452 12775 24508
rect 12775 24452 12779 24508
rect 12715 24448 12779 24452
rect 20157 24508 20221 24512
rect 20157 24452 20161 24508
rect 20161 24452 20217 24508
rect 20217 24452 20221 24508
rect 20157 24448 20221 24452
rect 20237 24508 20301 24512
rect 20237 24452 20241 24508
rect 20241 24452 20297 24508
rect 20297 24452 20301 24508
rect 20237 24448 20301 24452
rect 20317 24508 20381 24512
rect 20317 24452 20321 24508
rect 20321 24452 20377 24508
rect 20377 24452 20381 24508
rect 20317 24448 20381 24452
rect 20397 24508 20461 24512
rect 20397 24452 20401 24508
rect 20401 24452 20457 24508
rect 20457 24452 20461 24508
rect 20397 24448 20461 24452
rect 14044 24380 14108 24444
rect 16804 24380 16868 24444
rect 19012 24380 19076 24444
rect 7052 24244 7116 24308
rect 15332 24244 15396 24308
rect 19564 24440 19628 24444
rect 19564 24384 19578 24440
rect 19578 24384 19628 24440
rect 19564 24380 19628 24384
rect 21404 24380 21468 24444
rect 21588 24440 21652 24444
rect 21588 24384 21602 24440
rect 21602 24384 21652 24440
rect 21588 24380 21652 24384
rect 22876 24244 22940 24308
rect 25820 24440 25884 24444
rect 27108 24516 27172 24580
rect 32260 24652 32324 24716
rect 27839 24508 27903 24512
rect 27839 24452 27843 24508
rect 27843 24452 27899 24508
rect 27899 24452 27903 24508
rect 27839 24448 27903 24452
rect 27919 24508 27983 24512
rect 27919 24452 27923 24508
rect 27923 24452 27979 24508
rect 27979 24452 27983 24508
rect 27919 24448 27983 24452
rect 27999 24508 28063 24512
rect 27999 24452 28003 24508
rect 28003 24452 28059 24508
rect 28059 24452 28063 24508
rect 27999 24448 28063 24452
rect 28079 24508 28143 24512
rect 28079 24452 28083 24508
rect 28083 24452 28139 24508
rect 28139 24452 28143 24508
rect 28079 24448 28143 24452
rect 25820 24384 25870 24440
rect 25870 24384 25884 24440
rect 25820 24380 25884 24384
rect 29868 24380 29932 24444
rect 13860 24168 13924 24172
rect 13860 24112 13910 24168
rect 13910 24112 13924 24168
rect 13860 24108 13924 24112
rect 8634 23964 8698 23968
rect 8634 23908 8638 23964
rect 8638 23908 8694 23964
rect 8694 23908 8698 23964
rect 8634 23904 8698 23908
rect 8714 23964 8778 23968
rect 8714 23908 8718 23964
rect 8718 23908 8774 23964
rect 8774 23908 8778 23964
rect 8714 23904 8778 23908
rect 8794 23964 8858 23968
rect 8794 23908 8798 23964
rect 8798 23908 8854 23964
rect 8854 23908 8858 23964
rect 8794 23904 8858 23908
rect 8874 23964 8938 23968
rect 8874 23908 8878 23964
rect 8878 23908 8934 23964
rect 8934 23908 8938 23964
rect 8874 23904 8938 23908
rect 15148 23972 15212 24036
rect 16804 24032 16868 24036
rect 16804 23976 16818 24032
rect 16818 23976 16868 24032
rect 16804 23972 16868 23976
rect 17540 23972 17604 24036
rect 21772 24108 21836 24172
rect 22692 24108 22756 24172
rect 30052 24244 30116 24308
rect 27476 23972 27540 24036
rect 16316 23964 16380 23968
rect 16316 23908 16320 23964
rect 16320 23908 16376 23964
rect 16376 23908 16380 23964
rect 16316 23904 16380 23908
rect 16396 23964 16460 23968
rect 16396 23908 16400 23964
rect 16400 23908 16456 23964
rect 16456 23908 16460 23964
rect 16396 23904 16460 23908
rect 16476 23964 16540 23968
rect 16476 23908 16480 23964
rect 16480 23908 16536 23964
rect 16536 23908 16540 23964
rect 16476 23904 16540 23908
rect 16556 23964 16620 23968
rect 16556 23908 16560 23964
rect 16560 23908 16616 23964
rect 16616 23908 16620 23964
rect 16556 23904 16620 23908
rect 23998 23964 24062 23968
rect 23998 23908 24002 23964
rect 24002 23908 24058 23964
rect 24058 23908 24062 23964
rect 23998 23904 24062 23908
rect 24078 23964 24142 23968
rect 24078 23908 24082 23964
rect 24082 23908 24138 23964
rect 24138 23908 24142 23964
rect 24078 23904 24142 23908
rect 24158 23964 24222 23968
rect 24158 23908 24162 23964
rect 24162 23908 24218 23964
rect 24218 23908 24222 23964
rect 24158 23904 24222 23908
rect 24238 23964 24302 23968
rect 24238 23908 24242 23964
rect 24242 23908 24298 23964
rect 24298 23908 24302 23964
rect 24238 23904 24302 23908
rect 31680 23964 31744 23968
rect 31680 23908 31684 23964
rect 31684 23908 31740 23964
rect 31740 23908 31744 23964
rect 31680 23904 31744 23908
rect 31760 23964 31824 23968
rect 31760 23908 31764 23964
rect 31764 23908 31820 23964
rect 31820 23908 31824 23964
rect 31760 23904 31824 23908
rect 31840 23964 31904 23968
rect 31840 23908 31844 23964
rect 31844 23908 31900 23964
rect 31900 23908 31904 23964
rect 31840 23904 31904 23908
rect 31920 23964 31984 23968
rect 31920 23908 31924 23964
rect 31924 23908 31980 23964
rect 31980 23908 31984 23964
rect 31920 23904 31984 23908
rect 17172 23836 17236 23900
rect 17540 23896 17604 23900
rect 17540 23840 17590 23896
rect 17590 23840 17604 23896
rect 17540 23836 17604 23840
rect 17724 23836 17788 23900
rect 14596 23700 14660 23764
rect 23796 23896 23860 23900
rect 23796 23840 23810 23896
rect 23810 23840 23860 23896
rect 23796 23836 23860 23840
rect 22508 23700 22572 23764
rect 26740 23760 26804 23764
rect 26740 23704 26754 23760
rect 26754 23704 26804 23760
rect 26740 23700 26804 23704
rect 6316 23428 6380 23492
rect 13492 23428 13556 23492
rect 15516 23564 15580 23628
rect 4793 23420 4857 23424
rect 4793 23364 4797 23420
rect 4797 23364 4853 23420
rect 4853 23364 4857 23420
rect 4793 23360 4857 23364
rect 4873 23420 4937 23424
rect 4873 23364 4877 23420
rect 4877 23364 4933 23420
rect 4933 23364 4937 23420
rect 4873 23360 4937 23364
rect 4953 23420 5017 23424
rect 4953 23364 4957 23420
rect 4957 23364 5013 23420
rect 5013 23364 5017 23420
rect 4953 23360 5017 23364
rect 5033 23420 5097 23424
rect 5033 23364 5037 23420
rect 5037 23364 5093 23420
rect 5093 23364 5097 23420
rect 5033 23360 5097 23364
rect 12475 23420 12539 23424
rect 12475 23364 12479 23420
rect 12479 23364 12535 23420
rect 12535 23364 12539 23420
rect 12475 23360 12539 23364
rect 12555 23420 12619 23424
rect 12555 23364 12559 23420
rect 12559 23364 12615 23420
rect 12615 23364 12619 23420
rect 12555 23360 12619 23364
rect 12635 23420 12699 23424
rect 12635 23364 12639 23420
rect 12639 23364 12695 23420
rect 12695 23364 12699 23420
rect 12635 23360 12699 23364
rect 12715 23420 12779 23424
rect 12715 23364 12719 23420
rect 12719 23364 12775 23420
rect 12775 23364 12779 23420
rect 12715 23360 12779 23364
rect 9260 23292 9324 23356
rect 13308 23352 13372 23356
rect 13308 23296 13358 23352
rect 13358 23296 13372 23352
rect 13308 23292 13372 23296
rect 17540 23428 17604 23492
rect 14780 23352 14844 23356
rect 14780 23296 14830 23352
rect 14830 23296 14844 23352
rect 14780 23292 14844 23296
rect 15148 23292 15212 23356
rect 16988 23292 17052 23356
rect 19748 23428 19812 23492
rect 20668 23428 20732 23492
rect 20157 23420 20221 23424
rect 20157 23364 20161 23420
rect 20161 23364 20217 23420
rect 20217 23364 20221 23420
rect 20157 23360 20221 23364
rect 20237 23420 20301 23424
rect 20237 23364 20241 23420
rect 20241 23364 20297 23420
rect 20297 23364 20301 23420
rect 20237 23360 20301 23364
rect 20317 23420 20381 23424
rect 20317 23364 20321 23420
rect 20321 23364 20377 23420
rect 20377 23364 20381 23420
rect 20317 23360 20381 23364
rect 20397 23420 20461 23424
rect 20397 23364 20401 23420
rect 20401 23364 20457 23420
rect 20457 23364 20461 23420
rect 20397 23360 20461 23364
rect 20668 23292 20732 23356
rect 20852 23292 20916 23356
rect 27292 23564 27356 23628
rect 24532 23428 24596 23492
rect 26740 23428 26804 23492
rect 28396 23428 28460 23492
rect 27839 23420 27903 23424
rect 27839 23364 27843 23420
rect 27843 23364 27899 23420
rect 27899 23364 27903 23420
rect 27839 23360 27903 23364
rect 27919 23420 27983 23424
rect 27919 23364 27923 23420
rect 27923 23364 27979 23420
rect 27979 23364 27983 23420
rect 27919 23360 27983 23364
rect 27999 23420 28063 23424
rect 27999 23364 28003 23420
rect 28003 23364 28059 23420
rect 28059 23364 28063 23420
rect 27999 23360 28063 23364
rect 28079 23420 28143 23424
rect 28079 23364 28083 23420
rect 28083 23364 28139 23420
rect 28139 23364 28143 23420
rect 28079 23360 28143 23364
rect 27108 23292 27172 23356
rect 27660 23352 27724 23356
rect 27660 23296 27710 23352
rect 27710 23296 27724 23352
rect 27660 23292 27724 23296
rect 28396 23352 28460 23356
rect 28396 23296 28446 23352
rect 28446 23296 28460 23352
rect 28396 23292 28460 23296
rect 28764 23352 28828 23356
rect 28764 23296 28814 23352
rect 28814 23296 28828 23352
rect 28764 23292 28828 23296
rect 30236 23292 30300 23356
rect 31340 23292 31404 23356
rect 17908 23156 17972 23220
rect 13492 22884 13556 22948
rect 8634 22876 8698 22880
rect 8634 22820 8638 22876
rect 8638 22820 8694 22876
rect 8694 22820 8698 22876
rect 8634 22816 8698 22820
rect 8714 22876 8778 22880
rect 8714 22820 8718 22876
rect 8718 22820 8774 22876
rect 8774 22820 8778 22876
rect 8714 22816 8778 22820
rect 8794 22876 8858 22880
rect 8794 22820 8798 22876
rect 8798 22820 8854 22876
rect 8854 22820 8858 22876
rect 8794 22816 8858 22820
rect 8874 22876 8938 22880
rect 8874 22820 8878 22876
rect 8878 22820 8934 22876
rect 8934 22820 8938 22876
rect 8874 22816 8938 22820
rect 16316 22876 16380 22880
rect 16316 22820 16320 22876
rect 16320 22820 16376 22876
rect 16376 22820 16380 22876
rect 16316 22816 16380 22820
rect 16396 22876 16460 22880
rect 16396 22820 16400 22876
rect 16400 22820 16456 22876
rect 16456 22820 16460 22876
rect 16396 22816 16460 22820
rect 16476 22876 16540 22880
rect 16476 22820 16480 22876
rect 16480 22820 16536 22876
rect 16536 22820 16540 22876
rect 16476 22816 16540 22820
rect 16556 22876 16620 22880
rect 16556 22820 16560 22876
rect 16560 22820 16616 22876
rect 16616 22820 16620 22876
rect 16556 22816 16620 22820
rect 8156 22808 8220 22812
rect 8156 22752 8206 22808
rect 8206 22752 8220 22808
rect 8156 22748 8220 22752
rect 11468 22672 11532 22676
rect 11468 22616 11482 22672
rect 11482 22616 11532 22672
rect 11468 22612 11532 22616
rect 13860 22612 13924 22676
rect 17724 22944 17788 22948
rect 17724 22888 17774 22944
rect 17774 22888 17788 22944
rect 17724 22884 17788 22888
rect 18276 22884 18340 22948
rect 18644 22884 18708 22948
rect 23612 22884 23676 22948
rect 23998 22876 24062 22880
rect 23998 22820 24002 22876
rect 24002 22820 24058 22876
rect 24058 22820 24062 22876
rect 23998 22816 24062 22820
rect 24078 22876 24142 22880
rect 24078 22820 24082 22876
rect 24082 22820 24138 22876
rect 24138 22820 24142 22876
rect 24078 22816 24142 22820
rect 24158 22876 24222 22880
rect 24158 22820 24162 22876
rect 24162 22820 24218 22876
rect 24218 22820 24222 22876
rect 24158 22816 24222 22820
rect 24238 22876 24302 22880
rect 24238 22820 24242 22876
rect 24242 22820 24298 22876
rect 24298 22820 24302 22876
rect 24238 22816 24302 22820
rect 31680 22876 31744 22880
rect 31680 22820 31684 22876
rect 31684 22820 31740 22876
rect 31740 22820 31744 22876
rect 31680 22816 31744 22820
rect 31760 22876 31824 22880
rect 31760 22820 31764 22876
rect 31764 22820 31820 22876
rect 31820 22820 31824 22876
rect 31760 22816 31824 22820
rect 31840 22876 31904 22880
rect 31840 22820 31844 22876
rect 31844 22820 31900 22876
rect 31900 22820 31904 22876
rect 31840 22816 31904 22820
rect 31920 22876 31984 22880
rect 31920 22820 31924 22876
rect 31924 22820 31980 22876
rect 31980 22820 31984 22876
rect 31920 22816 31984 22820
rect 17172 22748 17236 22812
rect 16988 22612 17052 22676
rect 17724 22612 17788 22676
rect 23428 22748 23492 22812
rect 24716 22748 24780 22812
rect 29868 22748 29932 22812
rect 30236 22748 30300 22812
rect 21036 22612 21100 22676
rect 21404 22612 21468 22676
rect 18276 22476 18340 22540
rect 21036 22476 21100 22540
rect 21588 22476 21652 22540
rect 13308 22400 13372 22404
rect 13308 22344 13322 22400
rect 13322 22344 13372 22400
rect 13308 22340 13372 22344
rect 21956 22476 22020 22540
rect 26372 22476 26436 22540
rect 27476 22536 27540 22540
rect 27476 22480 27526 22536
rect 27526 22480 27540 22536
rect 27476 22476 27540 22480
rect 27660 22476 27724 22540
rect 22140 22340 22204 22404
rect 25084 22340 25148 22404
rect 4793 22332 4857 22336
rect 4793 22276 4797 22332
rect 4797 22276 4853 22332
rect 4853 22276 4857 22332
rect 4793 22272 4857 22276
rect 4873 22332 4937 22336
rect 4873 22276 4877 22332
rect 4877 22276 4933 22332
rect 4933 22276 4937 22332
rect 4873 22272 4937 22276
rect 4953 22332 5017 22336
rect 4953 22276 4957 22332
rect 4957 22276 5013 22332
rect 5013 22276 5017 22332
rect 4953 22272 5017 22276
rect 5033 22332 5097 22336
rect 5033 22276 5037 22332
rect 5037 22276 5093 22332
rect 5093 22276 5097 22332
rect 5033 22272 5097 22276
rect 12475 22332 12539 22336
rect 12475 22276 12479 22332
rect 12479 22276 12535 22332
rect 12535 22276 12539 22332
rect 12475 22272 12539 22276
rect 12555 22332 12619 22336
rect 12555 22276 12559 22332
rect 12559 22276 12615 22332
rect 12615 22276 12619 22332
rect 12555 22272 12619 22276
rect 12635 22332 12699 22336
rect 12635 22276 12639 22332
rect 12639 22276 12695 22332
rect 12695 22276 12699 22332
rect 12635 22272 12699 22276
rect 12715 22332 12779 22336
rect 12715 22276 12719 22332
rect 12719 22276 12775 22332
rect 12775 22276 12779 22332
rect 12715 22272 12779 22276
rect 20157 22332 20221 22336
rect 20157 22276 20161 22332
rect 20161 22276 20217 22332
rect 20217 22276 20221 22332
rect 20157 22272 20221 22276
rect 20237 22332 20301 22336
rect 20237 22276 20241 22332
rect 20241 22276 20297 22332
rect 20297 22276 20301 22332
rect 20237 22272 20301 22276
rect 20317 22332 20381 22336
rect 20317 22276 20321 22332
rect 20321 22276 20377 22332
rect 20377 22276 20381 22332
rect 20317 22272 20381 22276
rect 20397 22332 20461 22336
rect 20397 22276 20401 22332
rect 20401 22276 20457 22332
rect 20457 22276 20461 22332
rect 20397 22272 20461 22276
rect 27839 22332 27903 22336
rect 27839 22276 27843 22332
rect 27843 22276 27899 22332
rect 27899 22276 27903 22332
rect 27839 22272 27903 22276
rect 27919 22332 27983 22336
rect 27919 22276 27923 22332
rect 27923 22276 27979 22332
rect 27979 22276 27983 22332
rect 27919 22272 27983 22276
rect 27999 22332 28063 22336
rect 27999 22276 28003 22332
rect 28003 22276 28059 22332
rect 28059 22276 28063 22332
rect 27999 22272 28063 22276
rect 28079 22332 28143 22336
rect 28079 22276 28083 22332
rect 28083 22276 28139 22332
rect 28139 22276 28143 22332
rect 28079 22272 28143 22276
rect 12020 22264 12084 22268
rect 12020 22208 12034 22264
rect 12034 22208 12084 22264
rect 12020 22204 12084 22208
rect 13860 22204 13924 22268
rect 16804 22204 16868 22268
rect 18644 22204 18708 22268
rect 19380 22204 19444 22268
rect 20668 22204 20732 22268
rect 10180 21932 10244 21996
rect 6868 21796 6932 21860
rect 13124 21796 13188 21860
rect 15884 21796 15948 21860
rect 8634 21788 8698 21792
rect 8634 21732 8638 21788
rect 8638 21732 8694 21788
rect 8694 21732 8698 21788
rect 8634 21728 8698 21732
rect 8714 21788 8778 21792
rect 8714 21732 8718 21788
rect 8718 21732 8774 21788
rect 8774 21732 8778 21788
rect 8714 21728 8778 21732
rect 8794 21788 8858 21792
rect 8794 21732 8798 21788
rect 8798 21732 8854 21788
rect 8854 21732 8858 21788
rect 8794 21728 8858 21732
rect 8874 21788 8938 21792
rect 8874 21732 8878 21788
rect 8878 21732 8934 21788
rect 8934 21732 8938 21788
rect 8874 21728 8938 21732
rect 16316 21788 16380 21792
rect 16316 21732 16320 21788
rect 16320 21732 16376 21788
rect 16376 21732 16380 21788
rect 16316 21728 16380 21732
rect 16396 21788 16460 21792
rect 16396 21732 16400 21788
rect 16400 21732 16456 21788
rect 16456 21732 16460 21788
rect 16396 21728 16460 21732
rect 16476 21788 16540 21792
rect 16476 21732 16480 21788
rect 16480 21732 16536 21788
rect 16536 21732 16540 21788
rect 16476 21728 16540 21732
rect 16556 21788 16620 21792
rect 16556 21732 16560 21788
rect 16560 21732 16616 21788
rect 16616 21732 16620 21788
rect 16556 21728 16620 21732
rect 12204 21720 12268 21724
rect 12204 21664 12254 21720
rect 12254 21664 12268 21720
rect 12204 21660 12268 21664
rect 14228 21720 14292 21724
rect 14228 21664 14242 21720
rect 14242 21664 14292 21720
rect 14228 21660 14292 21664
rect 18644 22068 18708 22132
rect 25636 22068 25700 22132
rect 26188 22128 26252 22132
rect 26188 22072 26202 22128
rect 26202 22072 26252 22128
rect 26188 22068 26252 22072
rect 26372 22068 26436 22132
rect 28396 22264 28460 22268
rect 28396 22208 28410 22264
rect 28410 22208 28460 22264
rect 28396 22204 28460 22208
rect 28948 22204 29012 22268
rect 17908 21992 17972 21996
rect 17908 21936 17958 21992
rect 17958 21936 17972 21992
rect 17908 21932 17972 21936
rect 17724 21796 17788 21860
rect 30972 21932 31036 21996
rect 18828 21796 18892 21860
rect 21772 21796 21836 21860
rect 22692 21796 22756 21860
rect 26556 21796 26620 21860
rect 23998 21788 24062 21792
rect 23998 21732 24002 21788
rect 24002 21732 24058 21788
rect 24058 21732 24062 21788
rect 23998 21728 24062 21732
rect 24078 21788 24142 21792
rect 24078 21732 24082 21788
rect 24082 21732 24138 21788
rect 24138 21732 24142 21788
rect 24078 21728 24142 21732
rect 24158 21788 24222 21792
rect 24158 21732 24162 21788
rect 24162 21732 24218 21788
rect 24218 21732 24222 21788
rect 24158 21728 24222 21732
rect 24238 21788 24302 21792
rect 24238 21732 24242 21788
rect 24242 21732 24298 21788
rect 24298 21732 24302 21788
rect 24238 21728 24302 21732
rect 17356 21660 17420 21724
rect 18092 21660 18156 21724
rect 18460 21720 18524 21724
rect 18460 21664 18510 21720
rect 18510 21664 18524 21720
rect 18460 21660 18524 21664
rect 19380 21660 19444 21724
rect 29132 21796 29196 21860
rect 30972 21796 31036 21860
rect 31680 21788 31744 21792
rect 31680 21732 31684 21788
rect 31684 21732 31740 21788
rect 31740 21732 31744 21788
rect 31680 21728 31744 21732
rect 31760 21788 31824 21792
rect 31760 21732 31764 21788
rect 31764 21732 31820 21788
rect 31820 21732 31824 21788
rect 31760 21728 31824 21732
rect 31840 21788 31904 21792
rect 31840 21732 31844 21788
rect 31844 21732 31900 21788
rect 31900 21732 31904 21788
rect 31840 21728 31904 21732
rect 31920 21788 31984 21792
rect 31920 21732 31924 21788
rect 31924 21732 31980 21788
rect 31980 21732 31984 21788
rect 31920 21728 31984 21732
rect 30420 21660 30484 21724
rect 31156 21660 31220 21724
rect 17172 21524 17236 21588
rect 17540 21524 17604 21588
rect 12940 21388 13004 21452
rect 17540 21388 17604 21452
rect 30604 21388 30668 21452
rect 30788 21448 30852 21452
rect 30788 21392 30838 21448
rect 30838 21392 30852 21448
rect 30788 21388 30852 21392
rect 13308 21252 13372 21316
rect 26556 21252 26620 21316
rect 4793 21244 4857 21248
rect 4793 21188 4797 21244
rect 4797 21188 4853 21244
rect 4853 21188 4857 21244
rect 4793 21184 4857 21188
rect 4873 21244 4937 21248
rect 4873 21188 4877 21244
rect 4877 21188 4933 21244
rect 4933 21188 4937 21244
rect 4873 21184 4937 21188
rect 4953 21244 5017 21248
rect 4953 21188 4957 21244
rect 4957 21188 5013 21244
rect 5013 21188 5017 21244
rect 4953 21184 5017 21188
rect 5033 21244 5097 21248
rect 5033 21188 5037 21244
rect 5037 21188 5093 21244
rect 5093 21188 5097 21244
rect 5033 21184 5097 21188
rect 12475 21244 12539 21248
rect 12475 21188 12479 21244
rect 12479 21188 12535 21244
rect 12535 21188 12539 21244
rect 12475 21184 12539 21188
rect 12555 21244 12619 21248
rect 12555 21188 12559 21244
rect 12559 21188 12615 21244
rect 12615 21188 12619 21244
rect 12555 21184 12619 21188
rect 12635 21244 12699 21248
rect 12635 21188 12639 21244
rect 12639 21188 12695 21244
rect 12695 21188 12699 21244
rect 12635 21184 12699 21188
rect 12715 21244 12779 21248
rect 12715 21188 12719 21244
rect 12719 21188 12775 21244
rect 12775 21188 12779 21244
rect 12715 21184 12779 21188
rect 20157 21244 20221 21248
rect 20157 21188 20161 21244
rect 20161 21188 20217 21244
rect 20217 21188 20221 21244
rect 20157 21184 20221 21188
rect 20237 21244 20301 21248
rect 20237 21188 20241 21244
rect 20241 21188 20297 21244
rect 20297 21188 20301 21244
rect 20237 21184 20301 21188
rect 20317 21244 20381 21248
rect 20317 21188 20321 21244
rect 20321 21188 20377 21244
rect 20377 21188 20381 21244
rect 20317 21184 20381 21188
rect 20397 21244 20461 21248
rect 20397 21188 20401 21244
rect 20401 21188 20457 21244
rect 20457 21188 20461 21244
rect 20397 21184 20461 21188
rect 27839 21244 27903 21248
rect 27839 21188 27843 21244
rect 27843 21188 27899 21244
rect 27899 21188 27903 21244
rect 27839 21184 27903 21188
rect 27919 21244 27983 21248
rect 27919 21188 27923 21244
rect 27923 21188 27979 21244
rect 27979 21188 27983 21244
rect 27919 21184 27983 21188
rect 27999 21244 28063 21248
rect 27999 21188 28003 21244
rect 28003 21188 28059 21244
rect 28059 21188 28063 21244
rect 27999 21184 28063 21188
rect 28079 21244 28143 21248
rect 28079 21188 28083 21244
rect 28083 21188 28139 21244
rect 28139 21188 28143 21244
rect 28079 21184 28143 21188
rect 12020 21116 12084 21180
rect 16988 21116 17052 21180
rect 19564 21116 19628 21180
rect 20668 21116 20732 21180
rect 22324 21116 22388 21180
rect 10916 20768 10980 20772
rect 10916 20712 10930 20768
rect 10930 20712 10980 20768
rect 10916 20708 10980 20712
rect 11652 20708 11716 20772
rect 12204 20708 12268 20772
rect 26924 20980 26988 21044
rect 27476 21040 27540 21044
rect 27476 20984 27490 21040
rect 27490 20984 27540 21040
rect 27476 20980 27540 20984
rect 28396 21116 28460 21180
rect 30052 20980 30116 21044
rect 17540 20844 17604 20908
rect 29684 20844 29748 20908
rect 30420 20844 30484 20908
rect 17172 20708 17236 20772
rect 25084 20708 25148 20772
rect 29684 20768 29748 20772
rect 29684 20712 29698 20768
rect 29698 20712 29748 20768
rect 29684 20708 29748 20712
rect 31156 20708 31220 20772
rect 8634 20700 8698 20704
rect 8634 20644 8638 20700
rect 8638 20644 8694 20700
rect 8694 20644 8698 20700
rect 8634 20640 8698 20644
rect 8714 20700 8778 20704
rect 8714 20644 8718 20700
rect 8718 20644 8774 20700
rect 8774 20644 8778 20700
rect 8714 20640 8778 20644
rect 8794 20700 8858 20704
rect 8794 20644 8798 20700
rect 8798 20644 8854 20700
rect 8854 20644 8858 20700
rect 8794 20640 8858 20644
rect 8874 20700 8938 20704
rect 8874 20644 8878 20700
rect 8878 20644 8934 20700
rect 8934 20644 8938 20700
rect 8874 20640 8938 20644
rect 16316 20700 16380 20704
rect 16316 20644 16320 20700
rect 16320 20644 16376 20700
rect 16376 20644 16380 20700
rect 16316 20640 16380 20644
rect 16396 20700 16460 20704
rect 16396 20644 16400 20700
rect 16400 20644 16456 20700
rect 16456 20644 16460 20700
rect 16396 20640 16460 20644
rect 16476 20700 16540 20704
rect 16476 20644 16480 20700
rect 16480 20644 16536 20700
rect 16536 20644 16540 20700
rect 16476 20640 16540 20644
rect 16556 20700 16620 20704
rect 16556 20644 16560 20700
rect 16560 20644 16616 20700
rect 16616 20644 16620 20700
rect 16556 20640 16620 20644
rect 23998 20700 24062 20704
rect 23998 20644 24002 20700
rect 24002 20644 24058 20700
rect 24058 20644 24062 20700
rect 23998 20640 24062 20644
rect 24078 20700 24142 20704
rect 24078 20644 24082 20700
rect 24082 20644 24138 20700
rect 24138 20644 24142 20700
rect 24078 20640 24142 20644
rect 24158 20700 24222 20704
rect 24158 20644 24162 20700
rect 24162 20644 24218 20700
rect 24218 20644 24222 20700
rect 24158 20640 24222 20644
rect 24238 20700 24302 20704
rect 24238 20644 24242 20700
rect 24242 20644 24298 20700
rect 24298 20644 24302 20700
rect 24238 20640 24302 20644
rect 31680 20700 31744 20704
rect 31680 20644 31684 20700
rect 31684 20644 31740 20700
rect 31740 20644 31744 20700
rect 31680 20640 31744 20644
rect 31760 20700 31824 20704
rect 31760 20644 31764 20700
rect 31764 20644 31820 20700
rect 31820 20644 31824 20700
rect 31760 20640 31824 20644
rect 31840 20700 31904 20704
rect 31840 20644 31844 20700
rect 31844 20644 31900 20700
rect 31900 20644 31904 20700
rect 31840 20640 31904 20644
rect 31920 20700 31984 20704
rect 31920 20644 31924 20700
rect 31924 20644 31980 20700
rect 31980 20644 31984 20700
rect 31920 20640 31984 20644
rect 14596 20572 14660 20636
rect 19196 20572 19260 20636
rect 26740 20572 26804 20636
rect 27292 20572 27356 20636
rect 23060 20436 23124 20500
rect 30236 20436 30300 20500
rect 27108 20300 27172 20364
rect 27292 20300 27356 20364
rect 28396 20300 28460 20364
rect 27660 20164 27724 20228
rect 30052 20164 30116 20228
rect 4793 20156 4857 20160
rect 4793 20100 4797 20156
rect 4797 20100 4853 20156
rect 4853 20100 4857 20156
rect 4793 20096 4857 20100
rect 4873 20156 4937 20160
rect 4873 20100 4877 20156
rect 4877 20100 4933 20156
rect 4933 20100 4937 20156
rect 4873 20096 4937 20100
rect 4953 20156 5017 20160
rect 4953 20100 4957 20156
rect 4957 20100 5013 20156
rect 5013 20100 5017 20156
rect 4953 20096 5017 20100
rect 5033 20156 5097 20160
rect 5033 20100 5037 20156
rect 5037 20100 5093 20156
rect 5093 20100 5097 20156
rect 5033 20096 5097 20100
rect 12475 20156 12539 20160
rect 12475 20100 12479 20156
rect 12479 20100 12535 20156
rect 12535 20100 12539 20156
rect 12475 20096 12539 20100
rect 12555 20156 12619 20160
rect 12555 20100 12559 20156
rect 12559 20100 12615 20156
rect 12615 20100 12619 20156
rect 12555 20096 12619 20100
rect 12635 20156 12699 20160
rect 12635 20100 12639 20156
rect 12639 20100 12695 20156
rect 12695 20100 12699 20156
rect 12635 20096 12699 20100
rect 12715 20156 12779 20160
rect 12715 20100 12719 20156
rect 12719 20100 12775 20156
rect 12775 20100 12779 20156
rect 12715 20096 12779 20100
rect 20157 20156 20221 20160
rect 20157 20100 20161 20156
rect 20161 20100 20217 20156
rect 20217 20100 20221 20156
rect 20157 20096 20221 20100
rect 20237 20156 20301 20160
rect 20237 20100 20241 20156
rect 20241 20100 20297 20156
rect 20297 20100 20301 20156
rect 20237 20096 20301 20100
rect 20317 20156 20381 20160
rect 20317 20100 20321 20156
rect 20321 20100 20377 20156
rect 20377 20100 20381 20156
rect 20317 20096 20381 20100
rect 20397 20156 20461 20160
rect 20397 20100 20401 20156
rect 20401 20100 20457 20156
rect 20457 20100 20461 20156
rect 20397 20096 20461 20100
rect 27839 20156 27903 20160
rect 27839 20100 27843 20156
rect 27843 20100 27899 20156
rect 27899 20100 27903 20156
rect 27839 20096 27903 20100
rect 27919 20156 27983 20160
rect 27919 20100 27923 20156
rect 27923 20100 27979 20156
rect 27979 20100 27983 20156
rect 27919 20096 27983 20100
rect 27999 20156 28063 20160
rect 27999 20100 28003 20156
rect 28003 20100 28059 20156
rect 28059 20100 28063 20156
rect 27999 20096 28063 20100
rect 28079 20156 28143 20160
rect 28079 20100 28083 20156
rect 28083 20100 28139 20156
rect 28139 20100 28143 20156
rect 28079 20096 28143 20100
rect 12940 20028 13004 20092
rect 19012 20028 19076 20092
rect 19380 20028 19444 20092
rect 17172 19892 17236 19956
rect 18460 19892 18524 19956
rect 26004 20028 26068 20092
rect 26372 20028 26436 20092
rect 28580 20028 28644 20092
rect 28948 20028 29012 20092
rect 23060 19892 23124 19956
rect 23244 19892 23308 19956
rect 24900 19756 24964 19820
rect 25636 19816 25700 19820
rect 25636 19760 25686 19816
rect 25686 19760 25700 19816
rect 25636 19756 25700 19760
rect 26924 19816 26988 19820
rect 26924 19760 26938 19816
rect 26938 19760 26988 19816
rect 26924 19756 26988 19760
rect 27108 19756 27172 19820
rect 8634 19612 8698 19616
rect 8634 19556 8638 19612
rect 8638 19556 8694 19612
rect 8694 19556 8698 19612
rect 8634 19552 8698 19556
rect 8714 19612 8778 19616
rect 8714 19556 8718 19612
rect 8718 19556 8774 19612
rect 8774 19556 8778 19612
rect 8714 19552 8778 19556
rect 8794 19612 8858 19616
rect 8794 19556 8798 19612
rect 8798 19556 8854 19612
rect 8854 19556 8858 19612
rect 8794 19552 8858 19556
rect 8874 19612 8938 19616
rect 8874 19556 8878 19612
rect 8878 19556 8934 19612
rect 8934 19556 8938 19612
rect 8874 19552 8938 19556
rect 16316 19612 16380 19616
rect 16316 19556 16320 19612
rect 16320 19556 16376 19612
rect 16376 19556 16380 19612
rect 16316 19552 16380 19556
rect 16396 19612 16460 19616
rect 16396 19556 16400 19612
rect 16400 19556 16456 19612
rect 16456 19556 16460 19612
rect 16396 19552 16460 19556
rect 16476 19612 16540 19616
rect 16476 19556 16480 19612
rect 16480 19556 16536 19612
rect 16536 19556 16540 19612
rect 16476 19552 16540 19556
rect 16556 19612 16620 19616
rect 16556 19556 16560 19612
rect 16560 19556 16616 19612
rect 16616 19556 16620 19612
rect 16556 19552 16620 19556
rect 23998 19612 24062 19616
rect 23998 19556 24002 19612
rect 24002 19556 24058 19612
rect 24058 19556 24062 19612
rect 23998 19552 24062 19556
rect 24078 19612 24142 19616
rect 24078 19556 24082 19612
rect 24082 19556 24138 19612
rect 24138 19556 24142 19612
rect 24078 19552 24142 19556
rect 24158 19612 24222 19616
rect 24158 19556 24162 19612
rect 24162 19556 24218 19612
rect 24218 19556 24222 19612
rect 24158 19552 24222 19556
rect 24238 19612 24302 19616
rect 24238 19556 24242 19612
rect 24242 19556 24298 19612
rect 24298 19556 24302 19612
rect 24238 19552 24302 19556
rect 15516 19484 15580 19548
rect 15884 19484 15948 19548
rect 18644 19484 18708 19548
rect 19380 19484 19444 19548
rect 19932 19484 19996 19548
rect 29500 19484 29564 19548
rect 30420 19620 30484 19684
rect 31680 19612 31744 19616
rect 31680 19556 31684 19612
rect 31684 19556 31740 19612
rect 31740 19556 31744 19612
rect 31680 19552 31744 19556
rect 31760 19612 31824 19616
rect 31760 19556 31764 19612
rect 31764 19556 31820 19612
rect 31820 19556 31824 19612
rect 31760 19552 31824 19556
rect 31840 19612 31904 19616
rect 31840 19556 31844 19612
rect 31844 19556 31900 19612
rect 31900 19556 31904 19612
rect 31840 19552 31904 19556
rect 31920 19612 31984 19616
rect 31920 19556 31924 19612
rect 31924 19556 31980 19612
rect 31980 19556 31984 19612
rect 31920 19552 31984 19556
rect 30788 19484 30852 19548
rect 13308 19408 13372 19412
rect 13308 19352 13322 19408
rect 13322 19352 13372 19408
rect 13308 19348 13372 19352
rect 19380 19348 19444 19412
rect 20530 19348 20594 19412
rect 28212 19348 28276 19412
rect 29316 19348 29380 19412
rect 29868 19348 29932 19412
rect 30236 19408 30300 19412
rect 30236 19352 30286 19408
rect 30286 19352 30300 19408
rect 30236 19348 30300 19352
rect 4793 19068 4857 19072
rect 4793 19012 4797 19068
rect 4797 19012 4853 19068
rect 4853 19012 4857 19068
rect 4793 19008 4857 19012
rect 4873 19068 4937 19072
rect 4873 19012 4877 19068
rect 4877 19012 4933 19068
rect 4933 19012 4937 19068
rect 4873 19008 4937 19012
rect 4953 19068 5017 19072
rect 4953 19012 4957 19068
rect 4957 19012 5013 19068
rect 5013 19012 5017 19068
rect 4953 19008 5017 19012
rect 5033 19068 5097 19072
rect 5033 19012 5037 19068
rect 5037 19012 5093 19068
rect 5093 19012 5097 19068
rect 5033 19008 5097 19012
rect 12475 19068 12539 19072
rect 12475 19012 12479 19068
rect 12479 19012 12535 19068
rect 12535 19012 12539 19068
rect 12475 19008 12539 19012
rect 12555 19068 12619 19072
rect 12555 19012 12559 19068
rect 12559 19012 12615 19068
rect 12615 19012 12619 19068
rect 12555 19008 12619 19012
rect 12635 19068 12699 19072
rect 12635 19012 12639 19068
rect 12639 19012 12695 19068
rect 12695 19012 12699 19068
rect 12635 19008 12699 19012
rect 12715 19068 12779 19072
rect 12715 19012 12719 19068
rect 12719 19012 12775 19068
rect 12775 19012 12779 19068
rect 12715 19008 12779 19012
rect 12940 18804 13004 18868
rect 18828 19076 18892 19140
rect 21588 19076 21652 19140
rect 20157 19068 20221 19072
rect 20157 19012 20161 19068
rect 20161 19012 20217 19068
rect 20217 19012 20221 19068
rect 20157 19008 20221 19012
rect 20237 19068 20301 19072
rect 20237 19012 20241 19068
rect 20241 19012 20297 19068
rect 20297 19012 20301 19068
rect 20237 19008 20301 19012
rect 20317 19068 20381 19072
rect 20317 19012 20321 19068
rect 20321 19012 20377 19068
rect 20377 19012 20381 19068
rect 20317 19008 20381 19012
rect 20397 19068 20461 19072
rect 20397 19012 20401 19068
rect 20401 19012 20457 19068
rect 20457 19012 20461 19068
rect 20397 19008 20461 19012
rect 26188 19076 26252 19140
rect 26556 19076 26620 19140
rect 15700 18864 15764 18868
rect 15700 18808 15750 18864
rect 15750 18808 15764 18864
rect 15700 18804 15764 18808
rect 16068 18804 16132 18868
rect 17356 18804 17420 18868
rect 24900 18940 24964 19004
rect 26924 19136 26988 19140
rect 26924 19080 26974 19136
rect 26974 19080 26988 19136
rect 26924 19076 26988 19080
rect 28396 19076 28460 19140
rect 29316 19076 29380 19140
rect 27839 19068 27903 19072
rect 27839 19012 27843 19068
rect 27843 19012 27899 19068
rect 27899 19012 27903 19068
rect 27839 19008 27903 19012
rect 27919 19068 27983 19072
rect 27919 19012 27923 19068
rect 27923 19012 27979 19068
rect 27979 19012 27983 19068
rect 27919 19008 27983 19012
rect 27999 19068 28063 19072
rect 27999 19012 28003 19068
rect 28003 19012 28059 19068
rect 28059 19012 28063 19068
rect 27999 19008 28063 19012
rect 28079 19068 28143 19072
rect 28079 19012 28083 19068
rect 28083 19012 28139 19068
rect 28139 19012 28143 19068
rect 28079 19008 28143 19012
rect 19748 18668 19812 18732
rect 21956 18804 22020 18868
rect 21404 18668 21468 18732
rect 31340 18668 31404 18732
rect 16068 18532 16132 18596
rect 21588 18532 21652 18596
rect 30420 18532 30484 18596
rect 8634 18524 8698 18528
rect 8634 18468 8638 18524
rect 8638 18468 8694 18524
rect 8694 18468 8698 18524
rect 8634 18464 8698 18468
rect 8714 18524 8778 18528
rect 8714 18468 8718 18524
rect 8718 18468 8774 18524
rect 8774 18468 8778 18524
rect 8714 18464 8778 18468
rect 8794 18524 8858 18528
rect 8794 18468 8798 18524
rect 8798 18468 8854 18524
rect 8854 18468 8858 18524
rect 8794 18464 8858 18468
rect 8874 18524 8938 18528
rect 8874 18468 8878 18524
rect 8878 18468 8934 18524
rect 8934 18468 8938 18524
rect 8874 18464 8938 18468
rect 16316 18524 16380 18528
rect 16316 18468 16320 18524
rect 16320 18468 16376 18524
rect 16376 18468 16380 18524
rect 16316 18464 16380 18468
rect 16396 18524 16460 18528
rect 16396 18468 16400 18524
rect 16400 18468 16456 18524
rect 16456 18468 16460 18524
rect 16396 18464 16460 18468
rect 16476 18524 16540 18528
rect 16476 18468 16480 18524
rect 16480 18468 16536 18524
rect 16536 18468 16540 18524
rect 16476 18464 16540 18468
rect 16556 18524 16620 18528
rect 16556 18468 16560 18524
rect 16560 18468 16616 18524
rect 16616 18468 16620 18524
rect 16556 18464 16620 18468
rect 23998 18524 24062 18528
rect 23998 18468 24002 18524
rect 24002 18468 24058 18524
rect 24058 18468 24062 18524
rect 23998 18464 24062 18468
rect 24078 18524 24142 18528
rect 24078 18468 24082 18524
rect 24082 18468 24138 18524
rect 24138 18468 24142 18524
rect 24078 18464 24142 18468
rect 24158 18524 24222 18528
rect 24158 18468 24162 18524
rect 24162 18468 24218 18524
rect 24218 18468 24222 18524
rect 24158 18464 24222 18468
rect 24238 18524 24302 18528
rect 24238 18468 24242 18524
rect 24242 18468 24298 18524
rect 24298 18468 24302 18524
rect 24238 18464 24302 18468
rect 16804 18456 16868 18460
rect 16804 18400 16818 18456
rect 16818 18400 16868 18456
rect 16804 18396 16868 18400
rect 26004 18396 26068 18460
rect 29132 18260 29196 18324
rect 31680 18524 31744 18528
rect 31680 18468 31684 18524
rect 31684 18468 31740 18524
rect 31740 18468 31744 18524
rect 31680 18464 31744 18468
rect 31760 18524 31824 18528
rect 31760 18468 31764 18524
rect 31764 18468 31820 18524
rect 31820 18468 31824 18524
rect 31760 18464 31824 18468
rect 31840 18524 31904 18528
rect 31840 18468 31844 18524
rect 31844 18468 31900 18524
rect 31900 18468 31904 18524
rect 31840 18464 31904 18468
rect 31920 18524 31984 18528
rect 31920 18468 31924 18524
rect 31924 18468 31980 18524
rect 31980 18468 31984 18524
rect 31920 18464 31984 18468
rect 25452 18124 25516 18188
rect 26372 18184 26436 18188
rect 26372 18128 26386 18184
rect 26386 18128 26436 18184
rect 26372 18124 26436 18128
rect 24716 18048 24780 18052
rect 24716 17992 24766 18048
rect 24766 17992 24780 18048
rect 24716 17988 24780 17992
rect 27292 17988 27356 18052
rect 28396 18124 28460 18188
rect 29132 18124 29196 18188
rect 4793 17980 4857 17984
rect 4793 17924 4797 17980
rect 4797 17924 4853 17980
rect 4853 17924 4857 17980
rect 4793 17920 4857 17924
rect 4873 17980 4937 17984
rect 4873 17924 4877 17980
rect 4877 17924 4933 17980
rect 4933 17924 4937 17980
rect 4873 17920 4937 17924
rect 4953 17980 5017 17984
rect 4953 17924 4957 17980
rect 4957 17924 5013 17980
rect 5013 17924 5017 17980
rect 4953 17920 5017 17924
rect 5033 17980 5097 17984
rect 5033 17924 5037 17980
rect 5037 17924 5093 17980
rect 5093 17924 5097 17980
rect 5033 17920 5097 17924
rect 12475 17980 12539 17984
rect 12475 17924 12479 17980
rect 12479 17924 12535 17980
rect 12535 17924 12539 17980
rect 12475 17920 12539 17924
rect 12555 17980 12619 17984
rect 12555 17924 12559 17980
rect 12559 17924 12615 17980
rect 12615 17924 12619 17980
rect 12555 17920 12619 17924
rect 12635 17980 12699 17984
rect 12635 17924 12639 17980
rect 12639 17924 12695 17980
rect 12695 17924 12699 17980
rect 12635 17920 12699 17924
rect 12715 17980 12779 17984
rect 12715 17924 12719 17980
rect 12719 17924 12775 17980
rect 12775 17924 12779 17980
rect 12715 17920 12779 17924
rect 20157 17980 20221 17984
rect 20157 17924 20161 17980
rect 20161 17924 20217 17980
rect 20217 17924 20221 17980
rect 20157 17920 20221 17924
rect 20237 17980 20301 17984
rect 20237 17924 20241 17980
rect 20241 17924 20297 17980
rect 20297 17924 20301 17980
rect 20237 17920 20301 17924
rect 20317 17980 20381 17984
rect 20317 17924 20321 17980
rect 20321 17924 20377 17980
rect 20377 17924 20381 17980
rect 20317 17920 20381 17924
rect 20397 17980 20461 17984
rect 20397 17924 20401 17980
rect 20401 17924 20457 17980
rect 20457 17924 20461 17980
rect 20397 17920 20461 17924
rect 27839 17980 27903 17984
rect 27839 17924 27843 17980
rect 27843 17924 27899 17980
rect 27899 17924 27903 17980
rect 27839 17920 27903 17924
rect 27919 17980 27983 17984
rect 27919 17924 27923 17980
rect 27923 17924 27979 17980
rect 27979 17924 27983 17980
rect 27919 17920 27983 17924
rect 27999 17980 28063 17984
rect 27999 17924 28003 17980
rect 28003 17924 28059 17980
rect 28059 17924 28063 17980
rect 27999 17920 28063 17924
rect 28079 17980 28143 17984
rect 28079 17924 28083 17980
rect 28083 17924 28139 17980
rect 28139 17924 28143 17980
rect 28079 17920 28143 17924
rect 14044 17716 14108 17780
rect 16804 17852 16868 17916
rect 16988 17852 17052 17916
rect 21220 17852 21284 17916
rect 30236 17912 30300 17916
rect 30236 17856 30286 17912
rect 30286 17856 30300 17912
rect 30236 17852 30300 17856
rect 17172 17716 17236 17780
rect 24900 17716 24964 17780
rect 26188 17776 26252 17780
rect 26188 17720 26238 17776
rect 26238 17720 26252 17776
rect 26188 17716 26252 17720
rect 27476 17716 27540 17780
rect 28764 17716 28828 17780
rect 29684 17580 29748 17644
rect 8634 17436 8698 17440
rect 8634 17380 8638 17436
rect 8638 17380 8694 17436
rect 8694 17380 8698 17436
rect 8634 17376 8698 17380
rect 8714 17436 8778 17440
rect 8714 17380 8718 17436
rect 8718 17380 8774 17436
rect 8774 17380 8778 17436
rect 8714 17376 8778 17380
rect 8794 17436 8858 17440
rect 8794 17380 8798 17436
rect 8798 17380 8854 17436
rect 8854 17380 8858 17436
rect 8794 17376 8858 17380
rect 8874 17436 8938 17440
rect 8874 17380 8878 17436
rect 8878 17380 8934 17436
rect 8934 17380 8938 17436
rect 8874 17376 8938 17380
rect 16316 17436 16380 17440
rect 16316 17380 16320 17436
rect 16320 17380 16376 17436
rect 16376 17380 16380 17436
rect 16316 17376 16380 17380
rect 16396 17436 16460 17440
rect 16396 17380 16400 17436
rect 16400 17380 16456 17436
rect 16456 17380 16460 17436
rect 16396 17376 16460 17380
rect 16476 17436 16540 17440
rect 16476 17380 16480 17436
rect 16480 17380 16536 17436
rect 16536 17380 16540 17436
rect 16476 17376 16540 17380
rect 16556 17436 16620 17440
rect 16556 17380 16560 17436
rect 16560 17380 16616 17436
rect 16616 17380 16620 17436
rect 16556 17376 16620 17380
rect 17172 17308 17236 17372
rect 10916 17172 10980 17236
rect 10548 16960 10612 16964
rect 10548 16904 10562 16960
rect 10562 16904 10612 16960
rect 10548 16900 10612 16904
rect 27108 17444 27172 17508
rect 27660 17444 27724 17508
rect 28580 17444 28644 17508
rect 23998 17436 24062 17440
rect 23998 17380 24002 17436
rect 24002 17380 24058 17436
rect 24058 17380 24062 17436
rect 23998 17376 24062 17380
rect 24078 17436 24142 17440
rect 24078 17380 24082 17436
rect 24082 17380 24138 17436
rect 24138 17380 24142 17436
rect 24078 17376 24142 17380
rect 24158 17436 24222 17440
rect 24158 17380 24162 17436
rect 24162 17380 24218 17436
rect 24218 17380 24222 17436
rect 24158 17376 24222 17380
rect 24238 17436 24302 17440
rect 24238 17380 24242 17436
rect 24242 17380 24298 17436
rect 24298 17380 24302 17436
rect 24238 17376 24302 17380
rect 31680 17436 31744 17440
rect 31680 17380 31684 17436
rect 31684 17380 31740 17436
rect 31740 17380 31744 17436
rect 31680 17376 31744 17380
rect 31760 17436 31824 17440
rect 31760 17380 31764 17436
rect 31764 17380 31820 17436
rect 31820 17380 31824 17436
rect 31760 17376 31824 17380
rect 31840 17436 31904 17440
rect 31840 17380 31844 17436
rect 31844 17380 31900 17436
rect 31900 17380 31904 17436
rect 31840 17376 31904 17380
rect 31920 17436 31984 17440
rect 31920 17380 31924 17436
rect 31924 17380 31980 17436
rect 31980 17380 31984 17436
rect 31920 17376 31984 17380
rect 30236 17308 30300 17372
rect 26372 17172 26436 17236
rect 16068 16900 16132 16964
rect 31524 17036 31588 17100
rect 17356 16900 17420 16964
rect 26004 16900 26068 16964
rect 26924 16900 26988 16964
rect 4793 16892 4857 16896
rect 4793 16836 4797 16892
rect 4797 16836 4853 16892
rect 4853 16836 4857 16892
rect 4793 16832 4857 16836
rect 4873 16892 4937 16896
rect 4873 16836 4877 16892
rect 4877 16836 4933 16892
rect 4933 16836 4937 16892
rect 4873 16832 4937 16836
rect 4953 16892 5017 16896
rect 4953 16836 4957 16892
rect 4957 16836 5013 16892
rect 5013 16836 5017 16892
rect 4953 16832 5017 16836
rect 5033 16892 5097 16896
rect 5033 16836 5037 16892
rect 5037 16836 5093 16892
rect 5093 16836 5097 16892
rect 5033 16832 5097 16836
rect 12475 16892 12539 16896
rect 12475 16836 12479 16892
rect 12479 16836 12535 16892
rect 12535 16836 12539 16892
rect 12475 16832 12539 16836
rect 12555 16892 12619 16896
rect 12555 16836 12559 16892
rect 12559 16836 12615 16892
rect 12615 16836 12619 16892
rect 12555 16832 12619 16836
rect 12635 16892 12699 16896
rect 12635 16836 12639 16892
rect 12639 16836 12695 16892
rect 12695 16836 12699 16892
rect 12635 16832 12699 16836
rect 12715 16892 12779 16896
rect 12715 16836 12719 16892
rect 12719 16836 12775 16892
rect 12775 16836 12779 16892
rect 12715 16832 12779 16836
rect 20157 16892 20221 16896
rect 20157 16836 20161 16892
rect 20161 16836 20217 16892
rect 20217 16836 20221 16892
rect 20157 16832 20221 16836
rect 20237 16892 20301 16896
rect 20237 16836 20241 16892
rect 20241 16836 20297 16892
rect 20297 16836 20301 16892
rect 20237 16832 20301 16836
rect 20317 16892 20381 16896
rect 20317 16836 20321 16892
rect 20321 16836 20377 16892
rect 20377 16836 20381 16892
rect 20317 16832 20381 16836
rect 20397 16892 20461 16896
rect 20397 16836 20401 16892
rect 20401 16836 20457 16892
rect 20457 16836 20461 16892
rect 20397 16832 20461 16836
rect 27839 16892 27903 16896
rect 27839 16836 27843 16892
rect 27843 16836 27899 16892
rect 27899 16836 27903 16892
rect 27839 16832 27903 16836
rect 27919 16892 27983 16896
rect 27919 16836 27923 16892
rect 27923 16836 27979 16892
rect 27979 16836 27983 16892
rect 27919 16832 27983 16836
rect 27999 16892 28063 16896
rect 27999 16836 28003 16892
rect 28003 16836 28059 16892
rect 28059 16836 28063 16892
rect 27999 16832 28063 16836
rect 28079 16892 28143 16896
rect 28079 16836 28083 16892
rect 28083 16836 28139 16892
rect 28139 16836 28143 16892
rect 28079 16832 28143 16836
rect 23796 16824 23860 16828
rect 23796 16768 23810 16824
rect 23810 16768 23860 16824
rect 23796 16764 23860 16768
rect 26924 16824 26988 16828
rect 26924 16768 26974 16824
rect 26974 16768 26988 16824
rect 26924 16764 26988 16768
rect 23612 16628 23676 16692
rect 10732 16492 10796 16556
rect 12204 16552 12268 16556
rect 12204 16496 12218 16552
rect 12218 16496 12268 16552
rect 12204 16492 12268 16496
rect 25820 16492 25884 16556
rect 28396 16764 28460 16828
rect 29132 16900 29196 16964
rect 30604 16900 30668 16964
rect 28396 16628 28460 16692
rect 29132 16764 29196 16828
rect 29500 16628 29564 16692
rect 28948 16492 29012 16556
rect 29500 16492 29564 16556
rect 30052 16628 30116 16692
rect 30972 16628 31036 16692
rect 30052 16492 30116 16556
rect 8634 16348 8698 16352
rect 8634 16292 8638 16348
rect 8638 16292 8694 16348
rect 8694 16292 8698 16348
rect 8634 16288 8698 16292
rect 8714 16348 8778 16352
rect 8714 16292 8718 16348
rect 8718 16292 8774 16348
rect 8774 16292 8778 16348
rect 8714 16288 8778 16292
rect 8794 16348 8858 16352
rect 8794 16292 8798 16348
rect 8798 16292 8854 16348
rect 8854 16292 8858 16348
rect 8794 16288 8858 16292
rect 8874 16348 8938 16352
rect 8874 16292 8878 16348
rect 8878 16292 8934 16348
rect 8934 16292 8938 16348
rect 8874 16288 8938 16292
rect 15148 16280 15212 16284
rect 16316 16348 16380 16352
rect 16316 16292 16320 16348
rect 16320 16292 16376 16348
rect 16376 16292 16380 16348
rect 16316 16288 16380 16292
rect 16396 16348 16460 16352
rect 16396 16292 16400 16348
rect 16400 16292 16456 16348
rect 16456 16292 16460 16348
rect 16396 16288 16460 16292
rect 16476 16348 16540 16352
rect 16476 16292 16480 16348
rect 16480 16292 16536 16348
rect 16536 16292 16540 16348
rect 16476 16288 16540 16292
rect 16556 16348 16620 16352
rect 16556 16292 16560 16348
rect 16560 16292 16616 16348
rect 16616 16292 16620 16348
rect 16556 16288 16620 16292
rect 15148 16224 15198 16280
rect 15198 16224 15212 16280
rect 15148 16220 15212 16224
rect 19012 16280 19076 16284
rect 19012 16224 19062 16280
rect 19062 16224 19076 16280
rect 19012 16220 19076 16224
rect 23998 16348 24062 16352
rect 23998 16292 24002 16348
rect 24002 16292 24058 16348
rect 24058 16292 24062 16348
rect 23998 16288 24062 16292
rect 24078 16348 24142 16352
rect 24078 16292 24082 16348
rect 24082 16292 24138 16348
rect 24138 16292 24142 16348
rect 24078 16288 24142 16292
rect 24158 16348 24222 16352
rect 24158 16292 24162 16348
rect 24162 16292 24218 16348
rect 24218 16292 24222 16348
rect 24158 16288 24222 16292
rect 24238 16348 24302 16352
rect 24238 16292 24242 16348
rect 24242 16292 24298 16348
rect 24298 16292 24302 16348
rect 24238 16288 24302 16292
rect 31680 16348 31744 16352
rect 31680 16292 31684 16348
rect 31684 16292 31740 16348
rect 31740 16292 31744 16348
rect 31680 16288 31744 16292
rect 31760 16348 31824 16352
rect 31760 16292 31764 16348
rect 31764 16292 31820 16348
rect 31820 16292 31824 16348
rect 31760 16288 31824 16292
rect 31840 16348 31904 16352
rect 31840 16292 31844 16348
rect 31844 16292 31900 16348
rect 31900 16292 31904 16348
rect 31840 16288 31904 16292
rect 31920 16348 31984 16352
rect 31920 16292 31924 16348
rect 31924 16292 31980 16348
rect 31980 16292 31984 16348
rect 31920 16288 31984 16292
rect 30420 15948 30484 16012
rect 30788 16008 30852 16012
rect 30788 15952 30802 16008
rect 30802 15952 30852 16008
rect 30788 15948 30852 15952
rect 4793 15804 4857 15808
rect 4793 15748 4797 15804
rect 4797 15748 4853 15804
rect 4853 15748 4857 15804
rect 4793 15744 4857 15748
rect 4873 15804 4937 15808
rect 4873 15748 4877 15804
rect 4877 15748 4933 15804
rect 4933 15748 4937 15804
rect 4873 15744 4937 15748
rect 4953 15804 5017 15808
rect 4953 15748 4957 15804
rect 4957 15748 5013 15804
rect 5013 15748 5017 15804
rect 4953 15744 5017 15748
rect 5033 15804 5097 15808
rect 5033 15748 5037 15804
rect 5037 15748 5093 15804
rect 5093 15748 5097 15804
rect 5033 15744 5097 15748
rect 12475 15804 12539 15808
rect 12475 15748 12479 15804
rect 12479 15748 12535 15804
rect 12535 15748 12539 15804
rect 12475 15744 12539 15748
rect 12555 15804 12619 15808
rect 12555 15748 12559 15804
rect 12559 15748 12615 15804
rect 12615 15748 12619 15804
rect 12555 15744 12619 15748
rect 12635 15804 12699 15808
rect 12635 15748 12639 15804
rect 12639 15748 12695 15804
rect 12695 15748 12699 15804
rect 12635 15744 12699 15748
rect 12715 15804 12779 15808
rect 12715 15748 12719 15804
rect 12719 15748 12775 15804
rect 12775 15748 12779 15804
rect 12715 15744 12779 15748
rect 20157 15804 20221 15808
rect 20157 15748 20161 15804
rect 20161 15748 20217 15804
rect 20217 15748 20221 15804
rect 20157 15744 20221 15748
rect 20237 15804 20301 15808
rect 20237 15748 20241 15804
rect 20241 15748 20297 15804
rect 20297 15748 20301 15804
rect 20237 15744 20301 15748
rect 20317 15804 20381 15808
rect 20317 15748 20321 15804
rect 20321 15748 20377 15804
rect 20377 15748 20381 15804
rect 20317 15744 20381 15748
rect 20397 15804 20461 15808
rect 20397 15748 20401 15804
rect 20401 15748 20457 15804
rect 20457 15748 20461 15804
rect 20397 15744 20461 15748
rect 27839 15804 27903 15808
rect 27839 15748 27843 15804
rect 27843 15748 27899 15804
rect 27899 15748 27903 15804
rect 27839 15744 27903 15748
rect 27919 15804 27983 15808
rect 27919 15748 27923 15804
rect 27923 15748 27979 15804
rect 27979 15748 27983 15804
rect 27919 15744 27983 15748
rect 27999 15804 28063 15808
rect 27999 15748 28003 15804
rect 28003 15748 28059 15804
rect 28059 15748 28063 15804
rect 27999 15744 28063 15748
rect 28079 15804 28143 15808
rect 28079 15748 28083 15804
rect 28083 15748 28139 15804
rect 28139 15748 28143 15804
rect 28079 15744 28143 15748
rect 16804 15540 16868 15604
rect 29132 15540 29196 15604
rect 24532 15404 24596 15468
rect 26740 15404 26804 15468
rect 11652 15268 11716 15332
rect 16068 15268 16132 15332
rect 17908 15268 17972 15332
rect 21404 15268 21468 15332
rect 24900 15268 24964 15332
rect 25820 15268 25884 15332
rect 30236 15268 30300 15332
rect 8634 15260 8698 15264
rect 8634 15204 8638 15260
rect 8638 15204 8694 15260
rect 8694 15204 8698 15260
rect 8634 15200 8698 15204
rect 8714 15260 8778 15264
rect 8714 15204 8718 15260
rect 8718 15204 8774 15260
rect 8774 15204 8778 15260
rect 8714 15200 8778 15204
rect 8794 15260 8858 15264
rect 8794 15204 8798 15260
rect 8798 15204 8854 15260
rect 8854 15204 8858 15260
rect 8794 15200 8858 15204
rect 8874 15260 8938 15264
rect 8874 15204 8878 15260
rect 8878 15204 8934 15260
rect 8934 15204 8938 15260
rect 8874 15200 8938 15204
rect 16316 15260 16380 15264
rect 16316 15204 16320 15260
rect 16320 15204 16376 15260
rect 16376 15204 16380 15260
rect 16316 15200 16380 15204
rect 16396 15260 16460 15264
rect 16396 15204 16400 15260
rect 16400 15204 16456 15260
rect 16456 15204 16460 15260
rect 16396 15200 16460 15204
rect 16476 15260 16540 15264
rect 16476 15204 16480 15260
rect 16480 15204 16536 15260
rect 16536 15204 16540 15260
rect 16476 15200 16540 15204
rect 16556 15260 16620 15264
rect 16556 15204 16560 15260
rect 16560 15204 16616 15260
rect 16616 15204 16620 15260
rect 16556 15200 16620 15204
rect 23998 15260 24062 15264
rect 23998 15204 24002 15260
rect 24002 15204 24058 15260
rect 24058 15204 24062 15260
rect 23998 15200 24062 15204
rect 24078 15260 24142 15264
rect 24078 15204 24082 15260
rect 24082 15204 24138 15260
rect 24138 15204 24142 15260
rect 24078 15200 24142 15204
rect 24158 15260 24222 15264
rect 24158 15204 24162 15260
rect 24162 15204 24218 15260
rect 24218 15204 24222 15260
rect 24158 15200 24222 15204
rect 24238 15260 24302 15264
rect 24238 15204 24242 15260
rect 24242 15204 24298 15260
rect 24298 15204 24302 15260
rect 24238 15200 24302 15204
rect 31680 15260 31744 15264
rect 31680 15204 31684 15260
rect 31684 15204 31740 15260
rect 31740 15204 31744 15260
rect 31680 15200 31744 15204
rect 31760 15260 31824 15264
rect 31760 15204 31764 15260
rect 31764 15204 31820 15260
rect 31820 15204 31824 15260
rect 31760 15200 31824 15204
rect 31840 15260 31904 15264
rect 31840 15204 31844 15260
rect 31844 15204 31900 15260
rect 31900 15204 31904 15260
rect 31840 15200 31904 15204
rect 31920 15260 31984 15264
rect 31920 15204 31924 15260
rect 31924 15204 31980 15260
rect 31980 15204 31984 15260
rect 31920 15200 31984 15204
rect 21404 15132 21468 15196
rect 25636 15132 25700 15196
rect 31524 15132 31588 15196
rect 4793 14716 4857 14720
rect 4793 14660 4797 14716
rect 4797 14660 4853 14716
rect 4853 14660 4857 14716
rect 4793 14656 4857 14660
rect 4873 14716 4937 14720
rect 4873 14660 4877 14716
rect 4877 14660 4933 14716
rect 4933 14660 4937 14716
rect 4873 14656 4937 14660
rect 4953 14716 5017 14720
rect 4953 14660 4957 14716
rect 4957 14660 5013 14716
rect 5013 14660 5017 14716
rect 4953 14656 5017 14660
rect 5033 14716 5097 14720
rect 5033 14660 5037 14716
rect 5037 14660 5093 14716
rect 5093 14660 5097 14716
rect 5033 14656 5097 14660
rect 12475 14716 12539 14720
rect 12475 14660 12479 14716
rect 12479 14660 12535 14716
rect 12535 14660 12539 14716
rect 12475 14656 12539 14660
rect 12555 14716 12619 14720
rect 12555 14660 12559 14716
rect 12559 14660 12615 14716
rect 12615 14660 12619 14716
rect 12555 14656 12619 14660
rect 12635 14716 12699 14720
rect 12635 14660 12639 14716
rect 12639 14660 12695 14716
rect 12695 14660 12699 14716
rect 12635 14656 12699 14660
rect 12715 14716 12779 14720
rect 12715 14660 12719 14716
rect 12719 14660 12775 14716
rect 12775 14660 12779 14716
rect 12715 14656 12779 14660
rect 20852 14724 20916 14788
rect 29316 14724 29380 14788
rect 20157 14716 20221 14720
rect 20157 14660 20161 14716
rect 20161 14660 20217 14716
rect 20217 14660 20221 14716
rect 20157 14656 20221 14660
rect 20237 14716 20301 14720
rect 20237 14660 20241 14716
rect 20241 14660 20297 14716
rect 20297 14660 20301 14716
rect 20237 14656 20301 14660
rect 20317 14716 20381 14720
rect 20317 14660 20321 14716
rect 20321 14660 20377 14716
rect 20377 14660 20381 14716
rect 20317 14656 20381 14660
rect 20397 14716 20461 14720
rect 20397 14660 20401 14716
rect 20401 14660 20457 14716
rect 20457 14660 20461 14716
rect 20397 14656 20461 14660
rect 27839 14716 27903 14720
rect 27839 14660 27843 14716
rect 27843 14660 27899 14716
rect 27899 14660 27903 14716
rect 27839 14656 27903 14660
rect 27919 14716 27983 14720
rect 27919 14660 27923 14716
rect 27923 14660 27979 14716
rect 27979 14660 27983 14716
rect 27919 14656 27983 14660
rect 27999 14716 28063 14720
rect 27999 14660 28003 14716
rect 28003 14660 28059 14716
rect 28059 14660 28063 14716
rect 27999 14656 28063 14660
rect 28079 14716 28143 14720
rect 28079 14660 28083 14716
rect 28083 14660 28139 14716
rect 28139 14660 28143 14716
rect 28079 14656 28143 14660
rect 19564 14588 19628 14652
rect 29684 14588 29748 14652
rect 8634 14172 8698 14176
rect 8634 14116 8638 14172
rect 8638 14116 8694 14172
rect 8694 14116 8698 14172
rect 8634 14112 8698 14116
rect 8714 14172 8778 14176
rect 8714 14116 8718 14172
rect 8718 14116 8774 14172
rect 8774 14116 8778 14172
rect 8714 14112 8778 14116
rect 8794 14172 8858 14176
rect 8794 14116 8798 14172
rect 8798 14116 8854 14172
rect 8854 14116 8858 14172
rect 8794 14112 8858 14116
rect 8874 14172 8938 14176
rect 8874 14116 8878 14172
rect 8878 14116 8934 14172
rect 8934 14116 8938 14172
rect 8874 14112 8938 14116
rect 12020 14044 12084 14108
rect 25268 14452 25332 14516
rect 23060 14316 23124 14380
rect 15148 14180 15212 14244
rect 21588 14180 21652 14244
rect 16316 14172 16380 14176
rect 16316 14116 16320 14172
rect 16320 14116 16376 14172
rect 16376 14116 16380 14172
rect 16316 14112 16380 14116
rect 16396 14172 16460 14176
rect 16396 14116 16400 14172
rect 16400 14116 16456 14172
rect 16456 14116 16460 14172
rect 16396 14112 16460 14116
rect 16476 14172 16540 14176
rect 16476 14116 16480 14172
rect 16480 14116 16536 14172
rect 16536 14116 16540 14172
rect 16476 14112 16540 14116
rect 16556 14172 16620 14176
rect 16556 14116 16560 14172
rect 16560 14116 16616 14172
rect 16616 14116 16620 14172
rect 16556 14112 16620 14116
rect 23998 14172 24062 14176
rect 23998 14116 24002 14172
rect 24002 14116 24058 14172
rect 24058 14116 24062 14172
rect 23998 14112 24062 14116
rect 24078 14172 24142 14176
rect 24078 14116 24082 14172
rect 24082 14116 24138 14172
rect 24138 14116 24142 14172
rect 24078 14112 24142 14116
rect 24158 14172 24222 14176
rect 24158 14116 24162 14172
rect 24162 14116 24218 14172
rect 24218 14116 24222 14172
rect 24158 14112 24222 14116
rect 24238 14172 24302 14176
rect 24238 14116 24242 14172
rect 24242 14116 24298 14172
rect 24298 14116 24302 14172
rect 24238 14112 24302 14116
rect 15516 14044 15580 14108
rect 19012 13908 19076 13972
rect 31680 14172 31744 14176
rect 31680 14116 31684 14172
rect 31684 14116 31740 14172
rect 31740 14116 31744 14172
rect 31680 14112 31744 14116
rect 31760 14172 31824 14176
rect 31760 14116 31764 14172
rect 31764 14116 31820 14172
rect 31820 14116 31824 14172
rect 31760 14112 31824 14116
rect 31840 14172 31904 14176
rect 31840 14116 31844 14172
rect 31844 14116 31900 14172
rect 31900 14116 31904 14172
rect 31840 14112 31904 14116
rect 31920 14172 31984 14176
rect 31920 14116 31924 14172
rect 31924 14116 31980 14172
rect 31980 14116 31984 14172
rect 31920 14112 31984 14116
rect 26004 13908 26068 13972
rect 20852 13772 20916 13836
rect 25268 13772 25332 13836
rect 25820 13772 25884 13836
rect 26556 13772 26620 13836
rect 28212 13832 28276 13836
rect 28212 13776 28226 13832
rect 28226 13776 28276 13832
rect 28212 13772 28276 13776
rect 29868 13772 29932 13836
rect 4793 13628 4857 13632
rect 4793 13572 4797 13628
rect 4797 13572 4853 13628
rect 4853 13572 4857 13628
rect 4793 13568 4857 13572
rect 4873 13628 4937 13632
rect 4873 13572 4877 13628
rect 4877 13572 4933 13628
rect 4933 13572 4937 13628
rect 4873 13568 4937 13572
rect 4953 13628 5017 13632
rect 4953 13572 4957 13628
rect 4957 13572 5013 13628
rect 5013 13572 5017 13628
rect 4953 13568 5017 13572
rect 5033 13628 5097 13632
rect 5033 13572 5037 13628
rect 5037 13572 5093 13628
rect 5093 13572 5097 13628
rect 5033 13568 5097 13572
rect 12475 13628 12539 13632
rect 12475 13572 12479 13628
rect 12479 13572 12535 13628
rect 12535 13572 12539 13628
rect 12475 13568 12539 13572
rect 12555 13628 12619 13632
rect 12555 13572 12559 13628
rect 12559 13572 12615 13628
rect 12615 13572 12619 13628
rect 12555 13568 12619 13572
rect 12635 13628 12699 13632
rect 12635 13572 12639 13628
rect 12639 13572 12695 13628
rect 12695 13572 12699 13628
rect 12635 13568 12699 13572
rect 12715 13628 12779 13632
rect 12715 13572 12719 13628
rect 12719 13572 12775 13628
rect 12775 13572 12779 13628
rect 12715 13568 12779 13572
rect 20157 13628 20221 13632
rect 20157 13572 20161 13628
rect 20161 13572 20217 13628
rect 20217 13572 20221 13628
rect 20157 13568 20221 13572
rect 20237 13628 20301 13632
rect 20237 13572 20241 13628
rect 20241 13572 20297 13628
rect 20297 13572 20301 13628
rect 20237 13568 20301 13572
rect 20317 13628 20381 13632
rect 20317 13572 20321 13628
rect 20321 13572 20377 13628
rect 20377 13572 20381 13628
rect 20317 13568 20381 13572
rect 20397 13628 20461 13632
rect 20397 13572 20401 13628
rect 20401 13572 20457 13628
rect 20457 13572 20461 13628
rect 20397 13568 20461 13572
rect 27839 13628 27903 13632
rect 27839 13572 27843 13628
rect 27843 13572 27899 13628
rect 27899 13572 27903 13628
rect 27839 13568 27903 13572
rect 27919 13628 27983 13632
rect 27919 13572 27923 13628
rect 27923 13572 27979 13628
rect 27979 13572 27983 13628
rect 27919 13568 27983 13572
rect 27999 13628 28063 13632
rect 27999 13572 28003 13628
rect 28003 13572 28059 13628
rect 28059 13572 28063 13628
rect 27999 13568 28063 13572
rect 28079 13628 28143 13632
rect 28079 13572 28083 13628
rect 28083 13572 28139 13628
rect 28139 13572 28143 13628
rect 28079 13568 28143 13572
rect 6868 13364 6932 13428
rect 21036 13500 21100 13564
rect 31156 13560 31220 13564
rect 31156 13504 31170 13560
rect 31170 13504 31220 13560
rect 31156 13500 31220 13504
rect 21956 13092 22020 13156
rect 25452 13152 25516 13156
rect 25452 13096 25502 13152
rect 25502 13096 25516 13152
rect 25452 13092 25516 13096
rect 27660 13092 27724 13156
rect 8634 13084 8698 13088
rect 8634 13028 8638 13084
rect 8638 13028 8694 13084
rect 8694 13028 8698 13084
rect 8634 13024 8698 13028
rect 8714 13084 8778 13088
rect 8714 13028 8718 13084
rect 8718 13028 8774 13084
rect 8774 13028 8778 13084
rect 8714 13024 8778 13028
rect 8794 13084 8858 13088
rect 8794 13028 8798 13084
rect 8798 13028 8854 13084
rect 8854 13028 8858 13084
rect 8794 13024 8858 13028
rect 8874 13084 8938 13088
rect 8874 13028 8878 13084
rect 8878 13028 8934 13084
rect 8934 13028 8938 13084
rect 8874 13024 8938 13028
rect 16316 13084 16380 13088
rect 16316 13028 16320 13084
rect 16320 13028 16376 13084
rect 16376 13028 16380 13084
rect 16316 13024 16380 13028
rect 16396 13084 16460 13088
rect 16396 13028 16400 13084
rect 16400 13028 16456 13084
rect 16456 13028 16460 13084
rect 16396 13024 16460 13028
rect 16476 13084 16540 13088
rect 16476 13028 16480 13084
rect 16480 13028 16536 13084
rect 16536 13028 16540 13084
rect 16476 13024 16540 13028
rect 16556 13084 16620 13088
rect 16556 13028 16560 13084
rect 16560 13028 16616 13084
rect 16616 13028 16620 13084
rect 16556 13024 16620 13028
rect 23998 13084 24062 13088
rect 23998 13028 24002 13084
rect 24002 13028 24058 13084
rect 24058 13028 24062 13084
rect 23998 13024 24062 13028
rect 24078 13084 24142 13088
rect 24078 13028 24082 13084
rect 24082 13028 24138 13084
rect 24138 13028 24142 13084
rect 24078 13024 24142 13028
rect 24158 13084 24222 13088
rect 24158 13028 24162 13084
rect 24162 13028 24218 13084
rect 24218 13028 24222 13084
rect 24158 13024 24222 13028
rect 24238 13084 24302 13088
rect 24238 13028 24242 13084
rect 24242 13028 24298 13084
rect 24298 13028 24302 13084
rect 24238 13024 24302 13028
rect 31680 13084 31744 13088
rect 31680 13028 31684 13084
rect 31684 13028 31740 13084
rect 31740 13028 31744 13084
rect 31680 13024 31744 13028
rect 31760 13084 31824 13088
rect 31760 13028 31764 13084
rect 31764 13028 31820 13084
rect 31820 13028 31824 13084
rect 31760 13024 31824 13028
rect 31840 13084 31904 13088
rect 31840 13028 31844 13084
rect 31844 13028 31900 13084
rect 31900 13028 31904 13084
rect 31840 13024 31904 13028
rect 31920 13084 31984 13088
rect 31920 13028 31924 13084
rect 31924 13028 31980 13084
rect 31980 13028 31984 13084
rect 31920 13024 31984 13028
rect 26372 12956 26436 13020
rect 29500 12956 29564 13020
rect 23796 12820 23860 12884
rect 27292 12820 27356 12884
rect 28396 12820 28460 12884
rect 21404 12548 21468 12612
rect 28948 12684 29012 12748
rect 4793 12540 4857 12544
rect 4793 12484 4797 12540
rect 4797 12484 4853 12540
rect 4853 12484 4857 12540
rect 4793 12480 4857 12484
rect 4873 12540 4937 12544
rect 4873 12484 4877 12540
rect 4877 12484 4933 12540
rect 4933 12484 4937 12540
rect 4873 12480 4937 12484
rect 4953 12540 5017 12544
rect 4953 12484 4957 12540
rect 4957 12484 5013 12540
rect 5013 12484 5017 12540
rect 4953 12480 5017 12484
rect 5033 12540 5097 12544
rect 5033 12484 5037 12540
rect 5037 12484 5093 12540
rect 5093 12484 5097 12540
rect 5033 12480 5097 12484
rect 12475 12540 12539 12544
rect 12475 12484 12479 12540
rect 12479 12484 12535 12540
rect 12535 12484 12539 12540
rect 12475 12480 12539 12484
rect 12555 12540 12619 12544
rect 12555 12484 12559 12540
rect 12559 12484 12615 12540
rect 12615 12484 12619 12540
rect 12555 12480 12619 12484
rect 12635 12540 12699 12544
rect 12635 12484 12639 12540
rect 12639 12484 12695 12540
rect 12695 12484 12699 12540
rect 12635 12480 12699 12484
rect 12715 12540 12779 12544
rect 12715 12484 12719 12540
rect 12719 12484 12775 12540
rect 12775 12484 12779 12540
rect 12715 12480 12779 12484
rect 20157 12540 20221 12544
rect 20157 12484 20161 12540
rect 20161 12484 20217 12540
rect 20217 12484 20221 12540
rect 20157 12480 20221 12484
rect 20237 12540 20301 12544
rect 20237 12484 20241 12540
rect 20241 12484 20297 12540
rect 20297 12484 20301 12540
rect 20237 12480 20301 12484
rect 20317 12540 20381 12544
rect 20317 12484 20321 12540
rect 20321 12484 20377 12540
rect 20377 12484 20381 12540
rect 20317 12480 20381 12484
rect 20397 12540 20461 12544
rect 20397 12484 20401 12540
rect 20401 12484 20457 12540
rect 20457 12484 20461 12540
rect 20397 12480 20461 12484
rect 27839 12540 27903 12544
rect 27839 12484 27843 12540
rect 27843 12484 27899 12540
rect 27899 12484 27903 12540
rect 27839 12480 27903 12484
rect 27919 12540 27983 12544
rect 27919 12484 27923 12540
rect 27923 12484 27979 12540
rect 27979 12484 27983 12540
rect 27919 12480 27983 12484
rect 27999 12540 28063 12544
rect 27999 12484 28003 12540
rect 28003 12484 28059 12540
rect 28059 12484 28063 12540
rect 27999 12480 28063 12484
rect 28079 12540 28143 12544
rect 28079 12484 28083 12540
rect 28083 12484 28139 12540
rect 28139 12484 28143 12540
rect 28079 12480 28143 12484
rect 17908 12276 17972 12340
rect 18828 12140 18892 12204
rect 25084 12276 25148 12340
rect 19564 12064 19628 12068
rect 19564 12008 19578 12064
rect 19578 12008 19628 12064
rect 19564 12004 19628 12008
rect 24900 12140 24964 12204
rect 8634 11996 8698 12000
rect 8634 11940 8638 11996
rect 8638 11940 8694 11996
rect 8694 11940 8698 11996
rect 8634 11936 8698 11940
rect 8714 11996 8778 12000
rect 8714 11940 8718 11996
rect 8718 11940 8774 11996
rect 8774 11940 8778 11996
rect 8714 11936 8778 11940
rect 8794 11996 8858 12000
rect 8794 11940 8798 11996
rect 8798 11940 8854 11996
rect 8854 11940 8858 11996
rect 8794 11936 8858 11940
rect 8874 11996 8938 12000
rect 8874 11940 8878 11996
rect 8878 11940 8934 11996
rect 8934 11940 8938 11996
rect 8874 11936 8938 11940
rect 16316 11996 16380 12000
rect 16316 11940 16320 11996
rect 16320 11940 16376 11996
rect 16376 11940 16380 11996
rect 16316 11936 16380 11940
rect 16396 11996 16460 12000
rect 16396 11940 16400 11996
rect 16400 11940 16456 11996
rect 16456 11940 16460 11996
rect 16396 11936 16460 11940
rect 16476 11996 16540 12000
rect 16476 11940 16480 11996
rect 16480 11940 16536 11996
rect 16536 11940 16540 11996
rect 16476 11936 16540 11940
rect 16556 11996 16620 12000
rect 16556 11940 16560 11996
rect 16560 11940 16616 11996
rect 16616 11940 16620 11996
rect 16556 11936 16620 11940
rect 23998 11996 24062 12000
rect 23998 11940 24002 11996
rect 24002 11940 24058 11996
rect 24058 11940 24062 11996
rect 23998 11936 24062 11940
rect 24078 11996 24142 12000
rect 24078 11940 24082 11996
rect 24082 11940 24138 11996
rect 24138 11940 24142 11996
rect 24078 11936 24142 11940
rect 24158 11996 24222 12000
rect 24158 11940 24162 11996
rect 24162 11940 24218 11996
rect 24218 11940 24222 11996
rect 24158 11936 24222 11940
rect 24238 11996 24302 12000
rect 24238 11940 24242 11996
rect 24242 11940 24298 11996
rect 24298 11940 24302 11996
rect 24238 11936 24302 11940
rect 31680 11996 31744 12000
rect 31680 11940 31684 11996
rect 31684 11940 31740 11996
rect 31740 11940 31744 11996
rect 31680 11936 31744 11940
rect 31760 11996 31824 12000
rect 31760 11940 31764 11996
rect 31764 11940 31820 11996
rect 31820 11940 31824 11996
rect 31760 11936 31824 11940
rect 31840 11996 31904 12000
rect 31840 11940 31844 11996
rect 31844 11940 31900 11996
rect 31900 11940 31904 11996
rect 31840 11936 31904 11940
rect 31920 11996 31984 12000
rect 31920 11940 31924 11996
rect 31924 11940 31980 11996
rect 31980 11940 31984 11996
rect 31920 11936 31984 11940
rect 24716 11868 24780 11932
rect 26924 11928 26988 11932
rect 26924 11872 26974 11928
rect 26974 11872 26988 11928
rect 26924 11868 26988 11872
rect 20668 11732 20732 11796
rect 4793 11452 4857 11456
rect 4793 11396 4797 11452
rect 4797 11396 4853 11452
rect 4853 11396 4857 11452
rect 4793 11392 4857 11396
rect 4873 11452 4937 11456
rect 4873 11396 4877 11452
rect 4877 11396 4933 11452
rect 4933 11396 4937 11452
rect 4873 11392 4937 11396
rect 4953 11452 5017 11456
rect 4953 11396 4957 11452
rect 4957 11396 5013 11452
rect 5013 11396 5017 11452
rect 4953 11392 5017 11396
rect 5033 11452 5097 11456
rect 5033 11396 5037 11452
rect 5037 11396 5093 11452
rect 5093 11396 5097 11452
rect 5033 11392 5097 11396
rect 12475 11452 12539 11456
rect 12475 11396 12479 11452
rect 12479 11396 12535 11452
rect 12535 11396 12539 11452
rect 12475 11392 12539 11396
rect 12555 11452 12619 11456
rect 12555 11396 12559 11452
rect 12559 11396 12615 11452
rect 12615 11396 12619 11452
rect 12555 11392 12619 11396
rect 12635 11452 12699 11456
rect 12635 11396 12639 11452
rect 12639 11396 12695 11452
rect 12695 11396 12699 11452
rect 12635 11392 12699 11396
rect 12715 11452 12779 11456
rect 12715 11396 12719 11452
rect 12719 11396 12775 11452
rect 12775 11396 12779 11452
rect 12715 11392 12779 11396
rect 20157 11452 20221 11456
rect 20157 11396 20161 11452
rect 20161 11396 20217 11452
rect 20217 11396 20221 11452
rect 20157 11392 20221 11396
rect 20237 11452 20301 11456
rect 20237 11396 20241 11452
rect 20241 11396 20297 11452
rect 20297 11396 20301 11452
rect 20237 11392 20301 11396
rect 20317 11452 20381 11456
rect 20317 11396 20321 11452
rect 20321 11396 20377 11452
rect 20377 11396 20381 11452
rect 20317 11392 20381 11396
rect 20397 11452 20461 11456
rect 20397 11396 20401 11452
rect 20401 11396 20457 11452
rect 20457 11396 20461 11452
rect 20397 11392 20461 11396
rect 27839 11452 27903 11456
rect 27839 11396 27843 11452
rect 27843 11396 27899 11452
rect 27899 11396 27903 11452
rect 27839 11392 27903 11396
rect 27919 11452 27983 11456
rect 27919 11396 27923 11452
rect 27923 11396 27979 11452
rect 27979 11396 27983 11452
rect 27919 11392 27983 11396
rect 27999 11452 28063 11456
rect 27999 11396 28003 11452
rect 28003 11396 28059 11452
rect 28059 11396 28063 11452
rect 27999 11392 28063 11396
rect 28079 11452 28143 11456
rect 28079 11396 28083 11452
rect 28083 11396 28139 11452
rect 28139 11396 28143 11452
rect 28079 11392 28143 11396
rect 26188 11324 26252 11388
rect 28580 11112 28644 11116
rect 28580 11056 28594 11112
rect 28594 11056 28644 11112
rect 28580 11052 28644 11056
rect 27108 10916 27172 10980
rect 31340 10976 31404 10980
rect 31340 10920 31390 10976
rect 31390 10920 31404 10976
rect 31340 10916 31404 10920
rect 8634 10908 8698 10912
rect 8634 10852 8638 10908
rect 8638 10852 8694 10908
rect 8694 10852 8698 10908
rect 8634 10848 8698 10852
rect 8714 10908 8778 10912
rect 8714 10852 8718 10908
rect 8718 10852 8774 10908
rect 8774 10852 8778 10908
rect 8714 10848 8778 10852
rect 8794 10908 8858 10912
rect 8794 10852 8798 10908
rect 8798 10852 8854 10908
rect 8854 10852 8858 10908
rect 8794 10848 8858 10852
rect 8874 10908 8938 10912
rect 8874 10852 8878 10908
rect 8878 10852 8934 10908
rect 8934 10852 8938 10908
rect 8874 10848 8938 10852
rect 16316 10908 16380 10912
rect 16316 10852 16320 10908
rect 16320 10852 16376 10908
rect 16376 10852 16380 10908
rect 16316 10848 16380 10852
rect 16396 10908 16460 10912
rect 16396 10852 16400 10908
rect 16400 10852 16456 10908
rect 16456 10852 16460 10908
rect 16396 10848 16460 10852
rect 16476 10908 16540 10912
rect 16476 10852 16480 10908
rect 16480 10852 16536 10908
rect 16536 10852 16540 10908
rect 16476 10848 16540 10852
rect 16556 10908 16620 10912
rect 16556 10852 16560 10908
rect 16560 10852 16616 10908
rect 16616 10852 16620 10908
rect 16556 10848 16620 10852
rect 23998 10908 24062 10912
rect 23998 10852 24002 10908
rect 24002 10852 24058 10908
rect 24058 10852 24062 10908
rect 23998 10848 24062 10852
rect 24078 10908 24142 10912
rect 24078 10852 24082 10908
rect 24082 10852 24138 10908
rect 24138 10852 24142 10908
rect 24078 10848 24142 10852
rect 24158 10908 24222 10912
rect 24158 10852 24162 10908
rect 24162 10852 24218 10908
rect 24218 10852 24222 10908
rect 24158 10848 24222 10852
rect 24238 10908 24302 10912
rect 24238 10852 24242 10908
rect 24242 10852 24298 10908
rect 24298 10852 24302 10908
rect 24238 10848 24302 10852
rect 31680 10908 31744 10912
rect 31680 10852 31684 10908
rect 31684 10852 31740 10908
rect 31740 10852 31744 10908
rect 31680 10848 31744 10852
rect 31760 10908 31824 10912
rect 31760 10852 31764 10908
rect 31764 10852 31820 10908
rect 31820 10852 31824 10908
rect 31760 10848 31824 10852
rect 31840 10908 31904 10912
rect 31840 10852 31844 10908
rect 31844 10852 31900 10908
rect 31900 10852 31904 10908
rect 31840 10848 31904 10852
rect 31920 10908 31984 10912
rect 31920 10852 31924 10908
rect 31924 10852 31980 10908
rect 31980 10852 31984 10908
rect 31920 10848 31984 10852
rect 30420 10780 30484 10844
rect 20852 10704 20916 10708
rect 20852 10648 20902 10704
rect 20902 10648 20916 10704
rect 20852 10644 20916 10648
rect 23612 10644 23676 10708
rect 10548 10508 10612 10572
rect 4793 10364 4857 10368
rect 4793 10308 4797 10364
rect 4797 10308 4853 10364
rect 4853 10308 4857 10364
rect 4793 10304 4857 10308
rect 4873 10364 4937 10368
rect 4873 10308 4877 10364
rect 4877 10308 4933 10364
rect 4933 10308 4937 10364
rect 4873 10304 4937 10308
rect 4953 10364 5017 10368
rect 4953 10308 4957 10364
rect 4957 10308 5013 10364
rect 5013 10308 5017 10364
rect 4953 10304 5017 10308
rect 5033 10364 5097 10368
rect 5033 10308 5037 10364
rect 5037 10308 5093 10364
rect 5093 10308 5097 10364
rect 5033 10304 5097 10308
rect 12475 10364 12539 10368
rect 12475 10308 12479 10364
rect 12479 10308 12535 10364
rect 12535 10308 12539 10364
rect 12475 10304 12539 10308
rect 12555 10364 12619 10368
rect 12555 10308 12559 10364
rect 12559 10308 12615 10364
rect 12615 10308 12619 10364
rect 12555 10304 12619 10308
rect 12635 10364 12699 10368
rect 12635 10308 12639 10364
rect 12639 10308 12695 10364
rect 12695 10308 12699 10364
rect 12635 10304 12699 10308
rect 12715 10364 12779 10368
rect 12715 10308 12719 10364
rect 12719 10308 12775 10364
rect 12775 10308 12779 10364
rect 12715 10304 12779 10308
rect 20157 10364 20221 10368
rect 20157 10308 20161 10364
rect 20161 10308 20217 10364
rect 20217 10308 20221 10364
rect 20157 10304 20221 10308
rect 20237 10364 20301 10368
rect 20237 10308 20241 10364
rect 20241 10308 20297 10364
rect 20297 10308 20301 10364
rect 20237 10304 20301 10308
rect 20317 10364 20381 10368
rect 20317 10308 20321 10364
rect 20321 10308 20377 10364
rect 20377 10308 20381 10364
rect 20317 10304 20381 10308
rect 20397 10364 20461 10368
rect 20397 10308 20401 10364
rect 20401 10308 20457 10364
rect 20457 10308 20461 10364
rect 20397 10304 20461 10308
rect 27839 10364 27903 10368
rect 27839 10308 27843 10364
rect 27843 10308 27899 10364
rect 27899 10308 27903 10364
rect 27839 10304 27903 10308
rect 27919 10364 27983 10368
rect 27919 10308 27923 10364
rect 27923 10308 27979 10364
rect 27979 10308 27983 10364
rect 27919 10304 27983 10308
rect 27999 10364 28063 10368
rect 27999 10308 28003 10364
rect 28003 10308 28059 10364
rect 28059 10308 28063 10364
rect 27999 10304 28063 10308
rect 28079 10364 28143 10368
rect 28079 10308 28083 10364
rect 28083 10308 28139 10364
rect 28139 10308 28143 10364
rect 28079 10304 28143 10308
rect 6500 10100 6564 10164
rect 15884 9964 15948 10028
rect 8634 9820 8698 9824
rect 8634 9764 8638 9820
rect 8638 9764 8694 9820
rect 8694 9764 8698 9820
rect 8634 9760 8698 9764
rect 8714 9820 8778 9824
rect 8714 9764 8718 9820
rect 8718 9764 8774 9820
rect 8774 9764 8778 9820
rect 8714 9760 8778 9764
rect 8794 9820 8858 9824
rect 8794 9764 8798 9820
rect 8798 9764 8854 9820
rect 8854 9764 8858 9820
rect 8794 9760 8858 9764
rect 8874 9820 8938 9824
rect 8874 9764 8878 9820
rect 8878 9764 8934 9820
rect 8934 9764 8938 9820
rect 8874 9760 8938 9764
rect 16316 9820 16380 9824
rect 16316 9764 16320 9820
rect 16320 9764 16376 9820
rect 16376 9764 16380 9820
rect 16316 9760 16380 9764
rect 16396 9820 16460 9824
rect 16396 9764 16400 9820
rect 16400 9764 16456 9820
rect 16456 9764 16460 9820
rect 16396 9760 16460 9764
rect 16476 9820 16540 9824
rect 16476 9764 16480 9820
rect 16480 9764 16536 9820
rect 16536 9764 16540 9820
rect 16476 9760 16540 9764
rect 16556 9820 16620 9824
rect 16556 9764 16560 9820
rect 16560 9764 16616 9820
rect 16616 9764 16620 9820
rect 16556 9760 16620 9764
rect 23998 9820 24062 9824
rect 23998 9764 24002 9820
rect 24002 9764 24058 9820
rect 24058 9764 24062 9820
rect 23998 9760 24062 9764
rect 24078 9820 24142 9824
rect 24078 9764 24082 9820
rect 24082 9764 24138 9820
rect 24138 9764 24142 9820
rect 24078 9760 24142 9764
rect 24158 9820 24222 9824
rect 24158 9764 24162 9820
rect 24162 9764 24218 9820
rect 24218 9764 24222 9820
rect 24158 9760 24222 9764
rect 24238 9820 24302 9824
rect 24238 9764 24242 9820
rect 24242 9764 24298 9820
rect 24298 9764 24302 9820
rect 24238 9760 24302 9764
rect 31680 9820 31744 9824
rect 31680 9764 31684 9820
rect 31684 9764 31740 9820
rect 31740 9764 31744 9820
rect 31680 9760 31744 9764
rect 31760 9820 31824 9824
rect 31760 9764 31764 9820
rect 31764 9764 31820 9820
rect 31820 9764 31824 9820
rect 31760 9760 31824 9764
rect 31840 9820 31904 9824
rect 31840 9764 31844 9820
rect 31844 9764 31900 9820
rect 31900 9764 31904 9820
rect 31840 9760 31904 9764
rect 31920 9820 31984 9824
rect 31920 9764 31924 9820
rect 31924 9764 31980 9820
rect 31980 9764 31984 9820
rect 31920 9760 31984 9764
rect 27108 9692 27172 9756
rect 5396 9616 5460 9620
rect 5396 9560 5446 9616
rect 5446 9560 5460 9616
rect 5396 9556 5460 9560
rect 25820 9556 25884 9620
rect 26740 9284 26804 9348
rect 4793 9276 4857 9280
rect 4793 9220 4797 9276
rect 4797 9220 4853 9276
rect 4853 9220 4857 9276
rect 4793 9216 4857 9220
rect 4873 9276 4937 9280
rect 4873 9220 4877 9276
rect 4877 9220 4933 9276
rect 4933 9220 4937 9276
rect 4873 9216 4937 9220
rect 4953 9276 5017 9280
rect 4953 9220 4957 9276
rect 4957 9220 5013 9276
rect 5013 9220 5017 9276
rect 4953 9216 5017 9220
rect 5033 9276 5097 9280
rect 5033 9220 5037 9276
rect 5037 9220 5093 9276
rect 5093 9220 5097 9276
rect 5033 9216 5097 9220
rect 12475 9276 12539 9280
rect 12475 9220 12479 9276
rect 12479 9220 12535 9276
rect 12535 9220 12539 9276
rect 12475 9216 12539 9220
rect 12555 9276 12619 9280
rect 12555 9220 12559 9276
rect 12559 9220 12615 9276
rect 12615 9220 12619 9276
rect 12555 9216 12619 9220
rect 12635 9276 12699 9280
rect 12635 9220 12639 9276
rect 12639 9220 12695 9276
rect 12695 9220 12699 9276
rect 12635 9216 12699 9220
rect 12715 9276 12779 9280
rect 12715 9220 12719 9276
rect 12719 9220 12775 9276
rect 12775 9220 12779 9276
rect 12715 9216 12779 9220
rect 20157 9276 20221 9280
rect 20157 9220 20161 9276
rect 20161 9220 20217 9276
rect 20217 9220 20221 9276
rect 20157 9216 20221 9220
rect 20237 9276 20301 9280
rect 20237 9220 20241 9276
rect 20241 9220 20297 9276
rect 20297 9220 20301 9276
rect 20237 9216 20301 9220
rect 20317 9276 20381 9280
rect 20317 9220 20321 9276
rect 20321 9220 20377 9276
rect 20377 9220 20381 9276
rect 20317 9216 20381 9220
rect 20397 9276 20461 9280
rect 20397 9220 20401 9276
rect 20401 9220 20457 9276
rect 20457 9220 20461 9276
rect 20397 9216 20461 9220
rect 27839 9276 27903 9280
rect 27839 9220 27843 9276
rect 27843 9220 27899 9276
rect 27899 9220 27903 9276
rect 27839 9216 27903 9220
rect 27919 9276 27983 9280
rect 27919 9220 27923 9276
rect 27923 9220 27979 9276
rect 27979 9220 27983 9276
rect 27919 9216 27983 9220
rect 27999 9276 28063 9280
rect 27999 9220 28003 9276
rect 28003 9220 28059 9276
rect 28059 9220 28063 9276
rect 27999 9216 28063 9220
rect 28079 9276 28143 9280
rect 28079 9220 28083 9276
rect 28083 9220 28139 9276
rect 28139 9220 28143 9276
rect 28079 9216 28143 9220
rect 13308 9012 13372 9076
rect 15332 8876 15396 8940
rect 28948 8740 29012 8804
rect 8634 8732 8698 8736
rect 8634 8676 8638 8732
rect 8638 8676 8694 8732
rect 8694 8676 8698 8732
rect 8634 8672 8698 8676
rect 8714 8732 8778 8736
rect 8714 8676 8718 8732
rect 8718 8676 8774 8732
rect 8774 8676 8778 8732
rect 8714 8672 8778 8676
rect 8794 8732 8858 8736
rect 8794 8676 8798 8732
rect 8798 8676 8854 8732
rect 8854 8676 8858 8732
rect 8794 8672 8858 8676
rect 8874 8732 8938 8736
rect 8874 8676 8878 8732
rect 8878 8676 8934 8732
rect 8934 8676 8938 8732
rect 8874 8672 8938 8676
rect 16316 8732 16380 8736
rect 16316 8676 16320 8732
rect 16320 8676 16376 8732
rect 16376 8676 16380 8732
rect 16316 8672 16380 8676
rect 16396 8732 16460 8736
rect 16396 8676 16400 8732
rect 16400 8676 16456 8732
rect 16456 8676 16460 8732
rect 16396 8672 16460 8676
rect 16476 8732 16540 8736
rect 16476 8676 16480 8732
rect 16480 8676 16536 8732
rect 16536 8676 16540 8732
rect 16476 8672 16540 8676
rect 16556 8732 16620 8736
rect 16556 8676 16560 8732
rect 16560 8676 16616 8732
rect 16616 8676 16620 8732
rect 16556 8672 16620 8676
rect 23998 8732 24062 8736
rect 23998 8676 24002 8732
rect 24002 8676 24058 8732
rect 24058 8676 24062 8732
rect 23998 8672 24062 8676
rect 24078 8732 24142 8736
rect 24078 8676 24082 8732
rect 24082 8676 24138 8732
rect 24138 8676 24142 8732
rect 24078 8672 24142 8676
rect 24158 8732 24222 8736
rect 24158 8676 24162 8732
rect 24162 8676 24218 8732
rect 24218 8676 24222 8732
rect 24158 8672 24222 8676
rect 24238 8732 24302 8736
rect 24238 8676 24242 8732
rect 24242 8676 24298 8732
rect 24298 8676 24302 8732
rect 24238 8672 24302 8676
rect 31680 8732 31744 8736
rect 31680 8676 31684 8732
rect 31684 8676 31740 8732
rect 31740 8676 31744 8732
rect 31680 8672 31744 8676
rect 31760 8732 31824 8736
rect 31760 8676 31764 8732
rect 31764 8676 31820 8732
rect 31820 8676 31824 8732
rect 31760 8672 31824 8676
rect 31840 8732 31904 8736
rect 31840 8676 31844 8732
rect 31844 8676 31900 8732
rect 31900 8676 31904 8732
rect 31840 8672 31904 8676
rect 31920 8732 31984 8736
rect 31920 8676 31924 8732
rect 31924 8676 31980 8732
rect 31980 8676 31984 8732
rect 31920 8672 31984 8676
rect 17724 8604 17788 8668
rect 29684 8664 29748 8668
rect 29684 8608 29734 8664
rect 29734 8608 29748 8664
rect 29684 8604 29748 8608
rect 30052 8604 30116 8668
rect 13124 8468 13188 8532
rect 19380 8332 19444 8396
rect 4793 8188 4857 8192
rect 4793 8132 4797 8188
rect 4797 8132 4853 8188
rect 4853 8132 4857 8188
rect 4793 8128 4857 8132
rect 4873 8188 4937 8192
rect 4873 8132 4877 8188
rect 4877 8132 4933 8188
rect 4933 8132 4937 8188
rect 4873 8128 4937 8132
rect 4953 8188 5017 8192
rect 4953 8132 4957 8188
rect 4957 8132 5013 8188
rect 5013 8132 5017 8188
rect 4953 8128 5017 8132
rect 5033 8188 5097 8192
rect 5033 8132 5037 8188
rect 5037 8132 5093 8188
rect 5093 8132 5097 8188
rect 5033 8128 5097 8132
rect 12475 8188 12539 8192
rect 12475 8132 12479 8188
rect 12479 8132 12535 8188
rect 12535 8132 12539 8188
rect 12475 8128 12539 8132
rect 12555 8188 12619 8192
rect 12555 8132 12559 8188
rect 12559 8132 12615 8188
rect 12615 8132 12619 8188
rect 12555 8128 12619 8132
rect 12635 8188 12699 8192
rect 12635 8132 12639 8188
rect 12639 8132 12695 8188
rect 12695 8132 12699 8188
rect 12635 8128 12699 8132
rect 12715 8188 12779 8192
rect 12715 8132 12719 8188
rect 12719 8132 12775 8188
rect 12775 8132 12779 8188
rect 12715 8128 12779 8132
rect 20157 8188 20221 8192
rect 20157 8132 20161 8188
rect 20161 8132 20217 8188
rect 20217 8132 20221 8188
rect 20157 8128 20221 8132
rect 20237 8188 20301 8192
rect 20237 8132 20241 8188
rect 20241 8132 20297 8188
rect 20297 8132 20301 8188
rect 20237 8128 20301 8132
rect 20317 8188 20381 8192
rect 20317 8132 20321 8188
rect 20321 8132 20377 8188
rect 20377 8132 20381 8188
rect 20317 8128 20381 8132
rect 20397 8188 20461 8192
rect 20397 8132 20401 8188
rect 20401 8132 20457 8188
rect 20457 8132 20461 8188
rect 20397 8128 20461 8132
rect 27839 8188 27903 8192
rect 27839 8132 27843 8188
rect 27843 8132 27899 8188
rect 27899 8132 27903 8188
rect 27839 8128 27903 8132
rect 27919 8188 27983 8192
rect 27919 8132 27923 8188
rect 27923 8132 27979 8188
rect 27979 8132 27983 8188
rect 27919 8128 27983 8132
rect 27999 8188 28063 8192
rect 27999 8132 28003 8188
rect 28003 8132 28059 8188
rect 28059 8132 28063 8188
rect 27999 8128 28063 8132
rect 28079 8188 28143 8192
rect 28079 8132 28083 8188
rect 28083 8132 28139 8188
rect 28139 8132 28143 8188
rect 28079 8128 28143 8132
rect 21036 7924 21100 7988
rect 9444 7788 9508 7852
rect 8634 7644 8698 7648
rect 8634 7588 8638 7644
rect 8638 7588 8694 7644
rect 8694 7588 8698 7644
rect 8634 7584 8698 7588
rect 8714 7644 8778 7648
rect 8714 7588 8718 7644
rect 8718 7588 8774 7644
rect 8774 7588 8778 7644
rect 8714 7584 8778 7588
rect 8794 7644 8858 7648
rect 8794 7588 8798 7644
rect 8798 7588 8854 7644
rect 8854 7588 8858 7644
rect 8794 7584 8858 7588
rect 8874 7644 8938 7648
rect 8874 7588 8878 7644
rect 8878 7588 8934 7644
rect 8934 7588 8938 7644
rect 8874 7584 8938 7588
rect 16316 7644 16380 7648
rect 16316 7588 16320 7644
rect 16320 7588 16376 7644
rect 16376 7588 16380 7644
rect 16316 7584 16380 7588
rect 16396 7644 16460 7648
rect 16396 7588 16400 7644
rect 16400 7588 16456 7644
rect 16456 7588 16460 7644
rect 16396 7584 16460 7588
rect 16476 7644 16540 7648
rect 16476 7588 16480 7644
rect 16480 7588 16536 7644
rect 16536 7588 16540 7644
rect 16476 7584 16540 7588
rect 16556 7644 16620 7648
rect 16556 7588 16560 7644
rect 16560 7588 16616 7644
rect 16616 7588 16620 7644
rect 16556 7584 16620 7588
rect 23998 7644 24062 7648
rect 23998 7588 24002 7644
rect 24002 7588 24058 7644
rect 24058 7588 24062 7644
rect 23998 7584 24062 7588
rect 24078 7644 24142 7648
rect 24078 7588 24082 7644
rect 24082 7588 24138 7644
rect 24138 7588 24142 7644
rect 24078 7584 24142 7588
rect 24158 7644 24222 7648
rect 24158 7588 24162 7644
rect 24162 7588 24218 7644
rect 24218 7588 24222 7644
rect 24158 7584 24222 7588
rect 24238 7644 24302 7648
rect 24238 7588 24242 7644
rect 24242 7588 24298 7644
rect 24298 7588 24302 7644
rect 24238 7584 24302 7588
rect 31680 7644 31744 7648
rect 31680 7588 31684 7644
rect 31684 7588 31740 7644
rect 31740 7588 31744 7644
rect 31680 7584 31744 7588
rect 31760 7644 31824 7648
rect 31760 7588 31764 7644
rect 31764 7588 31820 7644
rect 31820 7588 31824 7644
rect 31760 7584 31824 7588
rect 31840 7644 31904 7648
rect 31840 7588 31844 7644
rect 31844 7588 31900 7644
rect 31900 7588 31904 7644
rect 31840 7584 31904 7588
rect 31920 7644 31984 7648
rect 31920 7588 31924 7644
rect 31924 7588 31980 7644
rect 31980 7588 31984 7644
rect 31920 7584 31984 7588
rect 14412 7380 14476 7444
rect 11836 7244 11900 7308
rect 4793 7100 4857 7104
rect 4793 7044 4797 7100
rect 4797 7044 4853 7100
rect 4853 7044 4857 7100
rect 4793 7040 4857 7044
rect 4873 7100 4937 7104
rect 4873 7044 4877 7100
rect 4877 7044 4933 7100
rect 4933 7044 4937 7100
rect 4873 7040 4937 7044
rect 4953 7100 5017 7104
rect 4953 7044 4957 7100
rect 4957 7044 5013 7100
rect 5013 7044 5017 7100
rect 4953 7040 5017 7044
rect 5033 7100 5097 7104
rect 5033 7044 5037 7100
rect 5037 7044 5093 7100
rect 5093 7044 5097 7100
rect 5033 7040 5097 7044
rect 12475 7100 12539 7104
rect 12475 7044 12479 7100
rect 12479 7044 12535 7100
rect 12535 7044 12539 7100
rect 12475 7040 12539 7044
rect 12555 7100 12619 7104
rect 12555 7044 12559 7100
rect 12559 7044 12615 7100
rect 12615 7044 12619 7100
rect 12555 7040 12619 7044
rect 12635 7100 12699 7104
rect 12635 7044 12639 7100
rect 12639 7044 12695 7100
rect 12695 7044 12699 7100
rect 12635 7040 12699 7044
rect 12715 7100 12779 7104
rect 12715 7044 12719 7100
rect 12719 7044 12775 7100
rect 12775 7044 12779 7100
rect 12715 7040 12779 7044
rect 20157 7100 20221 7104
rect 20157 7044 20161 7100
rect 20161 7044 20217 7100
rect 20217 7044 20221 7100
rect 20157 7040 20221 7044
rect 20237 7100 20301 7104
rect 20237 7044 20241 7100
rect 20241 7044 20297 7100
rect 20297 7044 20301 7100
rect 20237 7040 20301 7044
rect 20317 7100 20381 7104
rect 20317 7044 20321 7100
rect 20321 7044 20377 7100
rect 20377 7044 20381 7100
rect 20317 7040 20381 7044
rect 20397 7100 20461 7104
rect 20397 7044 20401 7100
rect 20401 7044 20457 7100
rect 20457 7044 20461 7100
rect 20397 7040 20461 7044
rect 27839 7100 27903 7104
rect 27839 7044 27843 7100
rect 27843 7044 27899 7100
rect 27899 7044 27903 7100
rect 27839 7040 27903 7044
rect 27919 7100 27983 7104
rect 27919 7044 27923 7100
rect 27923 7044 27979 7100
rect 27979 7044 27983 7100
rect 27919 7040 27983 7044
rect 27999 7100 28063 7104
rect 27999 7044 28003 7100
rect 28003 7044 28059 7100
rect 28059 7044 28063 7100
rect 27999 7040 28063 7044
rect 28079 7100 28143 7104
rect 28079 7044 28083 7100
rect 28083 7044 28139 7100
rect 28139 7044 28143 7100
rect 28079 7040 28143 7044
rect 14044 6836 14108 6900
rect 18644 6700 18708 6764
rect 8634 6556 8698 6560
rect 8634 6500 8638 6556
rect 8638 6500 8694 6556
rect 8694 6500 8698 6556
rect 8634 6496 8698 6500
rect 8714 6556 8778 6560
rect 8714 6500 8718 6556
rect 8718 6500 8774 6556
rect 8774 6500 8778 6556
rect 8714 6496 8778 6500
rect 8794 6556 8858 6560
rect 8794 6500 8798 6556
rect 8798 6500 8854 6556
rect 8854 6500 8858 6556
rect 8794 6496 8858 6500
rect 8874 6556 8938 6560
rect 8874 6500 8878 6556
rect 8878 6500 8934 6556
rect 8934 6500 8938 6556
rect 8874 6496 8938 6500
rect 16316 6556 16380 6560
rect 16316 6500 16320 6556
rect 16320 6500 16376 6556
rect 16376 6500 16380 6556
rect 16316 6496 16380 6500
rect 16396 6556 16460 6560
rect 16396 6500 16400 6556
rect 16400 6500 16456 6556
rect 16456 6500 16460 6556
rect 16396 6496 16460 6500
rect 16476 6556 16540 6560
rect 16476 6500 16480 6556
rect 16480 6500 16536 6556
rect 16536 6500 16540 6556
rect 16476 6496 16540 6500
rect 16556 6556 16620 6560
rect 16556 6500 16560 6556
rect 16560 6500 16616 6556
rect 16616 6500 16620 6556
rect 16556 6496 16620 6500
rect 23998 6556 24062 6560
rect 23998 6500 24002 6556
rect 24002 6500 24058 6556
rect 24058 6500 24062 6556
rect 23998 6496 24062 6500
rect 24078 6556 24142 6560
rect 24078 6500 24082 6556
rect 24082 6500 24138 6556
rect 24138 6500 24142 6556
rect 24078 6496 24142 6500
rect 24158 6556 24222 6560
rect 24158 6500 24162 6556
rect 24162 6500 24218 6556
rect 24218 6500 24222 6556
rect 24158 6496 24222 6500
rect 24238 6556 24302 6560
rect 24238 6500 24242 6556
rect 24242 6500 24298 6556
rect 24298 6500 24302 6556
rect 24238 6496 24302 6500
rect 31680 6556 31744 6560
rect 31680 6500 31684 6556
rect 31684 6500 31740 6556
rect 31740 6500 31744 6556
rect 31680 6496 31744 6500
rect 31760 6556 31824 6560
rect 31760 6500 31764 6556
rect 31764 6500 31820 6556
rect 31820 6500 31824 6556
rect 31760 6496 31824 6500
rect 31840 6556 31904 6560
rect 31840 6500 31844 6556
rect 31844 6500 31900 6556
rect 31900 6500 31904 6556
rect 31840 6496 31904 6500
rect 31920 6556 31984 6560
rect 31920 6500 31924 6556
rect 31924 6500 31980 6556
rect 31980 6500 31984 6556
rect 31920 6496 31984 6500
rect 28764 6216 28828 6220
rect 28764 6160 28778 6216
rect 28778 6160 28828 6216
rect 28764 6156 28828 6160
rect 4793 6012 4857 6016
rect 4793 5956 4797 6012
rect 4797 5956 4853 6012
rect 4853 5956 4857 6012
rect 4793 5952 4857 5956
rect 4873 6012 4937 6016
rect 4873 5956 4877 6012
rect 4877 5956 4933 6012
rect 4933 5956 4937 6012
rect 4873 5952 4937 5956
rect 4953 6012 5017 6016
rect 4953 5956 4957 6012
rect 4957 5956 5013 6012
rect 5013 5956 5017 6012
rect 4953 5952 5017 5956
rect 5033 6012 5097 6016
rect 5033 5956 5037 6012
rect 5037 5956 5093 6012
rect 5093 5956 5097 6012
rect 5033 5952 5097 5956
rect 12475 6012 12539 6016
rect 12475 5956 12479 6012
rect 12479 5956 12535 6012
rect 12535 5956 12539 6012
rect 12475 5952 12539 5956
rect 12555 6012 12619 6016
rect 12555 5956 12559 6012
rect 12559 5956 12615 6012
rect 12615 5956 12619 6012
rect 12555 5952 12619 5956
rect 12635 6012 12699 6016
rect 12635 5956 12639 6012
rect 12639 5956 12695 6012
rect 12695 5956 12699 6012
rect 12635 5952 12699 5956
rect 12715 6012 12779 6016
rect 12715 5956 12719 6012
rect 12719 5956 12775 6012
rect 12775 5956 12779 6012
rect 12715 5952 12779 5956
rect 20157 6012 20221 6016
rect 20157 5956 20161 6012
rect 20161 5956 20217 6012
rect 20217 5956 20221 6012
rect 20157 5952 20221 5956
rect 20237 6012 20301 6016
rect 20237 5956 20241 6012
rect 20241 5956 20297 6012
rect 20297 5956 20301 6012
rect 20237 5952 20301 5956
rect 20317 6012 20381 6016
rect 20317 5956 20321 6012
rect 20321 5956 20377 6012
rect 20377 5956 20381 6012
rect 20317 5952 20381 5956
rect 20397 6012 20461 6016
rect 20397 5956 20401 6012
rect 20401 5956 20457 6012
rect 20457 5956 20461 6012
rect 20397 5952 20461 5956
rect 27839 6012 27903 6016
rect 27839 5956 27843 6012
rect 27843 5956 27899 6012
rect 27899 5956 27903 6012
rect 27839 5952 27903 5956
rect 27919 6012 27983 6016
rect 27919 5956 27923 6012
rect 27923 5956 27979 6012
rect 27979 5956 27983 6012
rect 27919 5952 27983 5956
rect 27999 6012 28063 6016
rect 27999 5956 28003 6012
rect 28003 5956 28059 6012
rect 28059 5956 28063 6012
rect 27999 5952 28063 5956
rect 28079 6012 28143 6016
rect 28079 5956 28083 6012
rect 28083 5956 28139 6012
rect 28139 5956 28143 6012
rect 28079 5952 28143 5956
rect 8634 5468 8698 5472
rect 8634 5412 8638 5468
rect 8638 5412 8694 5468
rect 8694 5412 8698 5468
rect 8634 5408 8698 5412
rect 8714 5468 8778 5472
rect 8714 5412 8718 5468
rect 8718 5412 8774 5468
rect 8774 5412 8778 5468
rect 8714 5408 8778 5412
rect 8794 5468 8858 5472
rect 8794 5412 8798 5468
rect 8798 5412 8854 5468
rect 8854 5412 8858 5468
rect 8794 5408 8858 5412
rect 8874 5468 8938 5472
rect 8874 5412 8878 5468
rect 8878 5412 8934 5468
rect 8934 5412 8938 5468
rect 8874 5408 8938 5412
rect 16316 5468 16380 5472
rect 16316 5412 16320 5468
rect 16320 5412 16376 5468
rect 16376 5412 16380 5468
rect 16316 5408 16380 5412
rect 16396 5468 16460 5472
rect 16396 5412 16400 5468
rect 16400 5412 16456 5468
rect 16456 5412 16460 5468
rect 16396 5408 16460 5412
rect 16476 5468 16540 5472
rect 16476 5412 16480 5468
rect 16480 5412 16536 5468
rect 16536 5412 16540 5468
rect 16476 5408 16540 5412
rect 16556 5468 16620 5472
rect 16556 5412 16560 5468
rect 16560 5412 16616 5468
rect 16616 5412 16620 5468
rect 16556 5408 16620 5412
rect 23998 5468 24062 5472
rect 23998 5412 24002 5468
rect 24002 5412 24058 5468
rect 24058 5412 24062 5468
rect 23998 5408 24062 5412
rect 24078 5468 24142 5472
rect 24078 5412 24082 5468
rect 24082 5412 24138 5468
rect 24138 5412 24142 5468
rect 24078 5408 24142 5412
rect 24158 5468 24222 5472
rect 24158 5412 24162 5468
rect 24162 5412 24218 5468
rect 24218 5412 24222 5468
rect 24158 5408 24222 5412
rect 24238 5468 24302 5472
rect 24238 5412 24242 5468
rect 24242 5412 24298 5468
rect 24298 5412 24302 5468
rect 24238 5408 24302 5412
rect 31680 5468 31744 5472
rect 31680 5412 31684 5468
rect 31684 5412 31740 5468
rect 31740 5412 31744 5468
rect 31680 5408 31744 5412
rect 31760 5468 31824 5472
rect 31760 5412 31764 5468
rect 31764 5412 31820 5468
rect 31820 5412 31824 5468
rect 31760 5408 31824 5412
rect 31840 5468 31904 5472
rect 31840 5412 31844 5468
rect 31844 5412 31900 5468
rect 31900 5412 31904 5468
rect 31840 5408 31904 5412
rect 31920 5468 31984 5472
rect 31920 5412 31924 5468
rect 31924 5412 31980 5468
rect 31980 5412 31984 5468
rect 31920 5408 31984 5412
rect 28948 5204 29012 5268
rect 13492 5068 13556 5132
rect 4793 4924 4857 4928
rect 4793 4868 4797 4924
rect 4797 4868 4853 4924
rect 4853 4868 4857 4924
rect 4793 4864 4857 4868
rect 4873 4924 4937 4928
rect 4873 4868 4877 4924
rect 4877 4868 4933 4924
rect 4933 4868 4937 4924
rect 4873 4864 4937 4868
rect 4953 4924 5017 4928
rect 4953 4868 4957 4924
rect 4957 4868 5013 4924
rect 5013 4868 5017 4924
rect 4953 4864 5017 4868
rect 5033 4924 5097 4928
rect 5033 4868 5037 4924
rect 5037 4868 5093 4924
rect 5093 4868 5097 4924
rect 5033 4864 5097 4868
rect 12475 4924 12539 4928
rect 12475 4868 12479 4924
rect 12479 4868 12535 4924
rect 12535 4868 12539 4924
rect 12475 4864 12539 4868
rect 12555 4924 12619 4928
rect 12555 4868 12559 4924
rect 12559 4868 12615 4924
rect 12615 4868 12619 4924
rect 12555 4864 12619 4868
rect 12635 4924 12699 4928
rect 12635 4868 12639 4924
rect 12639 4868 12695 4924
rect 12695 4868 12699 4924
rect 12635 4864 12699 4868
rect 12715 4924 12779 4928
rect 12715 4868 12719 4924
rect 12719 4868 12775 4924
rect 12775 4868 12779 4924
rect 12715 4864 12779 4868
rect 20157 4924 20221 4928
rect 20157 4868 20161 4924
rect 20161 4868 20217 4924
rect 20217 4868 20221 4924
rect 20157 4864 20221 4868
rect 20237 4924 20301 4928
rect 20237 4868 20241 4924
rect 20241 4868 20297 4924
rect 20297 4868 20301 4924
rect 20237 4864 20301 4868
rect 20317 4924 20381 4928
rect 20317 4868 20321 4924
rect 20321 4868 20377 4924
rect 20377 4868 20381 4924
rect 20317 4864 20381 4868
rect 20397 4924 20461 4928
rect 20397 4868 20401 4924
rect 20401 4868 20457 4924
rect 20457 4868 20461 4924
rect 20397 4864 20461 4868
rect 27839 4924 27903 4928
rect 27839 4868 27843 4924
rect 27843 4868 27899 4924
rect 27899 4868 27903 4924
rect 27839 4864 27903 4868
rect 27919 4924 27983 4928
rect 27919 4868 27923 4924
rect 27923 4868 27979 4924
rect 27979 4868 27983 4924
rect 27919 4864 27983 4868
rect 27999 4924 28063 4928
rect 27999 4868 28003 4924
rect 28003 4868 28059 4924
rect 28059 4868 28063 4924
rect 27999 4864 28063 4868
rect 28079 4924 28143 4928
rect 28079 4868 28083 4924
rect 28083 4868 28139 4924
rect 28139 4868 28143 4924
rect 28079 4864 28143 4868
rect 15700 4660 15764 4724
rect 29684 4660 29748 4724
rect 8634 4380 8698 4384
rect 8634 4324 8638 4380
rect 8638 4324 8694 4380
rect 8694 4324 8698 4380
rect 8634 4320 8698 4324
rect 8714 4380 8778 4384
rect 8714 4324 8718 4380
rect 8718 4324 8774 4380
rect 8774 4324 8778 4380
rect 8714 4320 8778 4324
rect 8794 4380 8858 4384
rect 8794 4324 8798 4380
rect 8798 4324 8854 4380
rect 8854 4324 8858 4380
rect 8794 4320 8858 4324
rect 8874 4380 8938 4384
rect 8874 4324 8878 4380
rect 8878 4324 8934 4380
rect 8934 4324 8938 4380
rect 8874 4320 8938 4324
rect 16316 4380 16380 4384
rect 16316 4324 16320 4380
rect 16320 4324 16376 4380
rect 16376 4324 16380 4380
rect 16316 4320 16380 4324
rect 16396 4380 16460 4384
rect 16396 4324 16400 4380
rect 16400 4324 16456 4380
rect 16456 4324 16460 4380
rect 16396 4320 16460 4324
rect 16476 4380 16540 4384
rect 16476 4324 16480 4380
rect 16480 4324 16536 4380
rect 16536 4324 16540 4380
rect 16476 4320 16540 4324
rect 16556 4380 16620 4384
rect 16556 4324 16560 4380
rect 16560 4324 16616 4380
rect 16616 4324 16620 4380
rect 16556 4320 16620 4324
rect 23998 4380 24062 4384
rect 23998 4324 24002 4380
rect 24002 4324 24058 4380
rect 24058 4324 24062 4380
rect 23998 4320 24062 4324
rect 24078 4380 24142 4384
rect 24078 4324 24082 4380
rect 24082 4324 24138 4380
rect 24138 4324 24142 4380
rect 24078 4320 24142 4324
rect 24158 4380 24222 4384
rect 24158 4324 24162 4380
rect 24162 4324 24218 4380
rect 24218 4324 24222 4380
rect 24158 4320 24222 4324
rect 24238 4380 24302 4384
rect 24238 4324 24242 4380
rect 24242 4324 24298 4380
rect 24298 4324 24302 4380
rect 24238 4320 24302 4324
rect 31680 4380 31744 4384
rect 31680 4324 31684 4380
rect 31684 4324 31740 4380
rect 31740 4324 31744 4380
rect 31680 4320 31744 4324
rect 31760 4380 31824 4384
rect 31760 4324 31764 4380
rect 31764 4324 31820 4380
rect 31820 4324 31824 4380
rect 31760 4320 31824 4324
rect 31840 4380 31904 4384
rect 31840 4324 31844 4380
rect 31844 4324 31900 4380
rect 31900 4324 31904 4380
rect 31840 4320 31904 4324
rect 31920 4380 31984 4384
rect 31920 4324 31924 4380
rect 31924 4324 31980 4380
rect 31980 4324 31984 4380
rect 31920 4320 31984 4324
rect 4793 3836 4857 3840
rect 4793 3780 4797 3836
rect 4797 3780 4853 3836
rect 4853 3780 4857 3836
rect 4793 3776 4857 3780
rect 4873 3836 4937 3840
rect 4873 3780 4877 3836
rect 4877 3780 4933 3836
rect 4933 3780 4937 3836
rect 4873 3776 4937 3780
rect 4953 3836 5017 3840
rect 4953 3780 4957 3836
rect 4957 3780 5013 3836
rect 5013 3780 5017 3836
rect 4953 3776 5017 3780
rect 5033 3836 5097 3840
rect 5033 3780 5037 3836
rect 5037 3780 5093 3836
rect 5093 3780 5097 3836
rect 5033 3776 5097 3780
rect 12475 3836 12539 3840
rect 12475 3780 12479 3836
rect 12479 3780 12535 3836
rect 12535 3780 12539 3836
rect 12475 3776 12539 3780
rect 12555 3836 12619 3840
rect 12555 3780 12559 3836
rect 12559 3780 12615 3836
rect 12615 3780 12619 3836
rect 12555 3776 12619 3780
rect 12635 3836 12699 3840
rect 12635 3780 12639 3836
rect 12639 3780 12695 3836
rect 12695 3780 12699 3836
rect 12635 3776 12699 3780
rect 12715 3836 12779 3840
rect 12715 3780 12719 3836
rect 12719 3780 12775 3836
rect 12775 3780 12779 3836
rect 12715 3776 12779 3780
rect 20157 3836 20221 3840
rect 20157 3780 20161 3836
rect 20161 3780 20217 3836
rect 20217 3780 20221 3836
rect 20157 3776 20221 3780
rect 20237 3836 20301 3840
rect 20237 3780 20241 3836
rect 20241 3780 20297 3836
rect 20297 3780 20301 3836
rect 20237 3776 20301 3780
rect 20317 3836 20381 3840
rect 20317 3780 20321 3836
rect 20321 3780 20377 3836
rect 20377 3780 20381 3836
rect 20317 3776 20381 3780
rect 20397 3836 20461 3840
rect 20397 3780 20401 3836
rect 20401 3780 20457 3836
rect 20457 3780 20461 3836
rect 20397 3776 20461 3780
rect 27839 3836 27903 3840
rect 27839 3780 27843 3836
rect 27843 3780 27899 3836
rect 27899 3780 27903 3836
rect 27839 3776 27903 3780
rect 27919 3836 27983 3840
rect 27919 3780 27923 3836
rect 27923 3780 27979 3836
rect 27979 3780 27983 3836
rect 27919 3776 27983 3780
rect 27999 3836 28063 3840
rect 27999 3780 28003 3836
rect 28003 3780 28059 3836
rect 28059 3780 28063 3836
rect 27999 3776 28063 3780
rect 28079 3836 28143 3840
rect 28079 3780 28083 3836
rect 28083 3780 28139 3836
rect 28139 3780 28143 3836
rect 28079 3776 28143 3780
rect 8634 3292 8698 3296
rect 8634 3236 8638 3292
rect 8638 3236 8694 3292
rect 8694 3236 8698 3292
rect 8634 3232 8698 3236
rect 8714 3292 8778 3296
rect 8714 3236 8718 3292
rect 8718 3236 8774 3292
rect 8774 3236 8778 3292
rect 8714 3232 8778 3236
rect 8794 3292 8858 3296
rect 8794 3236 8798 3292
rect 8798 3236 8854 3292
rect 8854 3236 8858 3292
rect 8794 3232 8858 3236
rect 8874 3292 8938 3296
rect 8874 3236 8878 3292
rect 8878 3236 8934 3292
rect 8934 3236 8938 3292
rect 8874 3232 8938 3236
rect 16316 3292 16380 3296
rect 16316 3236 16320 3292
rect 16320 3236 16376 3292
rect 16376 3236 16380 3292
rect 16316 3232 16380 3236
rect 16396 3292 16460 3296
rect 16396 3236 16400 3292
rect 16400 3236 16456 3292
rect 16456 3236 16460 3292
rect 16396 3232 16460 3236
rect 16476 3292 16540 3296
rect 16476 3236 16480 3292
rect 16480 3236 16536 3292
rect 16536 3236 16540 3292
rect 16476 3232 16540 3236
rect 16556 3292 16620 3296
rect 16556 3236 16560 3292
rect 16560 3236 16616 3292
rect 16616 3236 16620 3292
rect 16556 3232 16620 3236
rect 23998 3292 24062 3296
rect 23998 3236 24002 3292
rect 24002 3236 24058 3292
rect 24058 3236 24062 3292
rect 23998 3232 24062 3236
rect 24078 3292 24142 3296
rect 24078 3236 24082 3292
rect 24082 3236 24138 3292
rect 24138 3236 24142 3292
rect 24078 3232 24142 3236
rect 24158 3292 24222 3296
rect 24158 3236 24162 3292
rect 24162 3236 24218 3292
rect 24218 3236 24222 3292
rect 24158 3232 24222 3236
rect 24238 3292 24302 3296
rect 24238 3236 24242 3292
rect 24242 3236 24298 3292
rect 24298 3236 24302 3292
rect 24238 3232 24302 3236
rect 31680 3292 31744 3296
rect 31680 3236 31684 3292
rect 31684 3236 31740 3292
rect 31740 3236 31744 3292
rect 31680 3232 31744 3236
rect 31760 3292 31824 3296
rect 31760 3236 31764 3292
rect 31764 3236 31820 3292
rect 31820 3236 31824 3292
rect 31760 3232 31824 3236
rect 31840 3292 31904 3296
rect 31840 3236 31844 3292
rect 31844 3236 31900 3292
rect 31900 3236 31904 3292
rect 31840 3232 31904 3236
rect 31920 3292 31984 3296
rect 31920 3236 31924 3292
rect 31924 3236 31980 3292
rect 31980 3236 31984 3292
rect 31920 3232 31984 3236
rect 4793 2748 4857 2752
rect 4793 2692 4797 2748
rect 4797 2692 4853 2748
rect 4853 2692 4857 2748
rect 4793 2688 4857 2692
rect 4873 2748 4937 2752
rect 4873 2692 4877 2748
rect 4877 2692 4933 2748
rect 4933 2692 4937 2748
rect 4873 2688 4937 2692
rect 4953 2748 5017 2752
rect 4953 2692 4957 2748
rect 4957 2692 5013 2748
rect 5013 2692 5017 2748
rect 4953 2688 5017 2692
rect 5033 2748 5097 2752
rect 5033 2692 5037 2748
rect 5037 2692 5093 2748
rect 5093 2692 5097 2748
rect 5033 2688 5097 2692
rect 12475 2748 12539 2752
rect 12475 2692 12479 2748
rect 12479 2692 12535 2748
rect 12535 2692 12539 2748
rect 12475 2688 12539 2692
rect 12555 2748 12619 2752
rect 12555 2692 12559 2748
rect 12559 2692 12615 2748
rect 12615 2692 12619 2748
rect 12555 2688 12619 2692
rect 12635 2748 12699 2752
rect 12635 2692 12639 2748
rect 12639 2692 12695 2748
rect 12695 2692 12699 2748
rect 12635 2688 12699 2692
rect 12715 2748 12779 2752
rect 12715 2692 12719 2748
rect 12719 2692 12775 2748
rect 12775 2692 12779 2748
rect 12715 2688 12779 2692
rect 20157 2748 20221 2752
rect 20157 2692 20161 2748
rect 20161 2692 20217 2748
rect 20217 2692 20221 2748
rect 20157 2688 20221 2692
rect 20237 2748 20301 2752
rect 20237 2692 20241 2748
rect 20241 2692 20297 2748
rect 20297 2692 20301 2748
rect 20237 2688 20301 2692
rect 20317 2748 20381 2752
rect 20317 2692 20321 2748
rect 20321 2692 20377 2748
rect 20377 2692 20381 2748
rect 20317 2688 20381 2692
rect 20397 2748 20461 2752
rect 20397 2692 20401 2748
rect 20401 2692 20457 2748
rect 20457 2692 20461 2748
rect 20397 2688 20461 2692
rect 27839 2748 27903 2752
rect 27839 2692 27843 2748
rect 27843 2692 27899 2748
rect 27899 2692 27903 2748
rect 27839 2688 27903 2692
rect 27919 2748 27983 2752
rect 27919 2692 27923 2748
rect 27923 2692 27979 2748
rect 27979 2692 27983 2748
rect 27919 2688 27983 2692
rect 27999 2748 28063 2752
rect 27999 2692 28003 2748
rect 28003 2692 28059 2748
rect 28059 2692 28063 2748
rect 27999 2688 28063 2692
rect 28079 2748 28143 2752
rect 28079 2692 28083 2748
rect 28083 2692 28139 2748
rect 28139 2692 28143 2748
rect 28079 2688 28143 2692
rect 8634 2204 8698 2208
rect 8634 2148 8638 2204
rect 8638 2148 8694 2204
rect 8694 2148 8698 2204
rect 8634 2144 8698 2148
rect 8714 2204 8778 2208
rect 8714 2148 8718 2204
rect 8718 2148 8774 2204
rect 8774 2148 8778 2204
rect 8714 2144 8778 2148
rect 8794 2204 8858 2208
rect 8794 2148 8798 2204
rect 8798 2148 8854 2204
rect 8854 2148 8858 2204
rect 8794 2144 8858 2148
rect 8874 2204 8938 2208
rect 8874 2148 8878 2204
rect 8878 2148 8934 2204
rect 8934 2148 8938 2204
rect 8874 2144 8938 2148
rect 16316 2204 16380 2208
rect 16316 2148 16320 2204
rect 16320 2148 16376 2204
rect 16376 2148 16380 2204
rect 16316 2144 16380 2148
rect 16396 2204 16460 2208
rect 16396 2148 16400 2204
rect 16400 2148 16456 2204
rect 16456 2148 16460 2204
rect 16396 2144 16460 2148
rect 16476 2204 16540 2208
rect 16476 2148 16480 2204
rect 16480 2148 16536 2204
rect 16536 2148 16540 2204
rect 16476 2144 16540 2148
rect 16556 2204 16620 2208
rect 16556 2148 16560 2204
rect 16560 2148 16616 2204
rect 16616 2148 16620 2204
rect 16556 2144 16620 2148
rect 23998 2204 24062 2208
rect 23998 2148 24002 2204
rect 24002 2148 24058 2204
rect 24058 2148 24062 2204
rect 23998 2144 24062 2148
rect 24078 2204 24142 2208
rect 24078 2148 24082 2204
rect 24082 2148 24138 2204
rect 24138 2148 24142 2204
rect 24078 2144 24142 2148
rect 24158 2204 24222 2208
rect 24158 2148 24162 2204
rect 24162 2148 24218 2204
rect 24218 2148 24222 2204
rect 24158 2144 24222 2148
rect 24238 2204 24302 2208
rect 24238 2148 24242 2204
rect 24242 2148 24298 2204
rect 24298 2148 24302 2204
rect 24238 2144 24302 2148
rect 31680 2204 31744 2208
rect 31680 2148 31684 2204
rect 31684 2148 31740 2204
rect 31740 2148 31744 2204
rect 31680 2144 31744 2148
rect 31760 2204 31824 2208
rect 31760 2148 31764 2204
rect 31764 2148 31820 2204
rect 31820 2148 31824 2204
rect 31760 2144 31824 2148
rect 31840 2204 31904 2208
rect 31840 2148 31844 2204
rect 31844 2148 31900 2204
rect 31900 2148 31904 2204
rect 31840 2144 31904 2148
rect 31920 2204 31984 2208
rect 31920 2148 31924 2204
rect 31924 2148 31980 2204
rect 31980 2148 31984 2204
rect 31920 2144 31984 2148
<< metal4 >>
rect 22139 34916 22205 34917
rect 22139 34852 22140 34916
rect 22204 34852 22205 34916
rect 22139 34851 22205 34852
rect 20851 34780 20917 34781
rect 20851 34716 20852 34780
rect 20916 34716 20917 34780
rect 20851 34715 20917 34716
rect 10179 34644 10245 34645
rect 10179 34580 10180 34644
rect 10244 34580 10245 34644
rect 10179 34579 10245 34580
rect 9259 34100 9325 34101
rect 9259 34036 9260 34100
rect 9324 34036 9325 34100
rect 9259 34035 9325 34036
rect 6315 33148 6381 33149
rect 6315 33084 6316 33148
rect 6380 33084 6381 33148
rect 6315 33083 6381 33084
rect 4785 32128 5105 32688
rect 4785 32064 4793 32128
rect 4857 32064 4873 32128
rect 4937 32064 4953 32128
rect 5017 32064 5033 32128
rect 5097 32064 5105 32128
rect 4785 31040 5105 32064
rect 4785 30976 4793 31040
rect 4857 30976 4873 31040
rect 4937 30976 4953 31040
rect 5017 30976 5033 31040
rect 5097 30976 5105 31040
rect 4785 29952 5105 30976
rect 4785 29888 4793 29952
rect 4857 29888 4873 29952
rect 4937 29888 4953 29952
rect 5017 29888 5033 29952
rect 5097 29888 5105 29952
rect 4785 28864 5105 29888
rect 4785 28800 4793 28864
rect 4857 28800 4873 28864
rect 4937 28800 4953 28864
rect 5017 28800 5033 28864
rect 5097 28800 5105 28864
rect 4785 27776 5105 28800
rect 4785 27712 4793 27776
rect 4857 27712 4873 27776
rect 4937 27712 4953 27776
rect 5017 27712 5033 27776
rect 5097 27712 5105 27776
rect 4785 26688 5105 27712
rect 4785 26624 4793 26688
rect 4857 26624 4873 26688
rect 4937 26624 4953 26688
rect 5017 26624 5033 26688
rect 5097 26624 5105 26688
rect 4785 25600 5105 26624
rect 4785 25536 4793 25600
rect 4857 25536 4873 25600
rect 4937 25536 4953 25600
rect 5017 25536 5033 25600
rect 5097 25536 5105 25600
rect 4785 24512 5105 25536
rect 5395 25532 5461 25533
rect 5395 25468 5396 25532
rect 5460 25468 5461 25532
rect 5395 25467 5461 25468
rect 4785 24448 4793 24512
rect 4857 24448 4873 24512
rect 4937 24448 4953 24512
rect 5017 24448 5033 24512
rect 5097 24448 5105 24512
rect 4785 23424 5105 24448
rect 4785 23360 4793 23424
rect 4857 23360 4873 23424
rect 4937 23360 4953 23424
rect 5017 23360 5033 23424
rect 5097 23360 5105 23424
rect 4785 22336 5105 23360
rect 4785 22272 4793 22336
rect 4857 22272 4873 22336
rect 4937 22272 4953 22336
rect 5017 22272 5033 22336
rect 5097 22272 5105 22336
rect 4785 21248 5105 22272
rect 4785 21184 4793 21248
rect 4857 21184 4873 21248
rect 4937 21184 4953 21248
rect 5017 21184 5033 21248
rect 5097 21184 5105 21248
rect 4785 20160 5105 21184
rect 4785 20096 4793 20160
rect 4857 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5105 20160
rect 4785 19072 5105 20096
rect 4785 19008 4793 19072
rect 4857 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5105 19072
rect 4785 17984 5105 19008
rect 4785 17920 4793 17984
rect 4857 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5105 17984
rect 4785 16896 5105 17920
rect 4785 16832 4793 16896
rect 4857 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5105 16896
rect 4785 15808 5105 16832
rect 4785 15744 4793 15808
rect 4857 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5105 15808
rect 4785 14720 5105 15744
rect 4785 14656 4793 14720
rect 4857 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5105 14720
rect 4785 13632 5105 14656
rect 4785 13568 4793 13632
rect 4857 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5105 13632
rect 4785 12544 5105 13568
rect 4785 12480 4793 12544
rect 4857 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5105 12544
rect 4785 11456 5105 12480
rect 4785 11392 4793 11456
rect 4857 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5105 11456
rect 4785 10368 5105 11392
rect 4785 10304 4793 10368
rect 4857 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5105 10368
rect 4785 9280 5105 10304
rect 5398 9621 5458 25467
rect 6318 23493 6378 33083
rect 8626 32672 8946 32688
rect 8626 32608 8634 32672
rect 8698 32608 8714 32672
rect 8778 32608 8794 32672
rect 8858 32608 8874 32672
rect 8938 32608 8946 32672
rect 8155 31924 8221 31925
rect 8155 31860 8156 31924
rect 8220 31860 8221 31924
rect 8155 31859 8221 31860
rect 6683 30836 6749 30837
rect 6683 30772 6684 30836
rect 6748 30772 6749 30836
rect 6683 30771 6749 30772
rect 6315 23492 6381 23493
rect 6315 23428 6316 23492
rect 6380 23428 6381 23492
rect 6315 23427 6381 23428
rect 6686 12450 6746 30771
rect 6867 30700 6933 30701
rect 6867 30636 6868 30700
rect 6932 30636 6933 30700
rect 6867 30635 6933 30636
rect 6870 24717 6930 30635
rect 7051 30156 7117 30157
rect 7051 30092 7052 30156
rect 7116 30092 7117 30156
rect 7051 30091 7117 30092
rect 6867 24716 6933 24717
rect 6867 24652 6868 24716
rect 6932 24652 6933 24716
rect 6867 24651 6933 24652
rect 7054 24309 7114 30091
rect 7051 24308 7117 24309
rect 7051 24244 7052 24308
rect 7116 24244 7117 24308
rect 7051 24243 7117 24244
rect 8158 22813 8218 31859
rect 8626 31584 8946 32608
rect 8626 31520 8634 31584
rect 8698 31520 8714 31584
rect 8778 31520 8794 31584
rect 8858 31520 8874 31584
rect 8938 31520 8946 31584
rect 8626 30496 8946 31520
rect 8626 30432 8634 30496
rect 8698 30432 8714 30496
rect 8778 30432 8794 30496
rect 8858 30432 8874 30496
rect 8938 30432 8946 30496
rect 8626 29408 8946 30432
rect 8626 29344 8634 29408
rect 8698 29344 8714 29408
rect 8778 29344 8794 29408
rect 8858 29344 8874 29408
rect 8938 29344 8946 29408
rect 8626 28320 8946 29344
rect 8626 28256 8634 28320
rect 8698 28256 8714 28320
rect 8778 28256 8794 28320
rect 8858 28256 8874 28320
rect 8938 28256 8946 28320
rect 8626 27232 8946 28256
rect 8626 27168 8634 27232
rect 8698 27168 8714 27232
rect 8778 27168 8794 27232
rect 8858 27168 8874 27232
rect 8938 27168 8946 27232
rect 8626 26144 8946 27168
rect 8626 26080 8634 26144
rect 8698 26080 8714 26144
rect 8778 26080 8794 26144
rect 8858 26080 8874 26144
rect 8938 26080 8946 26144
rect 8626 25056 8946 26080
rect 8626 24992 8634 25056
rect 8698 24992 8714 25056
rect 8778 24992 8794 25056
rect 8858 24992 8874 25056
rect 8938 24992 8946 25056
rect 8626 23968 8946 24992
rect 8626 23904 8634 23968
rect 8698 23904 8714 23968
rect 8778 23904 8794 23968
rect 8858 23904 8874 23968
rect 8938 23904 8946 23968
rect 8626 22880 8946 23904
rect 9262 23357 9322 34035
rect 9443 29068 9509 29069
rect 9443 29004 9444 29068
rect 9508 29004 9509 29068
rect 9443 29003 9509 29004
rect 9259 23356 9325 23357
rect 9259 23292 9260 23356
rect 9324 23292 9325 23356
rect 9259 23291 9325 23292
rect 8626 22816 8634 22880
rect 8698 22816 8714 22880
rect 8778 22816 8794 22880
rect 8858 22816 8874 22880
rect 8938 22816 8946 22880
rect 8155 22812 8221 22813
rect 8155 22748 8156 22812
rect 8220 22748 8221 22812
rect 8155 22747 8221 22748
rect 6867 21860 6933 21861
rect 6867 21796 6868 21860
rect 6932 21796 6933 21860
rect 6867 21795 6933 21796
rect 6870 13429 6930 21795
rect 8626 21792 8946 22816
rect 8626 21728 8634 21792
rect 8698 21728 8714 21792
rect 8778 21728 8794 21792
rect 8858 21728 8874 21792
rect 8938 21728 8946 21792
rect 8626 20704 8946 21728
rect 8626 20640 8634 20704
rect 8698 20640 8714 20704
rect 8778 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8946 20704
rect 8626 19616 8946 20640
rect 8626 19552 8634 19616
rect 8698 19552 8714 19616
rect 8778 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8946 19616
rect 8626 18528 8946 19552
rect 8626 18464 8634 18528
rect 8698 18464 8714 18528
rect 8778 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8946 18528
rect 8626 17440 8946 18464
rect 8626 17376 8634 17440
rect 8698 17376 8714 17440
rect 8778 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8946 17440
rect 8626 16352 8946 17376
rect 8626 16288 8634 16352
rect 8698 16288 8714 16352
rect 8778 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8946 16352
rect 8626 15264 8946 16288
rect 8626 15200 8634 15264
rect 8698 15200 8714 15264
rect 8778 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8946 15264
rect 8626 14176 8946 15200
rect 8626 14112 8634 14176
rect 8698 14112 8714 14176
rect 8778 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8946 14176
rect 6867 13428 6933 13429
rect 6867 13364 6868 13428
rect 6932 13364 6933 13428
rect 6867 13363 6933 13364
rect 6502 12390 6746 12450
rect 8626 13088 8946 14112
rect 8626 13024 8634 13088
rect 8698 13024 8714 13088
rect 8778 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8946 13088
rect 6502 10165 6562 12390
rect 8626 12000 8946 13024
rect 8626 11936 8634 12000
rect 8698 11936 8714 12000
rect 8778 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8946 12000
rect 8626 10912 8946 11936
rect 8626 10848 8634 10912
rect 8698 10848 8714 10912
rect 8778 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8946 10912
rect 6499 10164 6565 10165
rect 6499 10100 6500 10164
rect 6564 10100 6565 10164
rect 6499 10099 6565 10100
rect 8626 9824 8946 10848
rect 8626 9760 8634 9824
rect 8698 9760 8714 9824
rect 8778 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8946 9824
rect 5395 9620 5461 9621
rect 5395 9556 5396 9620
rect 5460 9556 5461 9620
rect 5395 9555 5461 9556
rect 4785 9216 4793 9280
rect 4857 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5105 9280
rect 4785 8192 5105 9216
rect 4785 8128 4793 8192
rect 4857 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5105 8192
rect 4785 7104 5105 8128
rect 4785 7040 4793 7104
rect 4857 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5105 7104
rect 4785 6016 5105 7040
rect 4785 5952 4793 6016
rect 4857 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5105 6016
rect 4785 4928 5105 5952
rect 4785 4864 4793 4928
rect 4857 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5105 4928
rect 4785 3840 5105 4864
rect 4785 3776 4793 3840
rect 4857 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5105 3840
rect 4785 2752 5105 3776
rect 4785 2688 4793 2752
rect 4857 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5105 2752
rect 4785 2128 5105 2688
rect 8626 8736 8946 9760
rect 8626 8672 8634 8736
rect 8698 8672 8714 8736
rect 8778 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8946 8736
rect 8626 7648 8946 8672
rect 9446 7853 9506 29003
rect 10182 21997 10242 34579
rect 12203 33828 12269 33829
rect 12203 33764 12204 33828
rect 12268 33764 12269 33828
rect 12203 33763 12269 33764
rect 10731 31244 10797 31245
rect 10731 31180 10732 31244
rect 10796 31180 10797 31244
rect 10731 31179 10797 31180
rect 10179 21996 10245 21997
rect 10179 21932 10180 21996
rect 10244 21932 10245 21996
rect 10179 21931 10245 21932
rect 10547 16964 10613 16965
rect 10547 16900 10548 16964
rect 10612 16900 10613 16964
rect 10547 16899 10613 16900
rect 10550 10573 10610 16899
rect 10734 16557 10794 31179
rect 11467 30700 11533 30701
rect 11467 30636 11468 30700
rect 11532 30636 11533 30700
rect 11467 30635 11533 30636
rect 11470 22677 11530 30635
rect 11835 30428 11901 30429
rect 11835 30364 11836 30428
rect 11900 30364 11901 30428
rect 11835 30363 11901 30364
rect 11467 22676 11533 22677
rect 11467 22612 11468 22676
rect 11532 22612 11533 22676
rect 11467 22611 11533 22612
rect 10915 20772 10981 20773
rect 10915 20708 10916 20772
rect 10980 20708 10981 20772
rect 10915 20707 10981 20708
rect 11651 20772 11717 20773
rect 11651 20708 11652 20772
rect 11716 20708 11717 20772
rect 11651 20707 11717 20708
rect 10918 17237 10978 20707
rect 10915 17236 10981 17237
rect 10915 17172 10916 17236
rect 10980 17172 10981 17236
rect 10915 17171 10981 17172
rect 10731 16556 10797 16557
rect 10731 16492 10732 16556
rect 10796 16492 10797 16556
rect 10731 16491 10797 16492
rect 11654 15333 11714 20707
rect 11651 15332 11717 15333
rect 11651 15268 11652 15332
rect 11716 15268 11717 15332
rect 11651 15267 11717 15268
rect 10547 10572 10613 10573
rect 10547 10508 10548 10572
rect 10612 10508 10613 10572
rect 10547 10507 10613 10508
rect 9443 7852 9509 7853
rect 9443 7788 9444 7852
rect 9508 7788 9509 7852
rect 9443 7787 9509 7788
rect 8626 7584 8634 7648
rect 8698 7584 8714 7648
rect 8778 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8946 7648
rect 8626 6560 8946 7584
rect 11838 7309 11898 30363
rect 12019 27572 12085 27573
rect 12019 27508 12020 27572
rect 12084 27508 12085 27572
rect 12019 27507 12085 27508
rect 12022 25533 12082 27507
rect 12019 25532 12085 25533
rect 12019 25468 12020 25532
rect 12084 25468 12085 25532
rect 12019 25467 12085 25468
rect 12022 22269 12082 25467
rect 12019 22268 12085 22269
rect 12019 22204 12020 22268
rect 12084 22204 12085 22268
rect 12019 22203 12085 22204
rect 12206 21725 12266 33763
rect 15147 33420 15213 33421
rect 15147 33356 15148 33420
rect 15212 33356 15213 33420
rect 15147 33355 15213 33356
rect 12467 32128 12787 32688
rect 12467 32064 12475 32128
rect 12539 32064 12555 32128
rect 12619 32064 12635 32128
rect 12699 32064 12715 32128
rect 12779 32064 12787 32128
rect 12467 31040 12787 32064
rect 12467 30976 12475 31040
rect 12539 30976 12555 31040
rect 12619 30976 12635 31040
rect 12699 30976 12715 31040
rect 12779 30976 12787 31040
rect 12467 29952 12787 30976
rect 14227 30972 14293 30973
rect 14227 30908 14228 30972
rect 14292 30908 14293 30972
rect 14227 30907 14293 30908
rect 12467 29888 12475 29952
rect 12539 29888 12555 29952
rect 12619 29888 12635 29952
rect 12699 29888 12715 29952
rect 12779 29888 12787 29952
rect 12467 28864 12787 29888
rect 12939 29748 13005 29749
rect 12939 29684 12940 29748
rect 13004 29684 13005 29748
rect 12939 29683 13005 29684
rect 12467 28800 12475 28864
rect 12539 28800 12555 28864
rect 12619 28800 12635 28864
rect 12699 28800 12715 28864
rect 12779 28800 12787 28864
rect 12467 27776 12787 28800
rect 12467 27712 12475 27776
rect 12539 27712 12555 27776
rect 12619 27712 12635 27776
rect 12699 27712 12715 27776
rect 12779 27712 12787 27776
rect 12467 26688 12787 27712
rect 12467 26624 12475 26688
rect 12539 26624 12555 26688
rect 12619 26624 12635 26688
rect 12699 26624 12715 26688
rect 12779 26624 12787 26688
rect 12467 25600 12787 26624
rect 12467 25536 12475 25600
rect 12539 25536 12555 25600
rect 12619 25536 12635 25600
rect 12699 25536 12715 25600
rect 12779 25536 12787 25600
rect 12467 24512 12787 25536
rect 12467 24448 12475 24512
rect 12539 24448 12555 24512
rect 12619 24448 12635 24512
rect 12699 24448 12715 24512
rect 12779 24448 12787 24512
rect 12467 23424 12787 24448
rect 12467 23360 12475 23424
rect 12539 23360 12555 23424
rect 12619 23360 12635 23424
rect 12699 23360 12715 23424
rect 12779 23360 12787 23424
rect 12467 22336 12787 23360
rect 12467 22272 12475 22336
rect 12539 22272 12555 22336
rect 12619 22272 12635 22336
rect 12699 22272 12715 22336
rect 12779 22272 12787 22336
rect 12203 21724 12269 21725
rect 12203 21660 12204 21724
rect 12268 21660 12269 21724
rect 12203 21659 12269 21660
rect 12467 21248 12787 22272
rect 12942 21453 13002 29683
rect 13491 29340 13557 29341
rect 13491 29276 13492 29340
rect 13556 29276 13557 29340
rect 13491 29275 13557 29276
rect 13307 27980 13373 27981
rect 13307 27916 13308 27980
rect 13372 27916 13373 27980
rect 13307 27915 13373 27916
rect 13310 23357 13370 27915
rect 13494 26077 13554 29275
rect 13675 27844 13741 27845
rect 13675 27780 13676 27844
rect 13740 27780 13741 27844
rect 13675 27779 13741 27780
rect 13678 26213 13738 27779
rect 14230 26757 14290 30907
rect 14411 30428 14477 30429
rect 14411 30364 14412 30428
rect 14476 30364 14477 30428
rect 14411 30363 14477 30364
rect 14227 26756 14293 26757
rect 14227 26692 14228 26756
rect 14292 26692 14293 26756
rect 14227 26691 14293 26692
rect 13675 26212 13741 26213
rect 13675 26148 13676 26212
rect 13740 26148 13741 26212
rect 13675 26147 13741 26148
rect 13491 26076 13557 26077
rect 13491 26012 13492 26076
rect 13556 26012 13557 26076
rect 13491 26011 13557 26012
rect 13494 23493 13554 26011
rect 13491 23492 13557 23493
rect 13491 23428 13492 23492
rect 13556 23428 13557 23492
rect 13491 23427 13557 23428
rect 13307 23356 13373 23357
rect 13307 23292 13308 23356
rect 13372 23292 13373 23356
rect 13307 23291 13373 23292
rect 13491 22948 13557 22949
rect 13491 22884 13492 22948
rect 13556 22884 13557 22948
rect 13491 22883 13557 22884
rect 13307 22404 13373 22405
rect 13307 22340 13308 22404
rect 13372 22340 13373 22404
rect 13307 22339 13373 22340
rect 13123 21860 13189 21861
rect 13123 21796 13124 21860
rect 13188 21796 13189 21860
rect 13123 21795 13189 21796
rect 12939 21452 13005 21453
rect 12939 21388 12940 21452
rect 13004 21388 13005 21452
rect 12939 21387 13005 21388
rect 12467 21184 12475 21248
rect 12539 21184 12555 21248
rect 12619 21184 12635 21248
rect 12699 21184 12715 21248
rect 12779 21184 12787 21248
rect 12019 21180 12085 21181
rect 12019 21116 12020 21180
rect 12084 21116 12085 21180
rect 12019 21115 12085 21116
rect 12022 14109 12082 21115
rect 12203 20772 12269 20773
rect 12203 20708 12204 20772
rect 12268 20708 12269 20772
rect 12203 20707 12269 20708
rect 12206 16557 12266 20707
rect 12467 20160 12787 21184
rect 12467 20096 12475 20160
rect 12539 20096 12555 20160
rect 12619 20096 12635 20160
rect 12699 20096 12715 20160
rect 12779 20096 12787 20160
rect 12467 19072 12787 20096
rect 12939 20092 13005 20093
rect 12939 20028 12940 20092
rect 13004 20028 13005 20092
rect 12939 20027 13005 20028
rect 12467 19008 12475 19072
rect 12539 19008 12555 19072
rect 12619 19008 12635 19072
rect 12699 19008 12715 19072
rect 12779 19008 12787 19072
rect 12467 17984 12787 19008
rect 12942 18869 13002 20027
rect 12939 18868 13005 18869
rect 12939 18804 12940 18868
rect 13004 18804 13005 18868
rect 12939 18803 13005 18804
rect 12467 17920 12475 17984
rect 12539 17920 12555 17984
rect 12619 17920 12635 17984
rect 12699 17920 12715 17984
rect 12779 17920 12787 17984
rect 12467 16896 12787 17920
rect 12467 16832 12475 16896
rect 12539 16832 12555 16896
rect 12619 16832 12635 16896
rect 12699 16832 12715 16896
rect 12779 16832 12787 16896
rect 12203 16556 12269 16557
rect 12203 16492 12204 16556
rect 12268 16492 12269 16556
rect 12203 16491 12269 16492
rect 12467 15808 12787 16832
rect 12467 15744 12475 15808
rect 12539 15744 12555 15808
rect 12619 15744 12635 15808
rect 12699 15744 12715 15808
rect 12779 15744 12787 15808
rect 12467 14720 12787 15744
rect 12467 14656 12475 14720
rect 12539 14656 12555 14720
rect 12619 14656 12635 14720
rect 12699 14656 12715 14720
rect 12779 14656 12787 14720
rect 12019 14108 12085 14109
rect 12019 14044 12020 14108
rect 12084 14044 12085 14108
rect 12019 14043 12085 14044
rect 12467 13632 12787 14656
rect 12467 13568 12475 13632
rect 12539 13568 12555 13632
rect 12619 13568 12635 13632
rect 12699 13568 12715 13632
rect 12779 13568 12787 13632
rect 12467 12544 12787 13568
rect 12467 12480 12475 12544
rect 12539 12480 12555 12544
rect 12619 12480 12635 12544
rect 12699 12480 12715 12544
rect 12779 12480 12787 12544
rect 12467 11456 12787 12480
rect 12467 11392 12475 11456
rect 12539 11392 12555 11456
rect 12619 11392 12635 11456
rect 12699 11392 12715 11456
rect 12779 11392 12787 11456
rect 12467 10368 12787 11392
rect 12467 10304 12475 10368
rect 12539 10304 12555 10368
rect 12619 10304 12635 10368
rect 12699 10304 12715 10368
rect 12779 10304 12787 10368
rect 12467 9280 12787 10304
rect 12467 9216 12475 9280
rect 12539 9216 12555 9280
rect 12619 9216 12635 9280
rect 12699 9216 12715 9280
rect 12779 9216 12787 9280
rect 12467 8192 12787 9216
rect 13126 8533 13186 21795
rect 13310 21317 13370 22339
rect 13307 21316 13373 21317
rect 13307 21252 13308 21316
rect 13372 21252 13373 21316
rect 13307 21251 13373 21252
rect 13307 19412 13373 19413
rect 13307 19348 13308 19412
rect 13372 19348 13373 19412
rect 13307 19347 13373 19348
rect 13310 9077 13370 19347
rect 13307 9076 13373 9077
rect 13307 9012 13308 9076
rect 13372 9012 13373 9076
rect 13307 9011 13373 9012
rect 13123 8532 13189 8533
rect 13123 8468 13124 8532
rect 13188 8468 13189 8532
rect 13123 8467 13189 8468
rect 12467 8128 12475 8192
rect 12539 8128 12555 8192
rect 12619 8128 12635 8192
rect 12699 8128 12715 8192
rect 12779 8128 12787 8192
rect 11835 7308 11901 7309
rect 11835 7244 11836 7308
rect 11900 7244 11901 7308
rect 11835 7243 11901 7244
rect 8626 6496 8634 6560
rect 8698 6496 8714 6560
rect 8778 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8946 6560
rect 8626 5472 8946 6496
rect 8626 5408 8634 5472
rect 8698 5408 8714 5472
rect 8778 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8946 5472
rect 8626 4384 8946 5408
rect 8626 4320 8634 4384
rect 8698 4320 8714 4384
rect 8778 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8946 4384
rect 8626 3296 8946 4320
rect 8626 3232 8634 3296
rect 8698 3232 8714 3296
rect 8778 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8946 3296
rect 8626 2208 8946 3232
rect 8626 2144 8634 2208
rect 8698 2144 8714 2208
rect 8778 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8946 2208
rect 8626 2128 8946 2144
rect 12467 7104 12787 8128
rect 12467 7040 12475 7104
rect 12539 7040 12555 7104
rect 12619 7040 12635 7104
rect 12699 7040 12715 7104
rect 12779 7040 12787 7104
rect 12467 6016 12787 7040
rect 12467 5952 12475 6016
rect 12539 5952 12555 6016
rect 12619 5952 12635 6016
rect 12699 5952 12715 6016
rect 12779 5952 12787 6016
rect 12467 4928 12787 5952
rect 13494 5133 13554 22883
rect 13678 19350 13738 26147
rect 14043 26076 14109 26077
rect 14043 26012 14044 26076
rect 14108 26012 14109 26076
rect 14043 26011 14109 26012
rect 13859 24580 13925 24581
rect 13859 24516 13860 24580
rect 13924 24516 13925 24580
rect 13859 24515 13925 24516
rect 13862 24306 13922 24515
rect 14046 24445 14106 26011
rect 14227 25532 14293 25533
rect 14227 25468 14228 25532
rect 14292 25468 14293 25532
rect 14227 25467 14293 25468
rect 14043 24444 14109 24445
rect 14043 24380 14044 24444
rect 14108 24380 14109 24444
rect 14043 24379 14109 24380
rect 13862 24246 14106 24306
rect 13859 24172 13925 24173
rect 13859 24108 13860 24172
rect 13924 24108 13925 24172
rect 13859 24107 13925 24108
rect 13862 22677 13922 24107
rect 13859 22676 13925 22677
rect 13859 22612 13860 22676
rect 13924 22612 13925 22676
rect 13859 22611 13925 22612
rect 13862 22269 13922 22611
rect 13859 22268 13925 22269
rect 13859 22204 13860 22268
rect 13924 22204 13925 22268
rect 13859 22203 13925 22204
rect 13678 19290 13922 19350
rect 13862 12450 13922 19290
rect 14046 17781 14106 24246
rect 14230 21725 14290 25467
rect 14227 21724 14293 21725
rect 14227 21660 14228 21724
rect 14292 21660 14293 21724
rect 14227 21659 14293 21660
rect 14043 17780 14109 17781
rect 14043 17716 14044 17780
rect 14108 17716 14109 17780
rect 14043 17715 14109 17716
rect 13862 12390 14106 12450
rect 14046 6901 14106 12390
rect 14414 7445 14474 30363
rect 15150 30157 15210 33355
rect 16067 33284 16133 33285
rect 16067 33220 16068 33284
rect 16132 33220 16133 33284
rect 16067 33219 16133 33220
rect 15515 30972 15581 30973
rect 15515 30908 15516 30972
rect 15580 30908 15581 30972
rect 15515 30907 15581 30908
rect 15147 30156 15213 30157
rect 15147 30092 15148 30156
rect 15212 30092 15213 30156
rect 15147 30091 15213 30092
rect 14779 28252 14845 28253
rect 14779 28188 14780 28252
rect 14844 28188 14845 28252
rect 14779 28187 14845 28188
rect 14595 28116 14661 28117
rect 14595 28052 14596 28116
rect 14660 28052 14661 28116
rect 14595 28051 14661 28052
rect 14598 25941 14658 28051
rect 14782 26485 14842 28187
rect 15147 26756 15213 26757
rect 15147 26692 15148 26756
rect 15212 26692 15213 26756
rect 15147 26691 15213 26692
rect 14779 26484 14845 26485
rect 14779 26420 14780 26484
rect 14844 26420 14845 26484
rect 14779 26419 14845 26420
rect 14595 25940 14661 25941
rect 14595 25876 14596 25940
rect 14660 25876 14661 25940
rect 14595 25875 14661 25876
rect 14595 25532 14661 25533
rect 14595 25468 14596 25532
rect 14660 25468 14661 25532
rect 14595 25467 14661 25468
rect 14598 25261 14658 25467
rect 14782 25261 14842 26419
rect 14963 26348 15029 26349
rect 14963 26284 14964 26348
rect 15028 26284 15029 26348
rect 14963 26283 15029 26284
rect 14595 25260 14661 25261
rect 14595 25196 14596 25260
rect 14660 25196 14661 25260
rect 14595 25195 14661 25196
rect 14779 25260 14845 25261
rect 14779 25196 14780 25260
rect 14844 25196 14845 25260
rect 14779 25195 14845 25196
rect 14779 24716 14845 24717
rect 14779 24652 14780 24716
rect 14844 24652 14845 24716
rect 14779 24651 14845 24652
rect 14595 23764 14661 23765
rect 14595 23700 14596 23764
rect 14660 23700 14661 23764
rect 14595 23699 14661 23700
rect 14598 20637 14658 23699
rect 14782 23357 14842 24651
rect 14779 23356 14845 23357
rect 14779 23292 14780 23356
rect 14844 23292 14845 23356
rect 14966 23354 15026 26283
rect 15150 24037 15210 26691
rect 15331 26484 15397 26485
rect 15331 26420 15332 26484
rect 15396 26420 15397 26484
rect 15331 26419 15397 26420
rect 15334 24581 15394 26419
rect 15518 24853 15578 30907
rect 15699 29068 15765 29069
rect 15699 29004 15700 29068
rect 15764 29004 15765 29068
rect 15699 29003 15765 29004
rect 15702 26349 15762 29003
rect 15883 28116 15949 28117
rect 15883 28052 15884 28116
rect 15948 28052 15949 28116
rect 15883 28051 15949 28052
rect 15699 26348 15765 26349
rect 15699 26284 15700 26348
rect 15764 26284 15765 26348
rect 15699 26283 15765 26284
rect 15515 24852 15581 24853
rect 15515 24788 15516 24852
rect 15580 24788 15581 24852
rect 15515 24787 15581 24788
rect 15515 24716 15581 24717
rect 15515 24652 15516 24716
rect 15580 24652 15581 24716
rect 15515 24651 15581 24652
rect 15331 24580 15397 24581
rect 15331 24516 15332 24580
rect 15396 24516 15397 24580
rect 15331 24515 15397 24516
rect 15331 24308 15397 24309
rect 15331 24244 15332 24308
rect 15396 24244 15397 24308
rect 15331 24243 15397 24244
rect 15147 24036 15213 24037
rect 15147 23972 15148 24036
rect 15212 23972 15213 24036
rect 15147 23971 15213 23972
rect 15147 23356 15213 23357
rect 15147 23354 15148 23356
rect 14966 23294 15148 23354
rect 14779 23291 14845 23292
rect 15147 23292 15148 23294
rect 15212 23292 15213 23356
rect 15147 23291 15213 23292
rect 14595 20636 14661 20637
rect 14595 20572 14596 20636
rect 14660 20572 14661 20636
rect 14595 20571 14661 20572
rect 15147 16284 15213 16285
rect 15147 16220 15148 16284
rect 15212 16220 15213 16284
rect 15147 16219 15213 16220
rect 15150 14245 15210 16219
rect 15147 14244 15213 14245
rect 15147 14180 15148 14244
rect 15212 14180 15213 14244
rect 15147 14179 15213 14180
rect 15334 8941 15394 24243
rect 15518 23629 15578 24651
rect 15515 23628 15581 23629
rect 15515 23564 15516 23628
rect 15580 23564 15581 23628
rect 15515 23563 15581 23564
rect 15515 19548 15581 19549
rect 15515 19484 15516 19548
rect 15580 19484 15581 19548
rect 15515 19483 15581 19484
rect 15518 14109 15578 19483
rect 15702 18869 15762 26283
rect 15886 24989 15946 28051
rect 16070 27573 16130 33219
rect 19931 32740 19997 32741
rect 16308 32672 16628 32688
rect 19931 32676 19932 32740
rect 19996 32676 19997 32740
rect 19931 32675 19997 32676
rect 16308 32608 16316 32672
rect 16380 32608 16396 32672
rect 16460 32608 16476 32672
rect 16540 32608 16556 32672
rect 16620 32608 16628 32672
rect 16308 31584 16628 32608
rect 16308 31520 16316 31584
rect 16380 31520 16396 31584
rect 16460 31520 16476 31584
rect 16540 31520 16556 31584
rect 16620 31520 16628 31584
rect 16308 30496 16628 31520
rect 17723 31380 17789 31381
rect 17723 31316 17724 31380
rect 17788 31316 17789 31380
rect 17723 31315 17789 31316
rect 16308 30432 16316 30496
rect 16380 30432 16396 30496
rect 16460 30432 16476 30496
rect 16540 30432 16556 30496
rect 16620 30432 16628 30496
rect 16308 29408 16628 30432
rect 17171 29884 17237 29885
rect 17171 29820 17172 29884
rect 17236 29820 17237 29884
rect 17171 29819 17237 29820
rect 16308 29344 16316 29408
rect 16380 29344 16396 29408
rect 16460 29344 16476 29408
rect 16540 29344 16556 29408
rect 16620 29344 16628 29408
rect 16308 28320 16628 29344
rect 16987 28524 17053 28525
rect 16987 28460 16988 28524
rect 17052 28460 17053 28524
rect 16987 28459 17053 28460
rect 16308 28256 16316 28320
rect 16380 28256 16396 28320
rect 16460 28256 16476 28320
rect 16540 28256 16556 28320
rect 16620 28256 16628 28320
rect 16067 27572 16133 27573
rect 16067 27508 16068 27572
rect 16132 27508 16133 27572
rect 16067 27507 16133 27508
rect 16308 27232 16628 28256
rect 16803 28252 16869 28253
rect 16803 28188 16804 28252
rect 16868 28188 16869 28252
rect 16803 28187 16869 28188
rect 16308 27168 16316 27232
rect 16380 27168 16396 27232
rect 16460 27168 16476 27232
rect 16540 27168 16556 27232
rect 16620 27168 16628 27232
rect 16067 27164 16133 27165
rect 16067 27100 16068 27164
rect 16132 27100 16133 27164
rect 16067 27099 16133 27100
rect 15883 24988 15949 24989
rect 15883 24924 15884 24988
rect 15948 24924 15949 24988
rect 15883 24923 15949 24924
rect 16070 24717 16130 27099
rect 16308 26144 16628 27168
rect 16806 26485 16866 28187
rect 16803 26484 16869 26485
rect 16803 26420 16804 26484
rect 16868 26420 16869 26484
rect 16803 26419 16869 26420
rect 16803 26348 16869 26349
rect 16803 26284 16804 26348
rect 16868 26284 16869 26348
rect 16803 26283 16869 26284
rect 16308 26080 16316 26144
rect 16380 26080 16396 26144
rect 16460 26080 16476 26144
rect 16540 26080 16556 26144
rect 16620 26080 16628 26144
rect 16308 25056 16628 26080
rect 16308 24992 16316 25056
rect 16380 24992 16396 25056
rect 16460 24992 16476 25056
rect 16540 24992 16556 25056
rect 16620 24992 16628 25056
rect 16067 24716 16133 24717
rect 16067 24652 16068 24716
rect 16132 24652 16133 24716
rect 16067 24651 16133 24652
rect 15883 21860 15949 21861
rect 15883 21796 15884 21860
rect 15948 21796 15949 21860
rect 15883 21795 15949 21796
rect 15886 19549 15946 21795
rect 15883 19548 15949 19549
rect 15883 19484 15884 19548
rect 15948 19484 15949 19548
rect 15883 19483 15949 19484
rect 16070 19350 16130 24651
rect 15886 19290 16130 19350
rect 16308 23968 16628 24992
rect 16806 24445 16866 26283
rect 16803 24444 16869 24445
rect 16803 24380 16804 24444
rect 16868 24380 16869 24444
rect 16803 24379 16869 24380
rect 16803 24036 16869 24037
rect 16803 23972 16804 24036
rect 16868 23972 16869 24036
rect 16803 23971 16869 23972
rect 16308 23904 16316 23968
rect 16380 23904 16396 23968
rect 16460 23904 16476 23968
rect 16540 23904 16556 23968
rect 16620 23904 16628 23968
rect 16308 22880 16628 23904
rect 16308 22816 16316 22880
rect 16380 22816 16396 22880
rect 16460 22816 16476 22880
rect 16540 22816 16556 22880
rect 16620 22816 16628 22880
rect 16308 21792 16628 22816
rect 16806 22269 16866 23971
rect 16990 23357 17050 28459
rect 17174 26893 17234 29819
rect 17539 29476 17605 29477
rect 17539 29412 17540 29476
rect 17604 29412 17605 29476
rect 17539 29411 17605 29412
rect 17355 27300 17421 27301
rect 17355 27236 17356 27300
rect 17420 27236 17421 27300
rect 17355 27235 17421 27236
rect 17171 26892 17237 26893
rect 17171 26828 17172 26892
rect 17236 26828 17237 26892
rect 17171 26827 17237 26828
rect 17171 26076 17237 26077
rect 17171 26012 17172 26076
rect 17236 26012 17237 26076
rect 17171 26011 17237 26012
rect 17174 23901 17234 26011
rect 17358 25533 17418 27235
rect 17542 25669 17602 29411
rect 17539 25668 17605 25669
rect 17539 25604 17540 25668
rect 17604 25604 17605 25668
rect 17539 25603 17605 25604
rect 17355 25532 17421 25533
rect 17355 25468 17356 25532
rect 17420 25468 17421 25532
rect 17355 25467 17421 25468
rect 17539 25124 17605 25125
rect 17539 25060 17540 25124
rect 17604 25060 17605 25124
rect 17539 25059 17605 25060
rect 17355 24716 17421 24717
rect 17355 24652 17356 24716
rect 17420 24652 17421 24716
rect 17355 24651 17421 24652
rect 17171 23900 17237 23901
rect 17171 23836 17172 23900
rect 17236 23836 17237 23900
rect 17171 23835 17237 23836
rect 16987 23356 17053 23357
rect 16987 23292 16988 23356
rect 17052 23292 17053 23356
rect 16987 23291 17053 23292
rect 17171 22812 17237 22813
rect 17171 22748 17172 22812
rect 17236 22748 17237 22812
rect 17171 22747 17237 22748
rect 16987 22676 17053 22677
rect 16987 22612 16988 22676
rect 17052 22612 17053 22676
rect 16987 22611 17053 22612
rect 16803 22268 16869 22269
rect 16803 22204 16804 22268
rect 16868 22204 16869 22268
rect 16803 22203 16869 22204
rect 16308 21728 16316 21792
rect 16380 21728 16396 21792
rect 16460 21728 16476 21792
rect 16540 21728 16556 21792
rect 16620 21728 16628 21792
rect 16308 20704 16628 21728
rect 16990 21450 17050 22611
rect 17174 21589 17234 22747
rect 17358 22674 17418 24651
rect 17542 24037 17602 25059
rect 17539 24036 17605 24037
rect 17539 23972 17540 24036
rect 17604 23972 17605 24036
rect 17539 23971 17605 23972
rect 17726 23901 17786 31315
rect 18091 31108 18157 31109
rect 18091 31044 18092 31108
rect 18156 31044 18157 31108
rect 18091 31043 18157 31044
rect 17907 30020 17973 30021
rect 17907 29956 17908 30020
rect 17972 29956 17973 30020
rect 17907 29955 17973 29956
rect 17910 26757 17970 29955
rect 17907 26756 17973 26757
rect 17907 26692 17908 26756
rect 17972 26692 17973 26756
rect 17907 26691 17973 26692
rect 18094 26485 18154 31043
rect 19747 30836 19813 30837
rect 19747 30772 19748 30836
rect 19812 30772 19813 30836
rect 19747 30771 19813 30772
rect 19195 30700 19261 30701
rect 19195 30636 19196 30700
rect 19260 30636 19261 30700
rect 19195 30635 19261 30636
rect 19011 30428 19077 30429
rect 19011 30390 19012 30428
rect 18830 30364 19012 30390
rect 19076 30364 19077 30428
rect 18830 30363 19077 30364
rect 18830 30330 19074 30363
rect 18275 29748 18341 29749
rect 18275 29684 18276 29748
rect 18340 29684 18341 29748
rect 18275 29683 18341 29684
rect 17907 26484 17973 26485
rect 17907 26420 17908 26484
rect 17972 26420 17973 26484
rect 17907 26419 17973 26420
rect 18091 26484 18157 26485
rect 18091 26420 18092 26484
rect 18156 26420 18157 26484
rect 18091 26419 18157 26420
rect 17539 23900 17605 23901
rect 17539 23836 17540 23900
rect 17604 23836 17605 23900
rect 17539 23835 17605 23836
rect 17723 23900 17789 23901
rect 17723 23836 17724 23900
rect 17788 23836 17789 23900
rect 17723 23835 17789 23836
rect 17542 23626 17602 23835
rect 17542 23566 17786 23626
rect 17539 23492 17605 23493
rect 17539 23428 17540 23492
rect 17604 23428 17605 23492
rect 17539 23427 17605 23428
rect 17542 22810 17602 23427
rect 17726 22949 17786 23566
rect 17910 23221 17970 26419
rect 18091 26348 18157 26349
rect 18091 26284 18092 26348
rect 18156 26346 18157 26348
rect 18278 26346 18338 29683
rect 18459 28252 18525 28253
rect 18459 28188 18460 28252
rect 18524 28188 18525 28252
rect 18459 28187 18525 28188
rect 18643 28252 18709 28253
rect 18643 28188 18644 28252
rect 18708 28188 18709 28252
rect 18643 28187 18709 28188
rect 18462 27573 18522 28187
rect 18459 27572 18525 27573
rect 18459 27508 18460 27572
rect 18524 27508 18525 27572
rect 18459 27507 18525 27508
rect 18459 27028 18525 27029
rect 18459 26964 18460 27028
rect 18524 26964 18525 27028
rect 18459 26963 18525 26964
rect 18156 26286 18338 26346
rect 18156 26284 18157 26286
rect 18091 26283 18157 26284
rect 18091 26076 18157 26077
rect 18091 26012 18092 26076
rect 18156 26012 18157 26076
rect 18091 26011 18157 26012
rect 17907 23220 17973 23221
rect 17907 23156 17908 23220
rect 17972 23156 17973 23220
rect 17907 23155 17973 23156
rect 17723 22948 17789 22949
rect 17723 22884 17724 22948
rect 17788 22884 17789 22948
rect 17723 22883 17789 22884
rect 17542 22750 17970 22810
rect 17723 22676 17789 22677
rect 17358 22614 17602 22674
rect 17355 21724 17421 21725
rect 17355 21660 17356 21724
rect 17420 21660 17421 21724
rect 17355 21659 17421 21660
rect 17171 21588 17237 21589
rect 17171 21524 17172 21588
rect 17236 21524 17237 21588
rect 17171 21523 17237 21524
rect 16308 20640 16316 20704
rect 16380 20640 16396 20704
rect 16460 20640 16476 20704
rect 16540 20640 16556 20704
rect 16620 20640 16628 20704
rect 16308 19616 16628 20640
rect 16308 19552 16316 19616
rect 16380 19552 16396 19616
rect 16460 19552 16476 19616
rect 16540 19552 16556 19616
rect 16620 19552 16628 19616
rect 15699 18868 15765 18869
rect 15699 18804 15700 18868
rect 15764 18804 15765 18868
rect 15699 18803 15765 18804
rect 15515 14108 15581 14109
rect 15515 14044 15516 14108
rect 15580 14044 15581 14108
rect 15515 14043 15581 14044
rect 15331 8940 15397 8941
rect 15331 8876 15332 8940
rect 15396 8876 15397 8940
rect 15331 8875 15397 8876
rect 14411 7444 14477 7445
rect 14411 7380 14412 7444
rect 14476 7380 14477 7444
rect 14411 7379 14477 7380
rect 14043 6900 14109 6901
rect 14043 6836 14044 6900
rect 14108 6836 14109 6900
rect 14043 6835 14109 6836
rect 13491 5132 13557 5133
rect 13491 5068 13492 5132
rect 13556 5068 13557 5132
rect 13491 5067 13557 5068
rect 12467 4864 12475 4928
rect 12539 4864 12555 4928
rect 12619 4864 12635 4928
rect 12699 4864 12715 4928
rect 12779 4864 12787 4928
rect 12467 3840 12787 4864
rect 15702 4725 15762 18803
rect 15886 10029 15946 19290
rect 16067 18868 16133 18869
rect 16067 18804 16068 18868
rect 16132 18804 16133 18868
rect 16067 18803 16133 18804
rect 16070 18597 16130 18803
rect 16067 18596 16133 18597
rect 16067 18532 16068 18596
rect 16132 18532 16133 18596
rect 16067 18531 16133 18532
rect 16308 18528 16628 19552
rect 16308 18464 16316 18528
rect 16380 18464 16396 18528
rect 16460 18464 16476 18528
rect 16540 18464 16556 18528
rect 16620 18464 16628 18528
rect 16308 17440 16628 18464
rect 16806 21390 17050 21450
rect 16806 18461 16866 21390
rect 16987 21180 17053 21181
rect 16987 21116 16988 21180
rect 17052 21116 17053 21180
rect 16987 21115 17053 21116
rect 16803 18460 16869 18461
rect 16803 18396 16804 18460
rect 16868 18396 16869 18460
rect 16803 18395 16869 18396
rect 16990 17917 17050 21115
rect 17174 20773 17234 21523
rect 17171 20772 17237 20773
rect 17171 20708 17172 20772
rect 17236 20708 17237 20772
rect 17171 20707 17237 20708
rect 17171 19956 17237 19957
rect 17171 19892 17172 19956
rect 17236 19892 17237 19956
rect 17171 19891 17237 19892
rect 16803 17916 16869 17917
rect 16803 17852 16804 17916
rect 16868 17852 16869 17916
rect 16803 17851 16869 17852
rect 16987 17916 17053 17917
rect 16987 17852 16988 17916
rect 17052 17852 17053 17916
rect 16987 17851 17053 17852
rect 16308 17376 16316 17440
rect 16380 17376 16396 17440
rect 16460 17376 16476 17440
rect 16540 17376 16556 17440
rect 16620 17376 16628 17440
rect 16067 16964 16133 16965
rect 16067 16900 16068 16964
rect 16132 16900 16133 16964
rect 16067 16899 16133 16900
rect 16070 15333 16130 16899
rect 16308 16352 16628 17376
rect 16308 16288 16316 16352
rect 16380 16288 16396 16352
rect 16460 16288 16476 16352
rect 16540 16288 16556 16352
rect 16620 16288 16628 16352
rect 16067 15332 16133 15333
rect 16067 15268 16068 15332
rect 16132 15268 16133 15332
rect 16067 15267 16133 15268
rect 16308 15264 16628 16288
rect 16806 15605 16866 17851
rect 17174 17781 17234 19891
rect 17358 18869 17418 21659
rect 17542 21589 17602 22614
rect 17723 22612 17724 22676
rect 17788 22612 17789 22676
rect 17723 22611 17789 22612
rect 17726 21861 17786 22611
rect 17910 21997 17970 22750
rect 17907 21996 17973 21997
rect 17907 21932 17908 21996
rect 17972 21932 17973 21996
rect 17907 21931 17973 21932
rect 17723 21860 17789 21861
rect 17723 21796 17724 21860
rect 17788 21796 17789 21860
rect 17723 21795 17789 21796
rect 17539 21588 17605 21589
rect 17539 21524 17540 21588
rect 17604 21524 17605 21588
rect 17539 21523 17605 21524
rect 17539 21452 17605 21453
rect 17539 21388 17540 21452
rect 17604 21388 17605 21452
rect 17539 21387 17605 21388
rect 17542 20909 17602 21387
rect 17539 20908 17605 20909
rect 17539 20844 17540 20908
rect 17604 20844 17605 20908
rect 17539 20843 17605 20844
rect 17355 18868 17421 18869
rect 17355 18804 17356 18868
rect 17420 18804 17421 18868
rect 17355 18803 17421 18804
rect 17171 17780 17237 17781
rect 17171 17716 17172 17780
rect 17236 17716 17237 17780
rect 17171 17715 17237 17716
rect 17171 17372 17237 17373
rect 17171 17308 17172 17372
rect 17236 17370 17237 17372
rect 17236 17310 17418 17370
rect 17236 17308 17237 17310
rect 17171 17307 17237 17308
rect 17358 16965 17418 17310
rect 17355 16964 17421 16965
rect 17355 16900 17356 16964
rect 17420 16900 17421 16964
rect 17355 16899 17421 16900
rect 16803 15604 16869 15605
rect 16803 15540 16804 15604
rect 16868 15540 16869 15604
rect 16803 15539 16869 15540
rect 16308 15200 16316 15264
rect 16380 15200 16396 15264
rect 16460 15200 16476 15264
rect 16540 15200 16556 15264
rect 16620 15200 16628 15264
rect 16308 14176 16628 15200
rect 16308 14112 16316 14176
rect 16380 14112 16396 14176
rect 16460 14112 16476 14176
rect 16540 14112 16556 14176
rect 16620 14112 16628 14176
rect 16308 13088 16628 14112
rect 16308 13024 16316 13088
rect 16380 13024 16396 13088
rect 16460 13024 16476 13088
rect 16540 13024 16556 13088
rect 16620 13024 16628 13088
rect 16308 12000 16628 13024
rect 16308 11936 16316 12000
rect 16380 11936 16396 12000
rect 16460 11936 16476 12000
rect 16540 11936 16556 12000
rect 16620 11936 16628 12000
rect 16308 10912 16628 11936
rect 16308 10848 16316 10912
rect 16380 10848 16396 10912
rect 16460 10848 16476 10912
rect 16540 10848 16556 10912
rect 16620 10848 16628 10912
rect 15883 10028 15949 10029
rect 15883 9964 15884 10028
rect 15948 9964 15949 10028
rect 15883 9963 15949 9964
rect 16308 9824 16628 10848
rect 16308 9760 16316 9824
rect 16380 9760 16396 9824
rect 16460 9760 16476 9824
rect 16540 9760 16556 9824
rect 16620 9760 16628 9824
rect 16308 8736 16628 9760
rect 16308 8672 16316 8736
rect 16380 8672 16396 8736
rect 16460 8672 16476 8736
rect 16540 8672 16556 8736
rect 16620 8672 16628 8736
rect 16308 7648 16628 8672
rect 17726 8669 17786 21795
rect 18094 21725 18154 26011
rect 18275 22948 18341 22949
rect 18275 22884 18276 22948
rect 18340 22884 18341 22948
rect 18275 22883 18341 22884
rect 18278 22541 18338 22883
rect 18275 22540 18341 22541
rect 18275 22476 18276 22540
rect 18340 22476 18341 22540
rect 18275 22475 18341 22476
rect 18091 21724 18157 21725
rect 18091 21660 18092 21724
rect 18156 21660 18157 21724
rect 18091 21659 18157 21660
rect 18278 19954 18338 22475
rect 18462 21725 18522 26963
rect 18646 26485 18706 28187
rect 18643 26484 18709 26485
rect 18643 26420 18644 26484
rect 18708 26420 18709 26484
rect 18643 26419 18709 26420
rect 18643 24988 18709 24989
rect 18643 24924 18644 24988
rect 18708 24924 18709 24988
rect 18643 24923 18709 24924
rect 18646 22949 18706 24923
rect 18830 23490 18890 30330
rect 19011 28660 19077 28661
rect 19011 28596 19012 28660
rect 19076 28596 19077 28660
rect 19011 28595 19077 28596
rect 19014 24445 19074 28595
rect 19198 27709 19258 30635
rect 19379 30292 19445 30293
rect 19379 30228 19380 30292
rect 19444 30228 19445 30292
rect 19379 30227 19445 30228
rect 19195 27708 19261 27709
rect 19195 27644 19196 27708
rect 19260 27644 19261 27708
rect 19195 27643 19261 27644
rect 19195 27572 19261 27573
rect 19195 27508 19196 27572
rect 19260 27508 19261 27572
rect 19195 27507 19261 27508
rect 19198 26482 19258 27507
rect 19382 26621 19442 30227
rect 19563 28932 19629 28933
rect 19563 28868 19564 28932
rect 19628 28868 19629 28932
rect 19563 28867 19629 28868
rect 19379 26620 19445 26621
rect 19379 26556 19380 26620
rect 19444 26556 19445 26620
rect 19379 26555 19445 26556
rect 19198 26422 19442 26482
rect 19195 25668 19261 25669
rect 19195 25604 19196 25668
rect 19260 25604 19261 25668
rect 19195 25603 19261 25604
rect 19011 24444 19077 24445
rect 19011 24380 19012 24444
rect 19076 24380 19077 24444
rect 19011 24379 19077 24380
rect 18830 23430 19074 23490
rect 18643 22948 18709 22949
rect 18643 22884 18644 22948
rect 18708 22884 18709 22948
rect 18643 22883 18709 22884
rect 18643 22268 18709 22269
rect 18643 22204 18644 22268
rect 18708 22266 18709 22268
rect 18708 22206 18890 22266
rect 18708 22204 18709 22206
rect 18643 22203 18709 22204
rect 18643 22132 18709 22133
rect 18643 22068 18644 22132
rect 18708 22068 18709 22132
rect 18643 22067 18709 22068
rect 18459 21724 18525 21725
rect 18459 21660 18460 21724
rect 18524 21660 18525 21724
rect 18459 21659 18525 21660
rect 18459 19956 18525 19957
rect 18459 19954 18460 19956
rect 18278 19894 18460 19954
rect 18459 19892 18460 19894
rect 18524 19892 18525 19956
rect 18459 19891 18525 19892
rect 18646 19549 18706 22067
rect 18830 21861 18890 22206
rect 18827 21860 18893 21861
rect 18827 21796 18828 21860
rect 18892 21796 18893 21860
rect 18827 21795 18893 21796
rect 19014 20093 19074 23430
rect 19198 20637 19258 25603
rect 19382 22269 19442 26422
rect 19566 25397 19626 28867
rect 19750 28661 19810 30771
rect 19934 30429 19994 32675
rect 20149 32128 20469 32688
rect 20667 32468 20733 32469
rect 20667 32404 20668 32468
rect 20732 32404 20733 32468
rect 20667 32403 20733 32404
rect 20149 32064 20157 32128
rect 20221 32064 20237 32128
rect 20301 32064 20317 32128
rect 20381 32064 20397 32128
rect 20461 32064 20469 32128
rect 20149 31040 20469 32064
rect 20149 30976 20157 31040
rect 20221 30976 20237 31040
rect 20301 30976 20317 31040
rect 20381 30976 20397 31040
rect 20461 30976 20469 31040
rect 19931 30428 19997 30429
rect 19931 30364 19932 30428
rect 19996 30364 19997 30428
rect 19931 30363 19997 30364
rect 20149 29952 20469 30976
rect 20149 29888 20157 29952
rect 20221 29888 20237 29952
rect 20301 29888 20317 29952
rect 20381 29888 20397 29952
rect 20461 29888 20469 29952
rect 19931 29204 19997 29205
rect 19931 29140 19932 29204
rect 19996 29140 19997 29204
rect 19931 29139 19997 29140
rect 19747 28660 19813 28661
rect 19747 28596 19748 28660
rect 19812 28596 19813 28660
rect 19747 28595 19813 28596
rect 19934 26754 19994 29139
rect 19750 26694 19994 26754
rect 20149 28864 20469 29888
rect 20149 28800 20157 28864
rect 20221 28800 20237 28864
rect 20301 28800 20317 28864
rect 20381 28800 20397 28864
rect 20461 28800 20469 28864
rect 20149 27776 20469 28800
rect 20670 28114 20730 32403
rect 20854 31770 20914 34715
rect 21955 31924 22021 31925
rect 21955 31860 21956 31924
rect 22020 31860 22021 31924
rect 21955 31859 22021 31860
rect 20854 31710 21650 31770
rect 21035 30428 21101 30429
rect 21035 30364 21036 30428
rect 21100 30364 21101 30428
rect 21035 30363 21101 30364
rect 20851 28796 20917 28797
rect 20851 28732 20852 28796
rect 20916 28732 20917 28796
rect 20851 28731 20917 28732
rect 20149 27712 20157 27776
rect 20221 27712 20237 27776
rect 20301 27712 20317 27776
rect 20381 27712 20397 27776
rect 20461 27712 20469 27776
rect 19563 25396 19629 25397
rect 19563 25332 19564 25396
rect 19628 25332 19629 25396
rect 19563 25331 19629 25332
rect 19563 24444 19629 24445
rect 19563 24380 19564 24444
rect 19628 24380 19629 24444
rect 19563 24379 19629 24380
rect 19379 22268 19445 22269
rect 19379 22204 19380 22268
rect 19444 22204 19445 22268
rect 19379 22203 19445 22204
rect 19379 21724 19445 21725
rect 19379 21660 19380 21724
rect 19444 21660 19445 21724
rect 19379 21659 19445 21660
rect 19382 20906 19442 21659
rect 19566 21181 19626 24379
rect 19750 23493 19810 26694
rect 20149 26688 20469 27712
rect 20149 26624 20157 26688
rect 20221 26624 20237 26688
rect 20301 26624 20317 26688
rect 20381 26624 20397 26688
rect 20461 26624 20469 26688
rect 19931 26620 19997 26621
rect 19931 26556 19932 26620
rect 19996 26556 19997 26620
rect 19931 26555 19997 26556
rect 19934 25941 19994 26555
rect 19931 25940 19997 25941
rect 19931 25876 19932 25940
rect 19996 25876 19997 25940
rect 19931 25875 19997 25876
rect 19747 23492 19813 23493
rect 19747 23428 19748 23492
rect 19812 23428 19813 23492
rect 19747 23427 19813 23428
rect 19563 21180 19629 21181
rect 19563 21116 19564 21180
rect 19628 21116 19629 21180
rect 19563 21115 19629 21116
rect 19382 20846 19626 20906
rect 19195 20636 19261 20637
rect 19195 20572 19196 20636
rect 19260 20572 19261 20636
rect 19195 20571 19261 20572
rect 19011 20092 19077 20093
rect 19011 20028 19012 20092
rect 19076 20028 19077 20092
rect 19011 20027 19077 20028
rect 19379 20092 19445 20093
rect 19379 20028 19380 20092
rect 19444 20028 19445 20092
rect 19379 20027 19445 20028
rect 19382 19549 19442 20027
rect 18643 19548 18709 19549
rect 18643 19484 18644 19548
rect 18708 19484 18709 19548
rect 18643 19483 18709 19484
rect 19379 19548 19445 19549
rect 19379 19484 19380 19548
rect 19444 19484 19445 19548
rect 19379 19483 19445 19484
rect 17907 15332 17973 15333
rect 17907 15268 17908 15332
rect 17972 15268 17973 15332
rect 17907 15267 17973 15268
rect 17910 12341 17970 15267
rect 17907 12340 17973 12341
rect 17907 12276 17908 12340
rect 17972 12276 17973 12340
rect 17907 12275 17973 12276
rect 17723 8668 17789 8669
rect 17723 8604 17724 8668
rect 17788 8604 17789 8668
rect 17723 8603 17789 8604
rect 16308 7584 16316 7648
rect 16380 7584 16396 7648
rect 16460 7584 16476 7648
rect 16540 7584 16556 7648
rect 16620 7584 16628 7648
rect 16308 6560 16628 7584
rect 18646 6765 18706 19483
rect 19379 19412 19445 19413
rect 19379 19348 19380 19412
rect 19444 19348 19445 19412
rect 19379 19347 19445 19348
rect 18827 19140 18893 19141
rect 18827 19076 18828 19140
rect 18892 19076 18893 19140
rect 18827 19075 18893 19076
rect 18830 12205 18890 19075
rect 19011 16284 19077 16285
rect 19011 16220 19012 16284
rect 19076 16220 19077 16284
rect 19011 16219 19077 16220
rect 19014 13973 19074 16219
rect 19011 13972 19077 13973
rect 19011 13908 19012 13972
rect 19076 13908 19077 13972
rect 19011 13907 19077 13908
rect 18827 12204 18893 12205
rect 18827 12140 18828 12204
rect 18892 12140 18893 12204
rect 18827 12139 18893 12140
rect 19382 8397 19442 19347
rect 19566 18730 19626 20846
rect 19934 19549 19994 25875
rect 20149 25600 20469 26624
rect 20532 28054 20730 28114
rect 20532 26618 20592 28054
rect 20667 27844 20733 27845
rect 20667 27780 20668 27844
rect 20732 27780 20733 27844
rect 20667 27779 20733 27780
rect 20670 26757 20730 27779
rect 20854 27709 20914 28731
rect 20851 27708 20917 27709
rect 20851 27644 20852 27708
rect 20916 27644 20917 27708
rect 20851 27643 20917 27644
rect 20667 26756 20733 26757
rect 20667 26692 20668 26756
rect 20732 26692 20733 26756
rect 20667 26691 20733 26692
rect 20532 26558 20914 26618
rect 20667 26484 20733 26485
rect 20667 26420 20668 26484
rect 20732 26420 20733 26484
rect 20667 26419 20733 26420
rect 20670 26210 20730 26419
rect 20854 26349 20914 26558
rect 20851 26348 20917 26349
rect 20851 26284 20852 26348
rect 20916 26284 20917 26348
rect 20851 26283 20917 26284
rect 20149 25536 20157 25600
rect 20221 25536 20237 25600
rect 20301 25536 20317 25600
rect 20381 25536 20397 25600
rect 20461 25536 20469 25600
rect 20149 24512 20469 25536
rect 20532 26150 20730 26210
rect 20851 26212 20917 26213
rect 20532 24989 20592 26150
rect 20851 26148 20852 26212
rect 20916 26148 20917 26212
rect 20851 26147 20917 26148
rect 20667 26076 20733 26077
rect 20667 26012 20668 26076
rect 20732 26012 20733 26076
rect 20667 26011 20733 26012
rect 20670 25533 20730 26011
rect 20667 25532 20733 25533
rect 20667 25468 20668 25532
rect 20732 25468 20733 25532
rect 20667 25467 20733 25468
rect 20667 25124 20733 25125
rect 20667 25060 20668 25124
rect 20732 25060 20733 25124
rect 20667 25059 20733 25060
rect 20529 24988 20595 24989
rect 20529 24924 20530 24988
rect 20594 24924 20595 24988
rect 20529 24923 20595 24924
rect 20149 24448 20157 24512
rect 20221 24448 20237 24512
rect 20301 24448 20317 24512
rect 20381 24448 20397 24512
rect 20461 24448 20469 24512
rect 20149 23424 20469 24448
rect 20670 23493 20730 25059
rect 20667 23492 20733 23493
rect 20667 23428 20668 23492
rect 20732 23428 20733 23492
rect 20667 23427 20733 23428
rect 20149 23360 20157 23424
rect 20221 23360 20237 23424
rect 20301 23360 20317 23424
rect 20381 23360 20397 23424
rect 20461 23360 20469 23424
rect 20149 22336 20469 23360
rect 20854 23357 20914 26147
rect 20667 23356 20733 23357
rect 20667 23292 20668 23356
rect 20732 23292 20733 23356
rect 20667 23291 20733 23292
rect 20851 23356 20917 23357
rect 20851 23292 20852 23356
rect 20916 23292 20917 23356
rect 20851 23291 20917 23292
rect 20670 22538 20730 23291
rect 21038 22677 21098 30363
rect 21403 29476 21469 29477
rect 21403 29412 21404 29476
rect 21468 29412 21469 29476
rect 21403 29411 21469 29412
rect 21219 29340 21285 29341
rect 21219 29276 21220 29340
rect 21284 29276 21285 29340
rect 21219 29275 21285 29276
rect 21222 27573 21282 29275
rect 21219 27572 21285 27573
rect 21219 27508 21220 27572
rect 21284 27508 21285 27572
rect 21219 27507 21285 27508
rect 21219 27436 21285 27437
rect 21219 27372 21220 27436
rect 21284 27372 21285 27436
rect 21219 27371 21285 27372
rect 21222 26213 21282 27371
rect 21219 26212 21285 26213
rect 21219 26148 21220 26212
rect 21284 26148 21285 26212
rect 21219 26147 21285 26148
rect 21219 25940 21285 25941
rect 21219 25876 21220 25940
rect 21284 25876 21285 25940
rect 21219 25875 21285 25876
rect 21035 22676 21101 22677
rect 21035 22612 21036 22676
rect 21100 22612 21101 22676
rect 21035 22611 21101 22612
rect 21035 22540 21101 22541
rect 21035 22538 21036 22540
rect 20670 22478 21036 22538
rect 21035 22476 21036 22478
rect 21100 22476 21101 22540
rect 21035 22475 21101 22476
rect 20149 22272 20157 22336
rect 20221 22272 20237 22336
rect 20301 22272 20317 22336
rect 20381 22272 20397 22336
rect 20461 22272 20469 22336
rect 20149 21248 20469 22272
rect 20667 22268 20733 22269
rect 20667 22204 20668 22268
rect 20732 22204 20733 22268
rect 20667 22203 20733 22204
rect 20670 21450 20730 22203
rect 20149 21184 20157 21248
rect 20221 21184 20237 21248
rect 20301 21184 20317 21248
rect 20381 21184 20397 21248
rect 20461 21184 20469 21248
rect 20149 20160 20469 21184
rect 20149 20096 20157 20160
rect 20221 20096 20237 20160
rect 20301 20096 20317 20160
rect 20381 20096 20397 20160
rect 20461 20096 20469 20160
rect 19931 19548 19997 19549
rect 19931 19484 19932 19548
rect 19996 19484 19997 19548
rect 19931 19483 19997 19484
rect 20149 19072 20469 20096
rect 20532 21390 20730 21450
rect 20532 19413 20592 21390
rect 20667 21180 20733 21181
rect 20667 21116 20668 21180
rect 20732 21116 20733 21180
rect 20667 21115 20733 21116
rect 20529 19412 20595 19413
rect 20529 19348 20530 19412
rect 20594 19348 20595 19412
rect 20529 19347 20595 19348
rect 20149 19008 20157 19072
rect 20221 19008 20237 19072
rect 20301 19008 20317 19072
rect 20381 19008 20397 19072
rect 20461 19008 20469 19072
rect 19747 18732 19813 18733
rect 19747 18730 19748 18732
rect 19566 18670 19748 18730
rect 19747 18668 19748 18670
rect 19812 18668 19813 18732
rect 19747 18667 19813 18668
rect 20149 17984 20469 19008
rect 20149 17920 20157 17984
rect 20221 17920 20237 17984
rect 20301 17920 20317 17984
rect 20381 17920 20397 17984
rect 20461 17920 20469 17984
rect 20149 16896 20469 17920
rect 20149 16832 20157 16896
rect 20221 16832 20237 16896
rect 20301 16832 20317 16896
rect 20381 16832 20397 16896
rect 20461 16832 20469 16896
rect 20149 15808 20469 16832
rect 20149 15744 20157 15808
rect 20221 15744 20237 15808
rect 20301 15744 20317 15808
rect 20381 15744 20397 15808
rect 20461 15744 20469 15808
rect 20149 14720 20469 15744
rect 20149 14656 20157 14720
rect 20221 14656 20237 14720
rect 20301 14656 20317 14720
rect 20381 14656 20397 14720
rect 20461 14656 20469 14720
rect 19563 14652 19629 14653
rect 19563 14588 19564 14652
rect 19628 14588 19629 14652
rect 19563 14587 19629 14588
rect 19566 12069 19626 14587
rect 20149 13632 20469 14656
rect 20149 13568 20157 13632
rect 20221 13568 20237 13632
rect 20301 13568 20317 13632
rect 20381 13568 20397 13632
rect 20461 13568 20469 13632
rect 20149 12544 20469 13568
rect 20149 12480 20157 12544
rect 20221 12480 20237 12544
rect 20301 12480 20317 12544
rect 20381 12480 20397 12544
rect 20461 12480 20469 12544
rect 19563 12068 19629 12069
rect 19563 12004 19564 12068
rect 19628 12004 19629 12068
rect 19563 12003 19629 12004
rect 20149 11456 20469 12480
rect 20670 11797 20730 21115
rect 21222 17917 21282 25875
rect 21406 24989 21466 29411
rect 21590 29341 21650 31710
rect 21771 29748 21837 29749
rect 21771 29684 21772 29748
rect 21836 29684 21837 29748
rect 21771 29683 21837 29684
rect 21587 29340 21653 29341
rect 21587 29276 21588 29340
rect 21652 29276 21653 29340
rect 21587 29275 21653 29276
rect 21774 27845 21834 29683
rect 21958 29341 22018 31859
rect 21955 29340 22021 29341
rect 21955 29276 21956 29340
rect 22020 29276 22021 29340
rect 21955 29275 22021 29276
rect 21955 29204 22021 29205
rect 21955 29140 21956 29204
rect 22020 29140 22021 29204
rect 21955 29139 22021 29140
rect 21958 28525 22018 29139
rect 21955 28524 22021 28525
rect 21955 28460 21956 28524
rect 22020 28460 22021 28524
rect 21955 28459 22021 28460
rect 21587 27844 21653 27845
rect 21587 27780 21588 27844
rect 21652 27780 21653 27844
rect 21587 27779 21653 27780
rect 21771 27844 21837 27845
rect 21771 27780 21772 27844
rect 21836 27780 21837 27844
rect 21771 27779 21837 27780
rect 21403 24988 21469 24989
rect 21403 24924 21404 24988
rect 21468 24924 21469 24988
rect 21403 24923 21469 24924
rect 21590 24445 21650 27779
rect 21771 26620 21837 26621
rect 21771 26556 21772 26620
rect 21836 26556 21837 26620
rect 21771 26555 21837 26556
rect 21774 24989 21834 26555
rect 21771 24988 21837 24989
rect 21771 24924 21772 24988
rect 21836 24924 21837 24988
rect 21771 24923 21837 24924
rect 21403 24444 21469 24445
rect 21403 24380 21404 24444
rect 21468 24380 21469 24444
rect 21403 24379 21469 24380
rect 21587 24444 21653 24445
rect 21587 24380 21588 24444
rect 21652 24380 21653 24444
rect 21587 24379 21653 24380
rect 21406 22677 21466 24379
rect 21590 23490 21650 24379
rect 21774 24173 21834 24923
rect 21771 24172 21837 24173
rect 21771 24108 21772 24172
rect 21836 24108 21837 24172
rect 21771 24107 21837 24108
rect 21590 23430 21834 23490
rect 21403 22676 21469 22677
rect 21403 22612 21404 22676
rect 21468 22612 21469 22676
rect 21403 22611 21469 22612
rect 21587 22540 21653 22541
rect 21587 22476 21588 22540
rect 21652 22476 21653 22540
rect 21587 22475 21653 22476
rect 21590 21858 21650 22475
rect 21774 22402 21834 23430
rect 21958 22541 22018 28459
rect 22142 27845 22202 34851
rect 26555 34236 26621 34237
rect 26555 34172 26556 34236
rect 26620 34172 26621 34236
rect 26555 34171 26621 34172
rect 23795 33828 23861 33829
rect 23795 33764 23796 33828
rect 23860 33764 23861 33828
rect 23795 33763 23861 33764
rect 22323 32604 22389 32605
rect 22323 32540 22324 32604
rect 22388 32540 22389 32604
rect 22323 32539 22389 32540
rect 22326 28253 22386 32539
rect 22507 31516 22573 31517
rect 22507 31452 22508 31516
rect 22572 31452 22573 31516
rect 22507 31451 22573 31452
rect 22510 29613 22570 31451
rect 22691 31244 22757 31245
rect 22691 31180 22692 31244
rect 22756 31180 22757 31244
rect 22691 31179 22757 31180
rect 22507 29612 22573 29613
rect 22507 29548 22508 29612
rect 22572 29548 22573 29612
rect 22507 29547 22573 29548
rect 22323 28252 22389 28253
rect 22323 28188 22324 28252
rect 22388 28188 22389 28252
rect 22323 28187 22389 28188
rect 22139 27844 22205 27845
rect 22139 27780 22140 27844
rect 22204 27780 22205 27844
rect 22139 27779 22205 27780
rect 22139 27708 22205 27709
rect 22139 27644 22140 27708
rect 22204 27644 22205 27708
rect 22139 27643 22205 27644
rect 21955 22540 22021 22541
rect 21955 22476 21956 22540
rect 22020 22476 22021 22540
rect 21955 22475 22021 22476
rect 22142 22405 22202 27643
rect 22139 22404 22205 22405
rect 21774 22342 22018 22402
rect 21771 21860 21837 21861
rect 21771 21858 21772 21860
rect 21590 21798 21772 21858
rect 21771 21796 21772 21798
rect 21836 21796 21837 21860
rect 21771 21795 21837 21796
rect 21587 19140 21653 19141
rect 21587 19076 21588 19140
rect 21652 19138 21653 19140
rect 21958 19138 22018 22342
rect 22139 22340 22140 22404
rect 22204 22340 22205 22404
rect 22139 22339 22205 22340
rect 22326 21181 22386 28187
rect 22510 27709 22570 29547
rect 22694 28933 22754 31179
rect 23427 30564 23493 30565
rect 23427 30500 23428 30564
rect 23492 30500 23493 30564
rect 23427 30499 23493 30500
rect 22875 30292 22941 30293
rect 22875 30228 22876 30292
rect 22940 30228 22941 30292
rect 22875 30227 22941 30228
rect 22691 28932 22757 28933
rect 22691 28868 22692 28932
rect 22756 28868 22757 28932
rect 22691 28867 22757 28868
rect 22878 28658 22938 30227
rect 23059 29476 23125 29477
rect 23059 29412 23060 29476
rect 23124 29412 23125 29476
rect 23059 29411 23125 29412
rect 22694 28598 22938 28658
rect 22694 28253 22754 28598
rect 22875 28524 22941 28525
rect 22875 28460 22876 28524
rect 22940 28460 22941 28524
rect 22875 28459 22941 28460
rect 22691 28252 22757 28253
rect 22691 28188 22692 28252
rect 22756 28188 22757 28252
rect 22691 28187 22757 28188
rect 22691 27844 22757 27845
rect 22691 27780 22692 27844
rect 22756 27780 22757 27844
rect 22691 27779 22757 27780
rect 22507 27708 22573 27709
rect 22507 27644 22508 27708
rect 22572 27644 22573 27708
rect 22507 27643 22573 27644
rect 22507 27572 22573 27573
rect 22507 27508 22508 27572
rect 22572 27508 22573 27572
rect 22507 27507 22573 27508
rect 22510 23765 22570 27507
rect 22694 24989 22754 27779
rect 22691 24988 22757 24989
rect 22691 24924 22692 24988
rect 22756 24924 22757 24988
rect 22691 24923 22757 24924
rect 22878 24309 22938 28459
rect 23062 26213 23122 29411
rect 23243 29340 23309 29341
rect 23243 29276 23244 29340
rect 23308 29276 23309 29340
rect 23243 29275 23309 29276
rect 23246 27573 23306 29275
rect 23430 27573 23490 30499
rect 23611 29340 23677 29341
rect 23611 29276 23612 29340
rect 23676 29276 23677 29340
rect 23611 29275 23677 29276
rect 23614 28253 23674 29275
rect 23611 28252 23677 28253
rect 23611 28188 23612 28252
rect 23676 28188 23677 28252
rect 23611 28187 23677 28188
rect 23243 27572 23309 27573
rect 23243 27508 23244 27572
rect 23308 27508 23309 27572
rect 23243 27507 23309 27508
rect 23427 27572 23493 27573
rect 23427 27508 23428 27572
rect 23492 27508 23493 27572
rect 23427 27507 23493 27508
rect 23611 27572 23677 27573
rect 23611 27508 23612 27572
rect 23676 27508 23677 27572
rect 23611 27507 23677 27508
rect 23614 27298 23674 27507
rect 23430 27238 23674 27298
rect 23243 27028 23309 27029
rect 23243 26964 23244 27028
rect 23308 26964 23309 27028
rect 23243 26963 23309 26964
rect 23059 26212 23125 26213
rect 23059 26148 23060 26212
rect 23124 26148 23125 26212
rect 23059 26147 23125 26148
rect 23059 26076 23125 26077
rect 23059 26012 23060 26076
rect 23124 26012 23125 26076
rect 23059 26011 23125 26012
rect 22875 24308 22941 24309
rect 22875 24244 22876 24308
rect 22940 24244 22941 24308
rect 22875 24243 22941 24244
rect 22691 24172 22757 24173
rect 22691 24108 22692 24172
rect 22756 24108 22757 24172
rect 22691 24107 22757 24108
rect 22507 23764 22573 23765
rect 22507 23700 22508 23764
rect 22572 23700 22573 23764
rect 22507 23699 22573 23700
rect 22694 21861 22754 24107
rect 22691 21860 22757 21861
rect 22691 21796 22692 21860
rect 22756 21796 22757 21860
rect 22691 21795 22757 21796
rect 22323 21180 22389 21181
rect 22323 21116 22324 21180
rect 22388 21116 22389 21180
rect 22323 21115 22389 21116
rect 23062 20501 23122 26011
rect 23059 20500 23125 20501
rect 23059 20436 23060 20500
rect 23124 20436 23125 20500
rect 23059 20435 23125 20436
rect 23246 19957 23306 26963
rect 23430 22813 23490 27238
rect 23611 27164 23677 27165
rect 23611 27100 23612 27164
rect 23676 27100 23677 27164
rect 23611 27099 23677 27100
rect 23614 25397 23674 27099
rect 23798 26621 23858 33763
rect 23990 32672 24310 32688
rect 23990 32608 23998 32672
rect 24062 32608 24078 32672
rect 24142 32608 24158 32672
rect 24222 32608 24238 32672
rect 24302 32608 24310 32672
rect 23990 31584 24310 32608
rect 26187 32060 26253 32061
rect 26187 31996 26188 32060
rect 26252 31996 26253 32060
rect 26187 31995 26253 31996
rect 25451 31788 25517 31789
rect 25451 31724 25452 31788
rect 25516 31724 25517 31788
rect 25451 31723 25517 31724
rect 24531 31652 24597 31653
rect 24531 31588 24532 31652
rect 24596 31588 24597 31652
rect 24531 31587 24597 31588
rect 23990 31520 23998 31584
rect 24062 31520 24078 31584
rect 24142 31520 24158 31584
rect 24222 31520 24238 31584
rect 24302 31520 24310 31584
rect 23990 30496 24310 31520
rect 23990 30432 23998 30496
rect 24062 30432 24078 30496
rect 24142 30432 24158 30496
rect 24222 30432 24238 30496
rect 24302 30432 24310 30496
rect 23990 29408 24310 30432
rect 23990 29344 23998 29408
rect 24062 29344 24078 29408
rect 24142 29344 24158 29408
rect 24222 29344 24238 29408
rect 24302 29344 24310 29408
rect 23990 28320 24310 29344
rect 24534 28522 24594 31587
rect 25267 31108 25333 31109
rect 25267 31044 25268 31108
rect 25332 31044 25333 31108
rect 25267 31043 25333 31044
rect 25083 30156 25149 30157
rect 25083 30154 25084 30156
rect 23990 28256 23998 28320
rect 24062 28256 24078 28320
rect 24142 28256 24158 28320
rect 24222 28256 24238 28320
rect 24302 28256 24310 28320
rect 23990 27232 24310 28256
rect 23990 27168 23998 27232
rect 24062 27168 24078 27232
rect 24142 27168 24158 27232
rect 24222 27168 24238 27232
rect 24302 27168 24310 27232
rect 23795 26620 23861 26621
rect 23795 26556 23796 26620
rect 23860 26556 23861 26620
rect 23795 26555 23861 26556
rect 23795 26212 23861 26213
rect 23795 26148 23796 26212
rect 23860 26148 23861 26212
rect 23795 26147 23861 26148
rect 23611 25396 23677 25397
rect 23611 25332 23612 25396
rect 23676 25332 23677 25396
rect 23611 25331 23677 25332
rect 23611 24988 23677 24989
rect 23611 24924 23612 24988
rect 23676 24924 23677 24988
rect 23611 24923 23677 24924
rect 23614 22949 23674 24923
rect 23798 23901 23858 26147
rect 23990 26144 24310 27168
rect 23990 26080 23998 26144
rect 24062 26080 24078 26144
rect 24142 26080 24158 26144
rect 24222 26080 24238 26144
rect 24302 26080 24310 26144
rect 23990 25056 24310 26080
rect 24396 28462 24594 28522
rect 24718 30094 25084 30154
rect 24396 25941 24456 28462
rect 24531 28388 24597 28389
rect 24531 28324 24532 28388
rect 24596 28324 24597 28388
rect 24531 28323 24597 28324
rect 24393 25940 24459 25941
rect 24393 25876 24394 25940
rect 24458 25876 24459 25940
rect 24393 25875 24459 25876
rect 24534 25397 24594 28323
rect 24718 27573 24778 30094
rect 25083 30092 25084 30094
rect 25148 30092 25149 30156
rect 25083 30091 25149 30092
rect 25083 29748 25149 29749
rect 25083 29684 25084 29748
rect 25148 29684 25149 29748
rect 25083 29683 25149 29684
rect 24899 29068 24965 29069
rect 24899 29004 24900 29068
rect 24964 29004 24965 29068
rect 24899 29003 24965 29004
rect 24902 28389 24962 29003
rect 25086 28389 25146 29683
rect 24899 28388 24965 28389
rect 24899 28324 24900 28388
rect 24964 28324 24965 28388
rect 24899 28323 24965 28324
rect 25083 28388 25149 28389
rect 25083 28324 25084 28388
rect 25148 28324 25149 28388
rect 25083 28323 25149 28324
rect 24899 27844 24965 27845
rect 24899 27780 24900 27844
rect 24964 27780 24965 27844
rect 24899 27779 24965 27780
rect 24715 27572 24781 27573
rect 24715 27508 24716 27572
rect 24780 27508 24781 27572
rect 24715 27507 24781 27508
rect 24902 26893 24962 27779
rect 25086 27437 25146 28323
rect 25270 27845 25330 31043
rect 25454 29749 25514 31723
rect 26003 31652 26069 31653
rect 26003 31588 26004 31652
rect 26068 31588 26069 31652
rect 26003 31587 26069 31588
rect 25819 30836 25885 30837
rect 25819 30772 25820 30836
rect 25884 30772 25885 30836
rect 25819 30771 25885 30772
rect 25635 30156 25701 30157
rect 25635 30092 25636 30156
rect 25700 30092 25701 30156
rect 25635 30091 25701 30092
rect 25451 29748 25517 29749
rect 25451 29684 25452 29748
rect 25516 29684 25517 29748
rect 25451 29683 25517 29684
rect 25638 29477 25698 30091
rect 25451 29476 25517 29477
rect 25451 29412 25452 29476
rect 25516 29412 25517 29476
rect 25451 29411 25517 29412
rect 25635 29476 25701 29477
rect 25635 29412 25636 29476
rect 25700 29412 25701 29476
rect 25635 29411 25701 29412
rect 25267 27844 25333 27845
rect 25267 27780 25268 27844
rect 25332 27780 25333 27844
rect 25267 27779 25333 27780
rect 25083 27436 25149 27437
rect 25083 27372 25084 27436
rect 25148 27372 25149 27436
rect 25083 27371 25149 27372
rect 25083 27164 25149 27165
rect 25083 27100 25084 27164
rect 25148 27100 25149 27164
rect 25083 27099 25149 27100
rect 24899 26892 24965 26893
rect 24899 26828 24900 26892
rect 24964 26828 24965 26892
rect 24899 26827 24965 26828
rect 24715 26620 24781 26621
rect 24715 26556 24716 26620
rect 24780 26618 24781 26620
rect 24780 26558 24962 26618
rect 24780 26556 24781 26558
rect 24715 26555 24781 26556
rect 24902 26349 24962 26558
rect 24715 26348 24781 26349
rect 24715 26284 24716 26348
rect 24780 26284 24781 26348
rect 24715 26283 24781 26284
rect 24899 26348 24965 26349
rect 24899 26284 24900 26348
rect 24964 26284 24965 26348
rect 24899 26283 24965 26284
rect 24531 25396 24597 25397
rect 24531 25332 24532 25396
rect 24596 25332 24597 25396
rect 24531 25331 24597 25332
rect 23990 24992 23998 25056
rect 24062 24992 24078 25056
rect 24142 24992 24158 25056
rect 24222 24992 24238 25056
rect 24302 24992 24310 25056
rect 23990 23968 24310 24992
rect 23990 23904 23998 23968
rect 24062 23904 24078 23968
rect 24142 23904 24158 23968
rect 24222 23904 24238 23968
rect 24302 23904 24310 23968
rect 23795 23900 23861 23901
rect 23795 23836 23796 23900
rect 23860 23836 23861 23900
rect 23795 23835 23861 23836
rect 23611 22948 23677 22949
rect 23611 22884 23612 22948
rect 23676 22884 23677 22948
rect 23611 22883 23677 22884
rect 23990 22880 24310 23904
rect 24531 23492 24597 23493
rect 24531 23428 24532 23492
rect 24596 23428 24597 23492
rect 24531 23427 24597 23428
rect 23990 22816 23998 22880
rect 24062 22816 24078 22880
rect 24142 22816 24158 22880
rect 24222 22816 24238 22880
rect 24302 22816 24310 22880
rect 23427 22812 23493 22813
rect 23427 22748 23428 22812
rect 23492 22748 23493 22812
rect 23427 22747 23493 22748
rect 23990 21792 24310 22816
rect 23990 21728 23998 21792
rect 24062 21728 24078 21792
rect 24142 21728 24158 21792
rect 24222 21728 24238 21792
rect 24302 21728 24310 21792
rect 23990 20704 24310 21728
rect 23990 20640 23998 20704
rect 24062 20640 24078 20704
rect 24142 20640 24158 20704
rect 24222 20640 24238 20704
rect 24302 20640 24310 20704
rect 23059 19956 23125 19957
rect 23059 19892 23060 19956
rect 23124 19892 23125 19956
rect 23059 19891 23125 19892
rect 23243 19956 23309 19957
rect 23243 19892 23244 19956
rect 23308 19892 23309 19956
rect 23243 19891 23309 19892
rect 21652 19078 22018 19138
rect 21652 19076 21653 19078
rect 21587 19075 21653 19076
rect 21955 18868 22021 18869
rect 21955 18804 21956 18868
rect 22020 18804 22021 18868
rect 21955 18803 22021 18804
rect 21403 18732 21469 18733
rect 21403 18668 21404 18732
rect 21468 18668 21469 18732
rect 21403 18667 21469 18668
rect 21219 17916 21285 17917
rect 21219 17852 21220 17916
rect 21284 17852 21285 17916
rect 21219 17851 21285 17852
rect 21406 15333 21466 18667
rect 21587 18596 21653 18597
rect 21587 18532 21588 18596
rect 21652 18532 21653 18596
rect 21587 18531 21653 18532
rect 21403 15332 21469 15333
rect 21403 15268 21404 15332
rect 21468 15268 21469 15332
rect 21403 15267 21469 15268
rect 21403 15196 21469 15197
rect 21403 15132 21404 15196
rect 21468 15132 21469 15196
rect 21403 15131 21469 15132
rect 20851 14788 20917 14789
rect 20851 14724 20852 14788
rect 20916 14724 20917 14788
rect 20851 14723 20917 14724
rect 20854 13837 20914 14723
rect 20851 13836 20917 13837
rect 20851 13772 20852 13836
rect 20916 13772 20917 13836
rect 20851 13771 20917 13772
rect 20667 11796 20733 11797
rect 20667 11732 20668 11796
rect 20732 11732 20733 11796
rect 20667 11731 20733 11732
rect 20149 11392 20157 11456
rect 20221 11392 20237 11456
rect 20301 11392 20317 11456
rect 20381 11392 20397 11456
rect 20461 11392 20469 11456
rect 20149 10368 20469 11392
rect 20854 10709 20914 13771
rect 21035 13564 21101 13565
rect 21035 13500 21036 13564
rect 21100 13500 21101 13564
rect 21035 13499 21101 13500
rect 20851 10708 20917 10709
rect 20851 10644 20852 10708
rect 20916 10644 20917 10708
rect 20851 10643 20917 10644
rect 20149 10304 20157 10368
rect 20221 10304 20237 10368
rect 20301 10304 20317 10368
rect 20381 10304 20397 10368
rect 20461 10304 20469 10368
rect 20149 9280 20469 10304
rect 20149 9216 20157 9280
rect 20221 9216 20237 9280
rect 20301 9216 20317 9280
rect 20381 9216 20397 9280
rect 20461 9216 20469 9280
rect 19379 8396 19445 8397
rect 19379 8332 19380 8396
rect 19444 8332 19445 8396
rect 19379 8331 19445 8332
rect 20149 8192 20469 9216
rect 20149 8128 20157 8192
rect 20221 8128 20237 8192
rect 20301 8128 20317 8192
rect 20381 8128 20397 8192
rect 20461 8128 20469 8192
rect 20149 7104 20469 8128
rect 21038 7989 21098 13499
rect 21406 12613 21466 15131
rect 21590 14245 21650 18531
rect 21587 14244 21653 14245
rect 21587 14180 21588 14244
rect 21652 14180 21653 14244
rect 21587 14179 21653 14180
rect 21958 13157 22018 18803
rect 23062 14381 23122 19891
rect 23990 19616 24310 20640
rect 23990 19552 23998 19616
rect 24062 19552 24078 19616
rect 24142 19552 24158 19616
rect 24222 19552 24238 19616
rect 24302 19552 24310 19616
rect 23990 18528 24310 19552
rect 23990 18464 23998 18528
rect 24062 18464 24078 18528
rect 24142 18464 24158 18528
rect 24222 18464 24238 18528
rect 24302 18464 24310 18528
rect 23990 17440 24310 18464
rect 23990 17376 23998 17440
rect 24062 17376 24078 17440
rect 24142 17376 24158 17440
rect 24222 17376 24238 17440
rect 24302 17376 24310 17440
rect 23795 16828 23861 16829
rect 23795 16764 23796 16828
rect 23860 16764 23861 16828
rect 23795 16763 23861 16764
rect 23611 16692 23677 16693
rect 23611 16628 23612 16692
rect 23676 16628 23677 16692
rect 23611 16627 23677 16628
rect 23059 14380 23125 14381
rect 23059 14316 23060 14380
rect 23124 14316 23125 14380
rect 23059 14315 23125 14316
rect 21955 13156 22021 13157
rect 21955 13092 21956 13156
rect 22020 13092 22021 13156
rect 21955 13091 22021 13092
rect 21403 12612 21469 12613
rect 21403 12548 21404 12612
rect 21468 12548 21469 12612
rect 21403 12547 21469 12548
rect 23614 10709 23674 16627
rect 23798 12885 23858 16763
rect 23990 16352 24310 17376
rect 23990 16288 23998 16352
rect 24062 16288 24078 16352
rect 24142 16288 24158 16352
rect 24222 16288 24238 16352
rect 24302 16288 24310 16352
rect 23990 15264 24310 16288
rect 24534 15469 24594 23427
rect 24718 22813 24778 26283
rect 24899 26076 24965 26077
rect 24899 26012 24900 26076
rect 24964 26012 24965 26076
rect 24899 26011 24965 26012
rect 24715 22812 24781 22813
rect 24715 22748 24716 22812
rect 24780 22748 24781 22812
rect 24715 22747 24781 22748
rect 24902 19821 24962 26011
rect 25086 25805 25146 27099
rect 25083 25804 25149 25805
rect 25083 25740 25084 25804
rect 25148 25740 25149 25804
rect 25083 25739 25149 25740
rect 25086 24989 25146 25739
rect 25270 25533 25330 27779
rect 25454 26349 25514 29411
rect 25822 28253 25882 30771
rect 26006 29477 26066 31587
rect 26003 29476 26069 29477
rect 26003 29412 26004 29476
rect 26068 29412 26069 29476
rect 26003 29411 26069 29412
rect 26003 28660 26069 28661
rect 26003 28596 26004 28660
rect 26068 28596 26069 28660
rect 26003 28595 26069 28596
rect 26006 28389 26066 28595
rect 26190 28389 26250 31995
rect 26558 30698 26618 34171
rect 30235 33420 30301 33421
rect 30235 33356 30236 33420
rect 30300 33356 30301 33420
rect 30235 33355 30301 33356
rect 30051 32876 30117 32877
rect 30051 32812 30052 32876
rect 30116 32812 30117 32876
rect 30051 32811 30117 32812
rect 27831 32128 28151 32688
rect 27831 32064 27839 32128
rect 27903 32064 27919 32128
rect 27983 32064 27999 32128
rect 28063 32064 28079 32128
rect 28143 32064 28151 32128
rect 27291 31652 27357 31653
rect 27291 31588 27292 31652
rect 27356 31588 27357 31652
rect 27291 31587 27357 31588
rect 27107 30700 27173 30701
rect 26558 30638 26986 30698
rect 26371 30020 26437 30021
rect 26371 29956 26372 30020
rect 26436 29956 26437 30020
rect 26371 29955 26437 29956
rect 26003 28388 26069 28389
rect 26003 28324 26004 28388
rect 26068 28324 26069 28388
rect 26003 28323 26069 28324
rect 26187 28388 26253 28389
rect 26187 28324 26188 28388
rect 26252 28324 26253 28388
rect 26187 28323 26253 28324
rect 25819 28252 25885 28253
rect 25819 28188 25820 28252
rect 25884 28188 25885 28252
rect 25819 28187 25885 28188
rect 26003 28252 26069 28253
rect 26003 28188 26004 28252
rect 26068 28188 26069 28252
rect 26374 28250 26434 29955
rect 26558 29205 26618 30638
rect 26926 30565 26986 30638
rect 27107 30636 27108 30700
rect 27172 30636 27173 30700
rect 27107 30635 27173 30636
rect 26739 30564 26805 30565
rect 26739 30500 26740 30564
rect 26804 30500 26805 30564
rect 26739 30499 26805 30500
rect 26923 30564 26989 30565
rect 26923 30500 26924 30564
rect 26988 30500 26989 30564
rect 26923 30499 26989 30500
rect 26555 29204 26621 29205
rect 26555 29140 26556 29204
rect 26620 29140 26621 29204
rect 26555 29139 26621 29140
rect 26003 28187 26069 28188
rect 26190 28190 26434 28250
rect 25635 28116 25701 28117
rect 25635 28052 25636 28116
rect 25700 28052 25701 28116
rect 25635 28051 25701 28052
rect 25451 26348 25517 26349
rect 25451 26284 25452 26348
rect 25516 26284 25517 26348
rect 25451 26283 25517 26284
rect 25267 25532 25333 25533
rect 25267 25468 25268 25532
rect 25332 25468 25333 25532
rect 25267 25467 25333 25468
rect 25267 25260 25333 25261
rect 25267 25196 25268 25260
rect 25332 25196 25333 25260
rect 25267 25195 25333 25196
rect 25083 24988 25149 24989
rect 25083 24924 25084 24988
rect 25148 24924 25149 24988
rect 25083 24923 25149 24924
rect 25083 22404 25149 22405
rect 25083 22340 25084 22404
rect 25148 22402 25149 22404
rect 25270 22402 25330 25195
rect 25148 22342 25330 22402
rect 25148 22340 25149 22342
rect 25083 22339 25149 22340
rect 25638 22133 25698 28051
rect 25822 24445 25882 28187
rect 26006 25941 26066 28187
rect 26003 25940 26069 25941
rect 26003 25876 26004 25940
rect 26068 25876 26069 25940
rect 26003 25875 26069 25876
rect 25819 24444 25885 24445
rect 25819 24380 25820 24444
rect 25884 24380 25885 24444
rect 25819 24379 25885 24380
rect 26190 22133 26250 28190
rect 26371 27844 26437 27845
rect 26371 27780 26372 27844
rect 26436 27780 26437 27844
rect 26371 27779 26437 27780
rect 26374 24853 26434 27779
rect 26558 25125 26618 29139
rect 26742 27301 26802 30499
rect 26923 29476 26989 29477
rect 26923 29412 26924 29476
rect 26988 29412 26989 29476
rect 26923 29411 26989 29412
rect 26926 29205 26986 29411
rect 26923 29204 26989 29205
rect 26923 29140 26924 29204
rect 26988 29140 26989 29204
rect 26923 29139 26989 29140
rect 26923 29068 26989 29069
rect 26923 29004 26924 29068
rect 26988 29004 26989 29068
rect 26923 29003 26989 29004
rect 26926 27845 26986 29003
rect 26923 27844 26989 27845
rect 26923 27780 26924 27844
rect 26988 27780 26989 27844
rect 26923 27779 26989 27780
rect 26923 27572 26989 27573
rect 26923 27508 26924 27572
rect 26988 27508 26989 27572
rect 26923 27507 26989 27508
rect 26739 27300 26805 27301
rect 26739 27236 26740 27300
rect 26804 27236 26805 27300
rect 26739 27235 26805 27236
rect 26742 26893 26802 27235
rect 26739 26892 26805 26893
rect 26739 26828 26740 26892
rect 26804 26828 26805 26892
rect 26739 26827 26805 26828
rect 26739 26620 26805 26621
rect 26739 26556 26740 26620
rect 26804 26556 26805 26620
rect 26739 26555 26805 26556
rect 26555 25124 26621 25125
rect 26555 25060 26556 25124
rect 26620 25060 26621 25124
rect 26555 25059 26621 25060
rect 26742 24853 26802 26555
rect 26371 24852 26437 24853
rect 26371 24788 26372 24852
rect 26436 24788 26437 24852
rect 26371 24787 26437 24788
rect 26739 24852 26805 24853
rect 26739 24788 26740 24852
rect 26804 24788 26805 24852
rect 26739 24787 26805 24788
rect 26739 23764 26805 23765
rect 26739 23700 26740 23764
rect 26804 23762 26805 23764
rect 26926 23762 26986 27507
rect 27110 24581 27170 30635
rect 27294 30021 27354 31587
rect 27831 31040 28151 32064
rect 28763 31652 28829 31653
rect 28763 31588 28764 31652
rect 28828 31588 28829 31652
rect 28763 31587 28829 31588
rect 27831 30976 27839 31040
rect 27903 30976 27919 31040
rect 27983 30976 27999 31040
rect 28063 30976 28079 31040
rect 28143 30976 28151 31040
rect 27475 30836 27541 30837
rect 27475 30772 27476 30836
rect 27540 30772 27541 30836
rect 27475 30771 27541 30772
rect 27291 30020 27357 30021
rect 27291 29956 27292 30020
rect 27356 29956 27357 30020
rect 27291 29955 27357 29956
rect 27291 29884 27357 29885
rect 27291 29820 27292 29884
rect 27356 29820 27357 29884
rect 27291 29819 27357 29820
rect 27294 29069 27354 29819
rect 27291 29068 27357 29069
rect 27291 29004 27292 29068
rect 27356 29004 27357 29068
rect 27291 29003 27357 29004
rect 27291 26348 27357 26349
rect 27291 26284 27292 26348
rect 27356 26284 27357 26348
rect 27291 26283 27357 26284
rect 27107 24580 27173 24581
rect 27107 24516 27108 24580
rect 27172 24516 27173 24580
rect 27107 24515 27173 24516
rect 26804 23702 26986 23762
rect 26804 23700 26805 23702
rect 26739 23699 26805 23700
rect 26739 23492 26805 23493
rect 26739 23428 26740 23492
rect 26804 23428 26805 23492
rect 26739 23427 26805 23428
rect 26371 22540 26437 22541
rect 26371 22476 26372 22540
rect 26436 22476 26437 22540
rect 26371 22475 26437 22476
rect 26374 22133 26434 22475
rect 25635 22132 25701 22133
rect 25635 22068 25636 22132
rect 25700 22068 25701 22132
rect 25635 22067 25701 22068
rect 26187 22132 26253 22133
rect 26187 22068 26188 22132
rect 26252 22068 26253 22132
rect 26187 22067 26253 22068
rect 26371 22132 26437 22133
rect 26371 22068 26372 22132
rect 26436 22068 26437 22132
rect 26371 22067 26437 22068
rect 26555 21860 26621 21861
rect 26555 21796 26556 21860
rect 26620 21796 26621 21860
rect 26555 21795 26621 21796
rect 26558 21317 26618 21795
rect 26555 21316 26621 21317
rect 26555 21252 26556 21316
rect 26620 21252 26621 21316
rect 26555 21251 26621 21252
rect 26742 21178 26802 23427
rect 27110 23357 27170 24515
rect 27294 23629 27354 26283
rect 27478 24037 27538 30771
rect 27659 30428 27725 30429
rect 27659 30364 27660 30428
rect 27724 30364 27725 30428
rect 27659 30363 27725 30364
rect 27662 27845 27722 30363
rect 27831 29952 28151 30976
rect 28395 30972 28461 30973
rect 28395 30908 28396 30972
rect 28460 30908 28461 30972
rect 28395 30907 28461 30908
rect 28257 30020 28323 30021
rect 28257 30018 28258 30020
rect 27831 29888 27839 29952
rect 27903 29888 27919 29952
rect 27983 29888 27999 29952
rect 28063 29888 28079 29952
rect 28143 29888 28151 29952
rect 27831 28864 28151 29888
rect 28214 29956 28258 30018
rect 28322 29956 28323 30020
rect 28214 29955 28323 29956
rect 28214 29341 28274 29955
rect 28211 29340 28277 29341
rect 28211 29276 28212 29340
rect 28276 29276 28277 29340
rect 28211 29275 28277 29276
rect 27831 28800 27839 28864
rect 27903 28800 27919 28864
rect 27983 28800 27999 28864
rect 28063 28800 28079 28864
rect 28143 28800 28151 28864
rect 27659 27844 27725 27845
rect 27659 27780 27660 27844
rect 27724 27780 27725 27844
rect 27659 27779 27725 27780
rect 27831 27776 28151 28800
rect 28211 28388 28277 28389
rect 28211 28324 28212 28388
rect 28276 28324 28277 28388
rect 28211 28323 28277 28324
rect 27831 27712 27839 27776
rect 27903 27712 27919 27776
rect 27983 27712 27999 27776
rect 28063 27712 28079 27776
rect 28143 27712 28151 27776
rect 27659 27708 27725 27709
rect 27659 27644 27660 27708
rect 27724 27644 27725 27708
rect 27659 27643 27725 27644
rect 27662 27165 27722 27643
rect 27659 27164 27725 27165
rect 27659 27100 27660 27164
rect 27724 27100 27725 27164
rect 27659 27099 27725 27100
rect 27831 26688 28151 27712
rect 28214 27709 28274 28323
rect 28214 27708 28323 27709
rect 28214 27646 28258 27708
rect 28257 27644 28258 27646
rect 28322 27644 28323 27708
rect 28257 27643 28323 27644
rect 27831 26624 27839 26688
rect 27903 26624 27919 26688
rect 27983 26624 27999 26688
rect 28063 26624 28079 26688
rect 28143 26624 28151 26688
rect 27659 26620 27725 26621
rect 27659 26556 27660 26620
rect 27724 26556 27725 26620
rect 27659 26555 27725 26556
rect 27662 25805 27722 26555
rect 27659 25804 27725 25805
rect 27659 25740 27660 25804
rect 27724 25740 27725 25804
rect 27659 25739 27725 25740
rect 27659 25668 27725 25669
rect 27659 25604 27660 25668
rect 27724 25604 27725 25668
rect 27659 25603 27725 25604
rect 27475 24036 27541 24037
rect 27475 23972 27476 24036
rect 27540 23972 27541 24036
rect 27475 23971 27541 23972
rect 27291 23628 27357 23629
rect 27291 23564 27292 23628
rect 27356 23564 27357 23628
rect 27291 23563 27357 23564
rect 27107 23356 27173 23357
rect 27107 23292 27108 23356
rect 27172 23292 27173 23356
rect 27107 23291 27173 23292
rect 26558 21118 26802 21178
rect 25083 20772 25149 20773
rect 25083 20708 25084 20772
rect 25148 20708 25149 20772
rect 25083 20707 25149 20708
rect 24899 19820 24965 19821
rect 24899 19756 24900 19820
rect 24964 19756 24965 19820
rect 24899 19755 24965 19756
rect 24899 19004 24965 19005
rect 24899 18940 24900 19004
rect 24964 18940 24965 19004
rect 24899 18939 24965 18940
rect 24715 18052 24781 18053
rect 24715 17988 24716 18052
rect 24780 17988 24781 18052
rect 24715 17987 24781 17988
rect 24531 15468 24597 15469
rect 24531 15404 24532 15468
rect 24596 15404 24597 15468
rect 24531 15403 24597 15404
rect 23990 15200 23998 15264
rect 24062 15200 24078 15264
rect 24142 15200 24158 15264
rect 24222 15200 24238 15264
rect 24302 15200 24310 15264
rect 23990 14176 24310 15200
rect 23990 14112 23998 14176
rect 24062 14112 24078 14176
rect 24142 14112 24158 14176
rect 24222 14112 24238 14176
rect 24302 14112 24310 14176
rect 23990 13088 24310 14112
rect 23990 13024 23998 13088
rect 24062 13024 24078 13088
rect 24142 13024 24158 13088
rect 24222 13024 24238 13088
rect 24302 13024 24310 13088
rect 23795 12884 23861 12885
rect 23795 12820 23796 12884
rect 23860 12820 23861 12884
rect 23795 12819 23861 12820
rect 23990 12000 24310 13024
rect 23990 11936 23998 12000
rect 24062 11936 24078 12000
rect 24142 11936 24158 12000
rect 24222 11936 24238 12000
rect 24302 11936 24310 12000
rect 23990 10912 24310 11936
rect 24718 11933 24778 17987
rect 24902 17781 24962 18939
rect 24899 17780 24965 17781
rect 24899 17716 24900 17780
rect 24964 17716 24965 17780
rect 24899 17715 24965 17716
rect 24899 15332 24965 15333
rect 24899 15268 24900 15332
rect 24964 15268 24965 15332
rect 24899 15267 24965 15268
rect 24902 12205 24962 15267
rect 25086 12341 25146 20707
rect 26003 20092 26069 20093
rect 26003 20028 26004 20092
rect 26068 20028 26069 20092
rect 26003 20027 26069 20028
rect 26371 20092 26437 20093
rect 26371 20028 26372 20092
rect 26436 20028 26437 20092
rect 26371 20027 26437 20028
rect 25635 19820 25701 19821
rect 25635 19756 25636 19820
rect 25700 19756 25701 19820
rect 25635 19755 25701 19756
rect 25451 18188 25517 18189
rect 25451 18124 25452 18188
rect 25516 18124 25517 18188
rect 25451 18123 25517 18124
rect 25267 14516 25333 14517
rect 25267 14452 25268 14516
rect 25332 14452 25333 14516
rect 25267 14451 25333 14452
rect 25270 13837 25330 14451
rect 25267 13836 25333 13837
rect 25267 13772 25268 13836
rect 25332 13772 25333 13836
rect 25267 13771 25333 13772
rect 25454 13157 25514 18123
rect 25638 15197 25698 19755
rect 26006 18461 26066 20027
rect 26187 19140 26253 19141
rect 26187 19076 26188 19140
rect 26252 19076 26253 19140
rect 26187 19075 26253 19076
rect 26003 18460 26069 18461
rect 26003 18396 26004 18460
rect 26068 18396 26069 18460
rect 26003 18395 26069 18396
rect 26190 18050 26250 19075
rect 26374 18189 26434 20027
rect 26558 19141 26618 21118
rect 26923 21044 26989 21045
rect 26923 20980 26924 21044
rect 26988 20980 26989 21044
rect 26923 20979 26989 20980
rect 26739 20636 26805 20637
rect 26739 20572 26740 20636
rect 26804 20572 26805 20636
rect 26739 20571 26805 20572
rect 26555 19140 26621 19141
rect 26555 19076 26556 19140
rect 26620 19076 26621 19140
rect 26555 19075 26621 19076
rect 26371 18188 26437 18189
rect 26371 18124 26372 18188
rect 26436 18124 26437 18188
rect 26371 18123 26437 18124
rect 26190 17990 26618 18050
rect 26187 17780 26253 17781
rect 26187 17716 26188 17780
rect 26252 17716 26253 17780
rect 26187 17715 26253 17716
rect 26003 16964 26069 16965
rect 26003 16900 26004 16964
rect 26068 16900 26069 16964
rect 26003 16899 26069 16900
rect 25819 16556 25885 16557
rect 25819 16492 25820 16556
rect 25884 16492 25885 16556
rect 25819 16491 25885 16492
rect 25822 15333 25882 16491
rect 25819 15332 25885 15333
rect 25819 15268 25820 15332
rect 25884 15268 25885 15332
rect 25819 15267 25885 15268
rect 25635 15196 25701 15197
rect 25635 15132 25636 15196
rect 25700 15132 25701 15196
rect 25635 15131 25701 15132
rect 26006 13973 26066 16899
rect 26003 13972 26069 13973
rect 26003 13908 26004 13972
rect 26068 13908 26069 13972
rect 26003 13907 26069 13908
rect 25819 13836 25885 13837
rect 25819 13772 25820 13836
rect 25884 13772 25885 13836
rect 25819 13771 25885 13772
rect 25451 13156 25517 13157
rect 25451 13092 25452 13156
rect 25516 13092 25517 13156
rect 25451 13091 25517 13092
rect 25083 12340 25149 12341
rect 25083 12276 25084 12340
rect 25148 12276 25149 12340
rect 25083 12275 25149 12276
rect 24899 12204 24965 12205
rect 24899 12140 24900 12204
rect 24964 12140 24965 12204
rect 24899 12139 24965 12140
rect 24715 11932 24781 11933
rect 24715 11868 24716 11932
rect 24780 11868 24781 11932
rect 24715 11867 24781 11868
rect 23990 10848 23998 10912
rect 24062 10848 24078 10912
rect 24142 10848 24158 10912
rect 24222 10848 24238 10912
rect 24302 10848 24310 10912
rect 23611 10708 23677 10709
rect 23611 10644 23612 10708
rect 23676 10644 23677 10708
rect 23611 10643 23677 10644
rect 23990 9824 24310 10848
rect 23990 9760 23998 9824
rect 24062 9760 24078 9824
rect 24142 9760 24158 9824
rect 24222 9760 24238 9824
rect 24302 9760 24310 9824
rect 23990 8736 24310 9760
rect 25822 9621 25882 13771
rect 26190 11389 26250 17715
rect 26371 17236 26437 17237
rect 26371 17172 26372 17236
rect 26436 17172 26437 17236
rect 26371 17171 26437 17172
rect 26374 13021 26434 17171
rect 26558 13837 26618 17990
rect 26742 15469 26802 20571
rect 26926 19821 26986 20979
rect 27110 20365 27170 23291
rect 27478 22541 27538 23971
rect 27662 23357 27722 25603
rect 27831 25600 28151 26624
rect 28398 26485 28458 30907
rect 28579 29748 28645 29749
rect 28579 29684 28580 29748
rect 28644 29684 28645 29748
rect 28579 29683 28645 29684
rect 28582 28389 28642 29683
rect 28766 28933 28826 31587
rect 29315 31108 29381 31109
rect 29315 31044 29316 31108
rect 29380 31044 29381 31108
rect 29315 31043 29381 31044
rect 28947 29612 29013 29613
rect 28947 29548 28948 29612
rect 29012 29548 29013 29612
rect 28947 29547 29013 29548
rect 28763 28932 28829 28933
rect 28763 28868 28764 28932
rect 28828 28868 28829 28932
rect 28763 28867 28829 28868
rect 28579 28388 28645 28389
rect 28579 28324 28580 28388
rect 28644 28324 28645 28388
rect 28579 28323 28645 28324
rect 28579 27980 28645 27981
rect 28579 27916 28580 27980
rect 28644 27916 28645 27980
rect 28579 27915 28645 27916
rect 28395 26484 28461 26485
rect 28395 26420 28396 26484
rect 28460 26420 28461 26484
rect 28395 26419 28461 26420
rect 28211 26348 28277 26349
rect 28211 26284 28212 26348
rect 28276 26284 28277 26348
rect 28211 26283 28277 26284
rect 27831 25536 27839 25600
rect 27903 25536 27919 25600
rect 27983 25536 27999 25600
rect 28063 25536 28079 25600
rect 28143 25536 28151 25600
rect 27831 24512 28151 25536
rect 27831 24448 27839 24512
rect 27903 24448 27919 24512
rect 27983 24448 27999 24512
rect 28063 24448 28079 24512
rect 28143 24448 28151 24512
rect 27831 23424 28151 24448
rect 27831 23360 27839 23424
rect 27903 23360 27919 23424
rect 27983 23360 27999 23424
rect 28063 23360 28079 23424
rect 28143 23360 28151 23424
rect 27659 23356 27725 23357
rect 27659 23292 27660 23356
rect 27724 23292 27725 23356
rect 27659 23291 27725 23292
rect 27475 22540 27541 22541
rect 27475 22476 27476 22540
rect 27540 22476 27541 22540
rect 27475 22475 27541 22476
rect 27659 22540 27725 22541
rect 27659 22476 27660 22540
rect 27724 22476 27725 22540
rect 27659 22475 27725 22476
rect 27475 21044 27541 21045
rect 27475 20980 27476 21044
rect 27540 20980 27541 21044
rect 27475 20979 27541 20980
rect 27291 20636 27357 20637
rect 27291 20572 27292 20636
rect 27356 20572 27357 20636
rect 27291 20571 27357 20572
rect 27294 20365 27354 20571
rect 27107 20364 27173 20365
rect 27107 20300 27108 20364
rect 27172 20300 27173 20364
rect 27107 20299 27173 20300
rect 27291 20364 27357 20365
rect 27291 20300 27292 20364
rect 27356 20300 27357 20364
rect 27291 20299 27357 20300
rect 26923 19820 26989 19821
rect 26923 19756 26924 19820
rect 26988 19756 26989 19820
rect 26923 19755 26989 19756
rect 27107 19820 27173 19821
rect 27107 19756 27108 19820
rect 27172 19756 27173 19820
rect 27107 19755 27173 19756
rect 26923 19140 26989 19141
rect 26923 19076 26924 19140
rect 26988 19076 26989 19140
rect 26923 19075 26989 19076
rect 26926 16965 26986 19075
rect 27110 17509 27170 19755
rect 27291 18052 27357 18053
rect 27291 17988 27292 18052
rect 27356 17988 27357 18052
rect 27291 17987 27357 17988
rect 27107 17508 27173 17509
rect 27107 17444 27108 17508
rect 27172 17444 27173 17508
rect 27107 17443 27173 17444
rect 26923 16964 26989 16965
rect 26923 16900 26924 16964
rect 26988 16900 26989 16964
rect 26923 16899 26989 16900
rect 26923 16828 26989 16829
rect 26923 16764 26924 16828
rect 26988 16764 26989 16828
rect 26923 16763 26989 16764
rect 26739 15468 26805 15469
rect 26739 15404 26740 15468
rect 26804 15404 26805 15468
rect 26739 15403 26805 15404
rect 26555 13836 26621 13837
rect 26555 13772 26556 13836
rect 26620 13772 26621 13836
rect 26555 13771 26621 13772
rect 26371 13020 26437 13021
rect 26371 12956 26372 13020
rect 26436 12956 26437 13020
rect 26371 12955 26437 12956
rect 26187 11388 26253 11389
rect 26187 11324 26188 11388
rect 26252 11324 26253 11388
rect 26187 11323 26253 11324
rect 25819 9620 25885 9621
rect 25819 9556 25820 9620
rect 25884 9556 25885 9620
rect 25819 9555 25885 9556
rect 26742 9349 26802 15403
rect 26926 11933 26986 16763
rect 26923 11932 26989 11933
rect 26923 11868 26924 11932
rect 26988 11868 26989 11932
rect 26923 11867 26989 11868
rect 27110 10981 27170 17443
rect 27294 12885 27354 17987
rect 27478 17781 27538 20979
rect 27662 20229 27722 22475
rect 27831 22336 28151 23360
rect 27831 22272 27839 22336
rect 27903 22272 27919 22336
rect 27983 22272 27999 22336
rect 28063 22272 28079 22336
rect 28143 22272 28151 22336
rect 27831 21248 28151 22272
rect 27831 21184 27839 21248
rect 27903 21184 27919 21248
rect 27983 21184 27999 21248
rect 28063 21184 28079 21248
rect 28143 21184 28151 21248
rect 27659 20228 27725 20229
rect 27659 20164 27660 20228
rect 27724 20164 27725 20228
rect 27659 20163 27725 20164
rect 27831 20160 28151 21184
rect 27831 20096 27839 20160
rect 27903 20096 27919 20160
rect 27983 20096 27999 20160
rect 28063 20096 28079 20160
rect 28143 20096 28151 20160
rect 27831 19072 28151 20096
rect 28214 19413 28274 26283
rect 28395 26076 28461 26077
rect 28395 26012 28396 26076
rect 28460 26012 28461 26076
rect 28395 26011 28461 26012
rect 28398 23493 28458 26011
rect 28395 23492 28461 23493
rect 28395 23428 28396 23492
rect 28460 23428 28461 23492
rect 28395 23427 28461 23428
rect 28395 23356 28461 23357
rect 28395 23292 28396 23356
rect 28460 23292 28461 23356
rect 28395 23291 28461 23292
rect 28398 22269 28458 23291
rect 28395 22268 28461 22269
rect 28395 22204 28396 22268
rect 28460 22204 28461 22268
rect 28395 22203 28461 22204
rect 28395 21180 28461 21181
rect 28395 21116 28396 21180
rect 28460 21116 28461 21180
rect 28395 21115 28461 21116
rect 28398 20365 28458 21115
rect 28395 20364 28461 20365
rect 28395 20300 28396 20364
rect 28460 20300 28461 20364
rect 28395 20299 28461 20300
rect 28582 20093 28642 27915
rect 28766 26621 28826 28867
rect 28763 26620 28829 26621
rect 28763 26556 28764 26620
rect 28828 26556 28829 26620
rect 28763 26555 28829 26556
rect 28763 26348 28829 26349
rect 28763 26284 28764 26348
rect 28828 26284 28829 26348
rect 28763 26283 28829 26284
rect 28766 23357 28826 26283
rect 28763 23356 28829 23357
rect 28763 23292 28764 23356
rect 28828 23292 28829 23356
rect 28763 23291 28829 23292
rect 28579 20092 28645 20093
rect 28579 20028 28580 20092
rect 28644 20028 28645 20092
rect 28579 20027 28645 20028
rect 28211 19412 28277 19413
rect 28211 19348 28212 19412
rect 28276 19348 28277 19412
rect 28211 19347 28277 19348
rect 28395 19140 28461 19141
rect 28395 19138 28396 19140
rect 27831 19008 27839 19072
rect 27903 19008 27919 19072
rect 27983 19008 27999 19072
rect 28063 19008 28079 19072
rect 28143 19008 28151 19072
rect 27831 17984 28151 19008
rect 27831 17920 27839 17984
rect 27903 17920 27919 17984
rect 27983 17920 27999 17984
rect 28063 17920 28079 17984
rect 28143 17920 28151 17984
rect 27475 17780 27541 17781
rect 27475 17716 27476 17780
rect 27540 17716 27541 17780
rect 27475 17715 27541 17716
rect 27478 17506 27538 17715
rect 27659 17508 27725 17509
rect 27659 17506 27660 17508
rect 27478 17446 27660 17506
rect 27659 17444 27660 17446
rect 27724 17444 27725 17508
rect 27659 17443 27725 17444
rect 27662 13157 27722 17443
rect 27831 16896 28151 17920
rect 27831 16832 27839 16896
rect 27903 16832 27919 16896
rect 27983 16832 27999 16896
rect 28063 16832 28079 16896
rect 28143 16832 28151 16896
rect 27831 15808 28151 16832
rect 27831 15744 27839 15808
rect 27903 15744 27919 15808
rect 27983 15744 27999 15808
rect 28063 15744 28079 15808
rect 28143 15744 28151 15808
rect 27831 14720 28151 15744
rect 27831 14656 27839 14720
rect 27903 14656 27919 14720
rect 27983 14656 27999 14720
rect 28063 14656 28079 14720
rect 28143 14656 28151 14720
rect 27831 13632 28151 14656
rect 28214 19078 28396 19138
rect 28214 13837 28274 19078
rect 28395 19076 28396 19078
rect 28460 19076 28461 19140
rect 28395 19075 28461 19076
rect 28395 18188 28461 18189
rect 28395 18124 28396 18188
rect 28460 18124 28461 18188
rect 28395 18123 28461 18124
rect 28398 16829 28458 18123
rect 28766 17781 28826 23291
rect 28950 22269 29010 29547
rect 29131 29476 29197 29477
rect 29131 29412 29132 29476
rect 29196 29412 29197 29476
rect 29131 29411 29197 29412
rect 29134 25669 29194 29411
rect 29318 28661 29378 31043
rect 29499 29884 29565 29885
rect 29499 29820 29500 29884
rect 29564 29820 29565 29884
rect 29499 29819 29565 29820
rect 29502 28661 29562 29819
rect 29683 29340 29749 29341
rect 29683 29276 29684 29340
rect 29748 29276 29749 29340
rect 29683 29275 29749 29276
rect 29315 28660 29381 28661
rect 29315 28596 29316 28660
rect 29380 28596 29381 28660
rect 29315 28595 29381 28596
rect 29499 28660 29565 28661
rect 29499 28596 29500 28660
rect 29564 28596 29565 28660
rect 29499 28595 29565 28596
rect 29499 28388 29565 28389
rect 29499 28324 29500 28388
rect 29564 28324 29565 28388
rect 29499 28323 29565 28324
rect 29315 28252 29381 28253
rect 29315 28188 29316 28252
rect 29380 28188 29381 28252
rect 29315 28187 29381 28188
rect 29131 25668 29197 25669
rect 29131 25604 29132 25668
rect 29196 25604 29197 25668
rect 29131 25603 29197 25604
rect 29131 25532 29197 25533
rect 29131 25468 29132 25532
rect 29196 25468 29197 25532
rect 29131 25467 29197 25468
rect 29134 24853 29194 25467
rect 29131 24852 29197 24853
rect 29131 24788 29132 24852
rect 29196 24788 29197 24852
rect 29131 24787 29197 24788
rect 28947 22268 29013 22269
rect 28947 22204 28948 22268
rect 29012 22204 29013 22268
rect 28947 22203 29013 22204
rect 29131 21860 29197 21861
rect 29131 21796 29132 21860
rect 29196 21796 29197 21860
rect 29131 21795 29197 21796
rect 28947 20092 29013 20093
rect 28947 20028 28948 20092
rect 29012 20028 29013 20092
rect 28947 20027 29013 20028
rect 28763 17780 28829 17781
rect 28763 17716 28764 17780
rect 28828 17716 28829 17780
rect 28763 17715 28829 17716
rect 28579 17508 28645 17509
rect 28579 17444 28580 17508
rect 28644 17444 28645 17508
rect 28579 17443 28645 17444
rect 28395 16828 28461 16829
rect 28395 16764 28396 16828
rect 28460 16764 28461 16828
rect 28395 16763 28461 16764
rect 28395 16692 28461 16693
rect 28395 16628 28396 16692
rect 28460 16628 28461 16692
rect 28395 16627 28461 16628
rect 28211 13836 28277 13837
rect 28211 13772 28212 13836
rect 28276 13772 28277 13836
rect 28211 13771 28277 13772
rect 27831 13568 27839 13632
rect 27903 13568 27919 13632
rect 27983 13568 27999 13632
rect 28063 13568 28079 13632
rect 28143 13568 28151 13632
rect 27659 13156 27725 13157
rect 27659 13092 27660 13156
rect 27724 13092 27725 13156
rect 27659 13091 27725 13092
rect 27291 12884 27357 12885
rect 27291 12820 27292 12884
rect 27356 12820 27357 12884
rect 27291 12819 27357 12820
rect 27831 12544 28151 13568
rect 28398 12885 28458 16627
rect 28395 12884 28461 12885
rect 28395 12820 28396 12884
rect 28460 12820 28461 12884
rect 28395 12819 28461 12820
rect 27831 12480 27839 12544
rect 27903 12480 27919 12544
rect 27983 12480 27999 12544
rect 28063 12480 28079 12544
rect 28143 12480 28151 12544
rect 27831 11456 28151 12480
rect 27831 11392 27839 11456
rect 27903 11392 27919 11456
rect 27983 11392 27999 11456
rect 28063 11392 28079 11456
rect 28143 11392 28151 11456
rect 27107 10980 27173 10981
rect 27107 10916 27108 10980
rect 27172 10916 27173 10980
rect 27107 10915 27173 10916
rect 27110 9757 27170 10915
rect 27831 10368 28151 11392
rect 28582 11117 28642 17443
rect 28950 16590 29010 20027
rect 29134 18325 29194 21795
rect 29318 19413 29378 28187
rect 29502 27709 29562 28323
rect 29499 27708 29565 27709
rect 29499 27644 29500 27708
rect 29564 27644 29565 27708
rect 29499 27643 29565 27644
rect 29686 27434 29746 29275
rect 29867 27844 29933 27845
rect 29867 27780 29868 27844
rect 29932 27780 29933 27844
rect 29867 27779 29933 27780
rect 29502 27374 29746 27434
rect 29502 26621 29562 27374
rect 29683 27300 29749 27301
rect 29683 27236 29684 27300
rect 29748 27236 29749 27300
rect 29683 27235 29749 27236
rect 29686 26893 29746 27235
rect 29683 26892 29749 26893
rect 29683 26828 29684 26892
rect 29748 26828 29749 26892
rect 29683 26827 29749 26828
rect 29499 26620 29565 26621
rect 29499 26556 29500 26620
rect 29564 26556 29565 26620
rect 29499 26555 29565 26556
rect 29499 26484 29565 26485
rect 29499 26420 29500 26484
rect 29564 26420 29565 26484
rect 29499 26419 29565 26420
rect 29502 19549 29562 26419
rect 29683 26348 29749 26349
rect 29683 26284 29684 26348
rect 29748 26284 29749 26348
rect 29683 26283 29749 26284
rect 29686 20909 29746 26283
rect 29870 25941 29930 27779
rect 30054 27301 30114 32811
rect 30051 27300 30117 27301
rect 30051 27236 30052 27300
rect 30116 27236 30117 27300
rect 30051 27235 30117 27236
rect 30238 27165 30298 33355
rect 31672 32672 31992 32688
rect 31672 32608 31680 32672
rect 31744 32608 31760 32672
rect 31824 32608 31840 32672
rect 31904 32608 31920 32672
rect 31984 32608 31992 32672
rect 31672 31584 31992 32608
rect 31672 31520 31680 31584
rect 31744 31520 31760 31584
rect 31824 31520 31840 31584
rect 31904 31520 31920 31584
rect 31984 31520 31992 31584
rect 30787 31244 30853 31245
rect 30787 31180 30788 31244
rect 30852 31180 30853 31244
rect 30787 31179 30853 31180
rect 30419 30836 30485 30837
rect 30419 30772 30420 30836
rect 30484 30772 30485 30836
rect 30419 30771 30485 30772
rect 30235 27164 30301 27165
rect 30235 27100 30236 27164
rect 30300 27100 30301 27164
rect 30235 27099 30301 27100
rect 30051 26620 30117 26621
rect 30051 26556 30052 26620
rect 30116 26556 30117 26620
rect 30051 26555 30117 26556
rect 29867 25940 29933 25941
rect 29867 25876 29868 25940
rect 29932 25876 29933 25940
rect 29867 25875 29933 25876
rect 29870 24989 29930 25875
rect 29867 24988 29933 24989
rect 29867 24924 29868 24988
rect 29932 24924 29933 24988
rect 29867 24923 29933 24924
rect 29867 24444 29933 24445
rect 29867 24380 29868 24444
rect 29932 24380 29933 24444
rect 29867 24379 29933 24380
rect 29870 22946 29930 24379
rect 30054 24309 30114 26555
rect 30051 24308 30117 24309
rect 30051 24244 30052 24308
rect 30116 24244 30117 24308
rect 30051 24243 30117 24244
rect 30238 23357 30298 27099
rect 30422 27029 30482 30771
rect 30603 30428 30669 30429
rect 30603 30364 30604 30428
rect 30668 30364 30669 30428
rect 30603 30363 30669 30364
rect 30419 27028 30485 27029
rect 30419 26964 30420 27028
rect 30484 26964 30485 27028
rect 30419 26963 30485 26964
rect 30606 26621 30666 30363
rect 30603 26620 30669 26621
rect 30603 26556 30604 26620
rect 30668 26556 30669 26620
rect 30603 26555 30669 26556
rect 30419 26484 30485 26485
rect 30419 26420 30420 26484
rect 30484 26420 30485 26484
rect 30419 26419 30485 26420
rect 30235 23356 30301 23357
rect 30235 23292 30236 23356
rect 30300 23292 30301 23356
rect 30235 23291 30301 23292
rect 29870 22886 30114 22946
rect 29867 22812 29933 22813
rect 29867 22748 29868 22812
rect 29932 22748 29933 22812
rect 29867 22747 29933 22748
rect 29683 20908 29749 20909
rect 29683 20844 29684 20908
rect 29748 20844 29749 20908
rect 29683 20843 29749 20844
rect 29683 20772 29749 20773
rect 29683 20708 29684 20772
rect 29748 20770 29749 20772
rect 29870 20770 29930 22747
rect 30054 21045 30114 22886
rect 30235 22812 30301 22813
rect 30235 22748 30236 22812
rect 30300 22748 30301 22812
rect 30235 22747 30301 22748
rect 30051 21044 30117 21045
rect 30051 20980 30052 21044
rect 30116 20980 30117 21044
rect 30051 20979 30117 20980
rect 29748 20710 29930 20770
rect 29748 20708 29749 20710
rect 29683 20707 29749 20708
rect 29499 19548 29565 19549
rect 29499 19484 29500 19548
rect 29564 19484 29565 19548
rect 29499 19483 29565 19484
rect 29315 19412 29381 19413
rect 29315 19348 29316 19412
rect 29380 19348 29381 19412
rect 29315 19347 29381 19348
rect 29315 19140 29381 19141
rect 29315 19076 29316 19140
rect 29380 19076 29381 19140
rect 29315 19075 29381 19076
rect 29131 18324 29197 18325
rect 29131 18260 29132 18324
rect 29196 18260 29197 18324
rect 29131 18259 29197 18260
rect 29131 18188 29197 18189
rect 29131 18124 29132 18188
rect 29196 18124 29197 18188
rect 29131 18123 29197 18124
rect 29134 16965 29194 18123
rect 29131 16964 29197 16965
rect 29131 16900 29132 16964
rect 29196 16900 29197 16964
rect 29131 16899 29197 16900
rect 29131 16828 29197 16829
rect 29131 16764 29132 16828
rect 29196 16764 29197 16828
rect 29131 16763 29197 16764
rect 28766 16557 29010 16590
rect 28766 16556 29013 16557
rect 28766 16530 28948 16556
rect 28579 11116 28645 11117
rect 28579 11052 28580 11116
rect 28644 11052 28645 11116
rect 28579 11051 28645 11052
rect 27831 10304 27839 10368
rect 27903 10304 27919 10368
rect 27983 10304 27999 10368
rect 28063 10304 28079 10368
rect 28143 10304 28151 10368
rect 27107 9756 27173 9757
rect 27107 9692 27108 9756
rect 27172 9692 27173 9756
rect 27107 9691 27173 9692
rect 26739 9348 26805 9349
rect 26739 9284 26740 9348
rect 26804 9284 26805 9348
rect 26739 9283 26805 9284
rect 23990 8672 23998 8736
rect 24062 8672 24078 8736
rect 24142 8672 24158 8736
rect 24222 8672 24238 8736
rect 24302 8672 24310 8736
rect 21035 7988 21101 7989
rect 21035 7924 21036 7988
rect 21100 7924 21101 7988
rect 21035 7923 21101 7924
rect 20149 7040 20157 7104
rect 20221 7040 20237 7104
rect 20301 7040 20317 7104
rect 20381 7040 20397 7104
rect 20461 7040 20469 7104
rect 18643 6764 18709 6765
rect 18643 6700 18644 6764
rect 18708 6700 18709 6764
rect 18643 6699 18709 6700
rect 16308 6496 16316 6560
rect 16380 6496 16396 6560
rect 16460 6496 16476 6560
rect 16540 6496 16556 6560
rect 16620 6496 16628 6560
rect 16308 5472 16628 6496
rect 16308 5408 16316 5472
rect 16380 5408 16396 5472
rect 16460 5408 16476 5472
rect 16540 5408 16556 5472
rect 16620 5408 16628 5472
rect 15699 4724 15765 4725
rect 15699 4660 15700 4724
rect 15764 4660 15765 4724
rect 15699 4659 15765 4660
rect 12467 3776 12475 3840
rect 12539 3776 12555 3840
rect 12619 3776 12635 3840
rect 12699 3776 12715 3840
rect 12779 3776 12787 3840
rect 12467 2752 12787 3776
rect 12467 2688 12475 2752
rect 12539 2688 12555 2752
rect 12619 2688 12635 2752
rect 12699 2688 12715 2752
rect 12779 2688 12787 2752
rect 12467 2128 12787 2688
rect 16308 4384 16628 5408
rect 16308 4320 16316 4384
rect 16380 4320 16396 4384
rect 16460 4320 16476 4384
rect 16540 4320 16556 4384
rect 16620 4320 16628 4384
rect 16308 3296 16628 4320
rect 16308 3232 16316 3296
rect 16380 3232 16396 3296
rect 16460 3232 16476 3296
rect 16540 3232 16556 3296
rect 16620 3232 16628 3296
rect 16308 2208 16628 3232
rect 16308 2144 16316 2208
rect 16380 2144 16396 2208
rect 16460 2144 16476 2208
rect 16540 2144 16556 2208
rect 16620 2144 16628 2208
rect 16308 2128 16628 2144
rect 20149 6016 20469 7040
rect 20149 5952 20157 6016
rect 20221 5952 20237 6016
rect 20301 5952 20317 6016
rect 20381 5952 20397 6016
rect 20461 5952 20469 6016
rect 20149 4928 20469 5952
rect 20149 4864 20157 4928
rect 20221 4864 20237 4928
rect 20301 4864 20317 4928
rect 20381 4864 20397 4928
rect 20461 4864 20469 4928
rect 20149 3840 20469 4864
rect 20149 3776 20157 3840
rect 20221 3776 20237 3840
rect 20301 3776 20317 3840
rect 20381 3776 20397 3840
rect 20461 3776 20469 3840
rect 20149 2752 20469 3776
rect 20149 2688 20157 2752
rect 20221 2688 20237 2752
rect 20301 2688 20317 2752
rect 20381 2688 20397 2752
rect 20461 2688 20469 2752
rect 20149 2128 20469 2688
rect 23990 7648 24310 8672
rect 23990 7584 23998 7648
rect 24062 7584 24078 7648
rect 24142 7584 24158 7648
rect 24222 7584 24238 7648
rect 24302 7584 24310 7648
rect 23990 6560 24310 7584
rect 23990 6496 23998 6560
rect 24062 6496 24078 6560
rect 24142 6496 24158 6560
rect 24222 6496 24238 6560
rect 24302 6496 24310 6560
rect 23990 5472 24310 6496
rect 23990 5408 23998 5472
rect 24062 5408 24078 5472
rect 24142 5408 24158 5472
rect 24222 5408 24238 5472
rect 24302 5408 24310 5472
rect 23990 4384 24310 5408
rect 23990 4320 23998 4384
rect 24062 4320 24078 4384
rect 24142 4320 24158 4384
rect 24222 4320 24238 4384
rect 24302 4320 24310 4384
rect 23990 3296 24310 4320
rect 23990 3232 23998 3296
rect 24062 3232 24078 3296
rect 24142 3232 24158 3296
rect 24222 3232 24238 3296
rect 24302 3232 24310 3296
rect 23990 2208 24310 3232
rect 23990 2144 23998 2208
rect 24062 2144 24078 2208
rect 24142 2144 24158 2208
rect 24222 2144 24238 2208
rect 24302 2144 24310 2208
rect 23990 2128 24310 2144
rect 27831 9280 28151 10304
rect 27831 9216 27839 9280
rect 27903 9216 27919 9280
rect 27983 9216 27999 9280
rect 28063 9216 28079 9280
rect 28143 9216 28151 9280
rect 27831 8192 28151 9216
rect 27831 8128 27839 8192
rect 27903 8128 27919 8192
rect 27983 8128 27999 8192
rect 28063 8128 28079 8192
rect 28143 8128 28151 8192
rect 27831 7104 28151 8128
rect 27831 7040 27839 7104
rect 27903 7040 27919 7104
rect 27983 7040 27999 7104
rect 28063 7040 28079 7104
rect 28143 7040 28151 7104
rect 27831 6016 28151 7040
rect 28766 6221 28826 16530
rect 28947 16492 28948 16530
rect 29012 16492 29013 16556
rect 28947 16491 29013 16492
rect 29134 15874 29194 16763
rect 28950 15814 29194 15874
rect 28950 12749 29010 15814
rect 29131 15604 29197 15605
rect 29131 15540 29132 15604
rect 29196 15540 29197 15604
rect 29131 15539 29197 15540
rect 28947 12748 29013 12749
rect 28947 12684 28948 12748
rect 29012 12684 29013 12748
rect 28947 12683 29013 12684
rect 29134 9210 29194 15539
rect 29318 14789 29378 19075
rect 29502 16693 29562 19483
rect 29686 17645 29746 20707
rect 30238 20501 30298 22747
rect 30422 21725 30482 26419
rect 30790 26077 30850 31179
rect 31672 30496 31992 31520
rect 32259 31380 32325 31381
rect 32259 31316 32260 31380
rect 32324 31316 32325 31380
rect 32259 31315 32325 31316
rect 31672 30432 31680 30496
rect 31744 30432 31760 30496
rect 31824 30432 31840 30496
rect 31904 30432 31920 30496
rect 31984 30432 31992 30496
rect 31155 29612 31221 29613
rect 31155 29548 31156 29612
rect 31220 29548 31221 29612
rect 31155 29547 31221 29548
rect 30971 27436 31037 27437
rect 30971 27372 30972 27436
rect 31036 27372 31037 27436
rect 30971 27371 31037 27372
rect 30787 26076 30853 26077
rect 30787 26012 30788 26076
rect 30852 26012 30853 26076
rect 30787 26011 30853 26012
rect 30603 25668 30669 25669
rect 30603 25604 30604 25668
rect 30668 25604 30669 25668
rect 30603 25603 30669 25604
rect 30606 25261 30666 25603
rect 30603 25260 30669 25261
rect 30603 25196 30604 25260
rect 30668 25196 30669 25260
rect 30603 25195 30669 25196
rect 30419 21724 30485 21725
rect 30419 21660 30420 21724
rect 30484 21660 30485 21724
rect 30419 21659 30485 21660
rect 30422 20909 30482 21659
rect 30790 21453 30850 26011
rect 30974 21997 31034 27371
rect 31158 25397 31218 29547
rect 31672 29408 31992 30432
rect 31672 29344 31680 29408
rect 31744 29344 31760 29408
rect 31824 29344 31840 29408
rect 31904 29344 31920 29408
rect 31984 29344 31992 29408
rect 31523 29068 31589 29069
rect 31523 29004 31524 29068
rect 31588 29004 31589 29068
rect 31523 29003 31589 29004
rect 31339 28388 31405 28389
rect 31339 28324 31340 28388
rect 31404 28324 31405 28388
rect 31339 28323 31405 28324
rect 31155 25396 31221 25397
rect 31155 25332 31156 25396
rect 31220 25332 31221 25396
rect 31155 25331 31221 25332
rect 31155 24988 31221 24989
rect 31155 24924 31156 24988
rect 31220 24924 31221 24988
rect 31155 24923 31221 24924
rect 30971 21996 31037 21997
rect 30971 21932 30972 21996
rect 31036 21932 31037 21996
rect 30971 21931 31037 21932
rect 30971 21860 31037 21861
rect 30971 21796 30972 21860
rect 31036 21796 31037 21860
rect 30971 21795 31037 21796
rect 30603 21452 30669 21453
rect 30603 21388 30604 21452
rect 30668 21388 30669 21452
rect 30603 21387 30669 21388
rect 30787 21452 30853 21453
rect 30787 21388 30788 21452
rect 30852 21388 30853 21452
rect 30787 21387 30853 21388
rect 30419 20908 30485 20909
rect 30419 20844 30420 20908
rect 30484 20844 30485 20908
rect 30419 20843 30485 20844
rect 30235 20500 30301 20501
rect 30235 20436 30236 20500
rect 30300 20436 30301 20500
rect 30235 20435 30301 20436
rect 30051 20228 30117 20229
rect 30051 20164 30052 20228
rect 30116 20164 30117 20228
rect 30051 20163 30117 20164
rect 29867 19412 29933 19413
rect 29867 19348 29868 19412
rect 29932 19348 29933 19412
rect 29867 19347 29933 19348
rect 29683 17644 29749 17645
rect 29683 17580 29684 17644
rect 29748 17580 29749 17644
rect 29683 17579 29749 17580
rect 29499 16692 29565 16693
rect 29499 16628 29500 16692
rect 29564 16690 29565 16692
rect 29564 16630 29746 16690
rect 29564 16628 29565 16630
rect 29499 16627 29565 16628
rect 29499 16556 29565 16557
rect 29499 16492 29500 16556
rect 29564 16492 29565 16556
rect 29499 16491 29565 16492
rect 29315 14788 29381 14789
rect 29315 14724 29316 14788
rect 29380 14724 29381 14788
rect 29315 14723 29381 14724
rect 29502 13021 29562 16491
rect 29686 14653 29746 16630
rect 29683 14652 29749 14653
rect 29683 14588 29684 14652
rect 29748 14588 29749 14652
rect 29683 14587 29749 14588
rect 29870 13837 29930 19347
rect 30054 16693 30114 20163
rect 30419 19684 30485 19685
rect 30419 19620 30420 19684
rect 30484 19620 30485 19684
rect 30419 19619 30485 19620
rect 30235 19412 30301 19413
rect 30235 19348 30236 19412
rect 30300 19348 30301 19412
rect 30235 19347 30301 19348
rect 30238 17917 30298 19347
rect 30422 18597 30482 19619
rect 30419 18596 30485 18597
rect 30419 18532 30420 18596
rect 30484 18532 30485 18596
rect 30419 18531 30485 18532
rect 30235 17916 30301 17917
rect 30235 17852 30236 17916
rect 30300 17852 30301 17916
rect 30235 17851 30301 17852
rect 30235 17372 30301 17373
rect 30235 17308 30236 17372
rect 30300 17308 30301 17372
rect 30235 17307 30301 17308
rect 30051 16692 30117 16693
rect 30051 16628 30052 16692
rect 30116 16628 30117 16692
rect 30051 16627 30117 16628
rect 30051 16556 30117 16557
rect 30051 16492 30052 16556
rect 30116 16492 30117 16556
rect 30051 16491 30117 16492
rect 29867 13836 29933 13837
rect 29867 13772 29868 13836
rect 29932 13772 29933 13836
rect 29867 13771 29933 13772
rect 29499 13020 29565 13021
rect 29499 12956 29500 13020
rect 29564 12956 29565 13020
rect 29499 12955 29565 12956
rect 28950 9150 29194 9210
rect 28950 8805 29010 9150
rect 28947 8804 29013 8805
rect 28947 8740 28948 8804
rect 29012 8740 29013 8804
rect 28947 8739 29013 8740
rect 28763 6220 28829 6221
rect 28763 6156 28764 6220
rect 28828 6156 28829 6220
rect 28763 6155 28829 6156
rect 27831 5952 27839 6016
rect 27903 5952 27919 6016
rect 27983 5952 27999 6016
rect 28063 5952 28079 6016
rect 28143 5952 28151 6016
rect 27831 4928 28151 5952
rect 28950 5269 29010 8739
rect 30054 8669 30114 16491
rect 30238 15333 30298 17307
rect 30422 16013 30482 18531
rect 30606 16965 30666 21387
rect 30790 19549 30850 21387
rect 30787 19548 30853 19549
rect 30787 19484 30788 19548
rect 30852 19484 30853 19548
rect 30787 19483 30853 19484
rect 30603 16964 30669 16965
rect 30603 16900 30604 16964
rect 30668 16900 30669 16964
rect 30603 16899 30669 16900
rect 30790 16013 30850 19483
rect 30974 16693 31034 21795
rect 31158 21725 31218 24923
rect 31342 23357 31402 28323
rect 31526 27573 31586 29003
rect 31672 28320 31992 29344
rect 31672 28256 31680 28320
rect 31744 28256 31760 28320
rect 31824 28256 31840 28320
rect 31904 28256 31920 28320
rect 31984 28256 31992 28320
rect 31523 27572 31589 27573
rect 31523 27508 31524 27572
rect 31588 27508 31589 27572
rect 31523 27507 31589 27508
rect 31339 23356 31405 23357
rect 31339 23292 31340 23356
rect 31404 23292 31405 23356
rect 31339 23291 31405 23292
rect 31155 21724 31221 21725
rect 31155 21660 31156 21724
rect 31220 21660 31221 21724
rect 31155 21659 31221 21660
rect 31155 20772 31221 20773
rect 31155 20708 31156 20772
rect 31220 20708 31221 20772
rect 31155 20707 31221 20708
rect 30971 16692 31037 16693
rect 30971 16628 30972 16692
rect 31036 16628 31037 16692
rect 30971 16627 31037 16628
rect 30419 16012 30485 16013
rect 30419 15948 30420 16012
rect 30484 15948 30485 16012
rect 30419 15947 30485 15948
rect 30787 16012 30853 16013
rect 30787 15948 30788 16012
rect 30852 15948 30853 16012
rect 30787 15947 30853 15948
rect 30235 15332 30301 15333
rect 30235 15268 30236 15332
rect 30300 15268 30301 15332
rect 30235 15267 30301 15268
rect 30422 10845 30482 15947
rect 31158 13565 31218 20707
rect 31339 18732 31405 18733
rect 31339 18668 31340 18732
rect 31404 18668 31405 18732
rect 31339 18667 31405 18668
rect 31155 13564 31221 13565
rect 31155 13500 31156 13564
rect 31220 13500 31221 13564
rect 31155 13499 31221 13500
rect 31342 10981 31402 18667
rect 31526 17101 31586 27507
rect 31672 27232 31992 28256
rect 32075 27980 32141 27981
rect 32075 27916 32076 27980
rect 32140 27916 32141 27980
rect 32075 27915 32141 27916
rect 31672 27168 31680 27232
rect 31744 27168 31760 27232
rect 31824 27168 31840 27232
rect 31904 27168 31920 27232
rect 31984 27168 31992 27232
rect 31672 26144 31992 27168
rect 31672 26080 31680 26144
rect 31744 26080 31760 26144
rect 31824 26080 31840 26144
rect 31904 26080 31920 26144
rect 31984 26080 31992 26144
rect 31672 25056 31992 26080
rect 32078 25533 32138 27915
rect 32075 25532 32141 25533
rect 32075 25468 32076 25532
rect 32140 25468 32141 25532
rect 32075 25467 32141 25468
rect 31672 24992 31680 25056
rect 31744 24992 31760 25056
rect 31824 24992 31840 25056
rect 31904 24992 31920 25056
rect 31984 24992 31992 25056
rect 31672 23968 31992 24992
rect 32262 24717 32322 31315
rect 32627 30020 32693 30021
rect 32627 29956 32628 30020
rect 32692 29956 32693 30020
rect 32627 29955 32693 29956
rect 32443 28796 32509 28797
rect 32443 28732 32444 28796
rect 32508 28732 32509 28796
rect 32443 28731 32509 28732
rect 32446 25397 32506 28731
rect 32443 25396 32509 25397
rect 32443 25332 32444 25396
rect 32508 25332 32509 25396
rect 32443 25331 32509 25332
rect 32630 25261 32690 29955
rect 32627 25260 32693 25261
rect 32627 25196 32628 25260
rect 32692 25196 32693 25260
rect 32627 25195 32693 25196
rect 32259 24716 32325 24717
rect 32259 24652 32260 24716
rect 32324 24652 32325 24716
rect 32259 24651 32325 24652
rect 31672 23904 31680 23968
rect 31744 23904 31760 23968
rect 31824 23904 31840 23968
rect 31904 23904 31920 23968
rect 31984 23904 31992 23968
rect 31672 22880 31992 23904
rect 31672 22816 31680 22880
rect 31744 22816 31760 22880
rect 31824 22816 31840 22880
rect 31904 22816 31920 22880
rect 31984 22816 31992 22880
rect 31672 21792 31992 22816
rect 31672 21728 31680 21792
rect 31744 21728 31760 21792
rect 31824 21728 31840 21792
rect 31904 21728 31920 21792
rect 31984 21728 31992 21792
rect 31672 20704 31992 21728
rect 31672 20640 31680 20704
rect 31744 20640 31760 20704
rect 31824 20640 31840 20704
rect 31904 20640 31920 20704
rect 31984 20640 31992 20704
rect 31672 19616 31992 20640
rect 31672 19552 31680 19616
rect 31744 19552 31760 19616
rect 31824 19552 31840 19616
rect 31904 19552 31920 19616
rect 31984 19552 31992 19616
rect 31672 18528 31992 19552
rect 31672 18464 31680 18528
rect 31744 18464 31760 18528
rect 31824 18464 31840 18528
rect 31904 18464 31920 18528
rect 31984 18464 31992 18528
rect 31672 17440 31992 18464
rect 31672 17376 31680 17440
rect 31744 17376 31760 17440
rect 31824 17376 31840 17440
rect 31904 17376 31920 17440
rect 31984 17376 31992 17440
rect 31523 17100 31589 17101
rect 31523 17036 31524 17100
rect 31588 17036 31589 17100
rect 31523 17035 31589 17036
rect 31526 15197 31586 17035
rect 31672 16352 31992 17376
rect 31672 16288 31680 16352
rect 31744 16288 31760 16352
rect 31824 16288 31840 16352
rect 31904 16288 31920 16352
rect 31984 16288 31992 16352
rect 31672 15264 31992 16288
rect 31672 15200 31680 15264
rect 31744 15200 31760 15264
rect 31824 15200 31840 15264
rect 31904 15200 31920 15264
rect 31984 15200 31992 15264
rect 31523 15196 31589 15197
rect 31523 15132 31524 15196
rect 31588 15132 31589 15196
rect 31523 15131 31589 15132
rect 31672 14176 31992 15200
rect 31672 14112 31680 14176
rect 31744 14112 31760 14176
rect 31824 14112 31840 14176
rect 31904 14112 31920 14176
rect 31984 14112 31992 14176
rect 31672 13088 31992 14112
rect 31672 13024 31680 13088
rect 31744 13024 31760 13088
rect 31824 13024 31840 13088
rect 31904 13024 31920 13088
rect 31984 13024 31992 13088
rect 31672 12000 31992 13024
rect 31672 11936 31680 12000
rect 31744 11936 31760 12000
rect 31824 11936 31840 12000
rect 31904 11936 31920 12000
rect 31984 11936 31992 12000
rect 31339 10980 31405 10981
rect 31339 10916 31340 10980
rect 31404 10916 31405 10980
rect 31339 10915 31405 10916
rect 31672 10912 31992 11936
rect 31672 10848 31680 10912
rect 31744 10848 31760 10912
rect 31824 10848 31840 10912
rect 31904 10848 31920 10912
rect 31984 10848 31992 10912
rect 30419 10844 30485 10845
rect 30419 10780 30420 10844
rect 30484 10780 30485 10844
rect 30419 10779 30485 10780
rect 31672 9824 31992 10848
rect 31672 9760 31680 9824
rect 31744 9760 31760 9824
rect 31824 9760 31840 9824
rect 31904 9760 31920 9824
rect 31984 9760 31992 9824
rect 31672 8736 31992 9760
rect 31672 8672 31680 8736
rect 31744 8672 31760 8736
rect 31824 8672 31840 8736
rect 31904 8672 31920 8736
rect 31984 8672 31992 8736
rect 29683 8668 29749 8669
rect 29683 8604 29684 8668
rect 29748 8604 29749 8668
rect 29683 8603 29749 8604
rect 30051 8668 30117 8669
rect 30051 8604 30052 8668
rect 30116 8604 30117 8668
rect 30051 8603 30117 8604
rect 28947 5268 29013 5269
rect 28947 5204 28948 5268
rect 29012 5204 29013 5268
rect 28947 5203 29013 5204
rect 27831 4864 27839 4928
rect 27903 4864 27919 4928
rect 27983 4864 27999 4928
rect 28063 4864 28079 4928
rect 28143 4864 28151 4928
rect 27831 3840 28151 4864
rect 29686 4725 29746 8603
rect 31672 7648 31992 8672
rect 31672 7584 31680 7648
rect 31744 7584 31760 7648
rect 31824 7584 31840 7648
rect 31904 7584 31920 7648
rect 31984 7584 31992 7648
rect 31672 6560 31992 7584
rect 31672 6496 31680 6560
rect 31744 6496 31760 6560
rect 31824 6496 31840 6560
rect 31904 6496 31920 6560
rect 31984 6496 31992 6560
rect 31672 5472 31992 6496
rect 31672 5408 31680 5472
rect 31744 5408 31760 5472
rect 31824 5408 31840 5472
rect 31904 5408 31920 5472
rect 31984 5408 31992 5472
rect 29683 4724 29749 4725
rect 29683 4660 29684 4724
rect 29748 4660 29749 4724
rect 29683 4659 29749 4660
rect 27831 3776 27839 3840
rect 27903 3776 27919 3840
rect 27983 3776 27999 3840
rect 28063 3776 28079 3840
rect 28143 3776 28151 3840
rect 27831 2752 28151 3776
rect 27831 2688 27839 2752
rect 27903 2688 27919 2752
rect 27983 2688 27999 2752
rect 28063 2688 28079 2752
rect 28143 2688 28151 2752
rect 27831 2128 28151 2688
rect 31672 4384 31992 5408
rect 31672 4320 31680 4384
rect 31744 4320 31760 4384
rect 31824 4320 31840 4384
rect 31904 4320 31920 4384
rect 31984 4320 31992 4384
rect 31672 3296 31992 4320
rect 31672 3232 31680 3296
rect 31744 3232 31760 3296
rect 31824 3232 31840 3296
rect 31904 3232 31920 3296
rect 31984 3232 31992 3296
rect 31672 2208 31992 3232
rect 31672 2144 31680 2208
rect 31744 2144 31760 2208
rect 31824 2144 31840 2208
rect 31904 2144 31920 2208
rect 31984 2144 31992 2208
rect 31672 2128 31992 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13616 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0439__B
timestamp 1666464484
transform -1 0 15824 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0440__B
timestamp 1666464484
transform 1 0 17388 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0442__B
timestamp 1666464484
transform 1 0 14352 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0445__A
timestamp 1666464484
transform 1 0 12052 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__A
timestamp 1666464484
transform 1 0 15088 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__A
timestamp 1666464484
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__B
timestamp 1666464484
transform 1 0 16192 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0449__A
timestamp 1666464484
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__A
timestamp 1666464484
transform 1 0 17480 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0453__A
timestamp 1666464484
transform 1 0 17572 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0453__B
timestamp 1666464484
transform 1 0 17940 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__A
timestamp 1666464484
transform -1 0 13248 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__B
timestamp 1666464484
transform -1 0 12144 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__A
timestamp 1666464484
transform 1 0 10488 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__B
timestamp 1666464484
transform -1 0 28336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__D
timestamp 1666464484
transform -1 0 29072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__A1
timestamp 1666464484
transform 1 0 18216 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__B1
timestamp 1666464484
transform -1 0 19136 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__A
timestamp 1666464484
transform -1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__B
timestamp 1666464484
transform 1 0 11960 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__C
timestamp 1666464484
transform 1 0 13064 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__B
timestamp 1666464484
transform 1 0 8832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__A1
timestamp 1666464484
transform 1 0 16744 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0461__A
timestamp 1666464484
transform 1 0 15824 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__A
timestamp 1666464484
transform 1 0 14444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__A
timestamp 1666464484
transform 1 0 14628 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__B
timestamp 1666464484
transform 1 0 13616 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__A1
timestamp 1666464484
transform 1 0 8280 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__A2
timestamp 1666464484
transform -1 0 9016 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__C1
timestamp 1666464484
transform -1 0 8096 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__A
timestamp 1666464484
transform 1 0 9384 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__A
timestamp 1666464484
transform 1 0 14536 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__B
timestamp 1666464484
transform 1 0 9752 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__D
timestamp 1666464484
transform 1 0 10856 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__A1
timestamp 1666464484
transform -1 0 20700 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__A2
timestamp 1666464484
transform -1 0 21252 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__A3
timestamp 1666464484
transform -1 0 19872 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__B
timestamp 1666464484
transform 1 0 8280 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0472__B1
timestamp 1666464484
transform 1 0 10488 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__B
timestamp 1666464484
transform 1 0 11408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0474__B
timestamp 1666464484
transform -1 0 10120 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__B
timestamp 1666464484
transform 1 0 12512 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__A
timestamp 1666464484
transform 1 0 10304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__B
timestamp 1666464484
transform 1 0 9936 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__A
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__C
timestamp 1666464484
transform 1 0 28244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__A
timestamp 1666464484
transform 1 0 11040 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__A
timestamp 1666464484
transform 1 0 9200 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__B
timestamp 1666464484
transform 1 0 8832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__C
timestamp 1666464484
transform 1 0 10488 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__A
timestamp 1666464484
transform 1 0 28796 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__B
timestamp 1666464484
transform -1 0 29532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__A1
timestamp 1666464484
transform -1 0 5336 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__A2
timestamp 1666464484
transform -1 0 30452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A1
timestamp 1666464484
transform 1 0 11776 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__B1
timestamp 1666464484
transform -1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__A
timestamp 1666464484
transform -1 0 27784 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__B
timestamp 1666464484
transform 1 0 26036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__A
timestamp 1666464484
transform -1 0 28888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__A
timestamp 1666464484
transform 1 0 29716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__A1
timestamp 1666464484
transform 1 0 25484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__B1
timestamp 1666464484
transform 1 0 25852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1666464484
transform -1 0 28336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__B
timestamp 1666464484
transform 1 0 27140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__B1
timestamp 1666464484
transform 1 0 27232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A
timestamp 1666464484
transform -1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A
timestamp 1666464484
transform -1 0 31188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__A1
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__B1
timestamp 1666464484
transform 1 0 26404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1666464484
transform -1 0 29532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__B
timestamp 1666464484
transform -1 0 28336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__A
timestamp 1666464484
transform -1 0 9016 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__C
timestamp 1666464484
transform 1 0 20148 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__D
timestamp 1666464484
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__A
timestamp 1666464484
transform -1 0 7544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__C
timestamp 1666464484
transform 1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__D
timestamp 1666464484
transform 1 0 9292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__C
timestamp 1666464484
transform -1 0 27324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A
timestamp 1666464484
transform -1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__A
timestamp 1666464484
transform -1 0 30636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__B
timestamp 1666464484
transform -1 0 30084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__A1
timestamp 1666464484
transform 1 0 7636 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__A2
timestamp 1666464484
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__B1
timestamp 1666464484
transform -1 0 8372 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__A
timestamp 1666464484
transform -1 0 7544 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__B
timestamp 1666464484
transform 1 0 9292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__C
timestamp 1666464484
transform -1 0 8924 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1666464484
transform -1 0 25484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__B
timestamp 1666464484
transform -1 0 26036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__A
timestamp 1666464484
transform 1 0 23736 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__A1
timestamp 1666464484
transform -1 0 7268 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__A2
timestamp 1666464484
transform 1 0 7912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__B1
timestamp 1666464484
transform 1 0 6808 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A1
timestamp 1666464484
transform 1 0 7912 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A2
timestamp 1666464484
transform 1 0 7360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A1
timestamp 1666464484
transform -1 0 6440 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A2
timestamp 1666464484
transform -1 0 5520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__B1
timestamp 1666464484
transform -1 0 6440 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A1
timestamp 1666464484
transform 1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A2
timestamp 1666464484
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1666464484
transform 1 0 12880 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A1
timestamp 1666464484
transform 1 0 18032 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__B1
timestamp 1666464484
transform 1 0 10764 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__A
timestamp 1666464484
transform -1 0 18400 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__B
timestamp 1666464484
transform 1 0 18768 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1666464484
transform 1 0 9752 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__B
timestamp 1666464484
transform 1 0 10764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1666464484
transform 1 0 26772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1666464484
transform -1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__A
timestamp 1666464484
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__B
timestamp 1666464484
transform -1 0 9384 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1666464484
transform -1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__B
timestamp 1666464484
transform -1 0 7544 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__B2
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A1
timestamp 1666464484
transform 1 0 10396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A2
timestamp 1666464484
transform 1 0 10948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A3
timestamp 1666464484
transform -1 0 19596 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A
timestamp 1666464484
transform 1 0 9384 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__B
timestamp 1666464484
transform 1 0 9016 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__D
timestamp 1666464484
transform 1 0 9936 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__C
timestamp 1666464484
transform 1 0 23920 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A
timestamp 1666464484
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A
timestamp 1666464484
transform -1 0 24748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A
timestamp 1666464484
transform -1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__B
timestamp 1666464484
transform -1 0 31096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A1
timestamp 1666464484
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__C1
timestamp 1666464484
transform 1 0 10948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__C1
timestamp 1666464484
transform -1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1666464484
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B
timestamp 1666464484
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1666464484
transform -1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A2
timestamp 1666464484
transform 1 0 24472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__B
timestamp 1666464484
transform -1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A1
timestamp 1666464484
transform 1 0 27784 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A2
timestamp 1666464484
transform 1 0 25116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A2
timestamp 1666464484
transform -1 0 10488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A3
timestamp 1666464484
transform -1 0 10672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__B
timestamp 1666464484
transform 1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__C
timestamp 1666464484
transform 1 0 17480 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A2
timestamp 1666464484
transform 1 0 25300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A3
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C
timestamp 1666464484
transform 1 0 26220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A2
timestamp 1666464484
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B1
timestamp 1666464484
transform 1 0 12880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1666464484
transform -1 0 28980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__C
timestamp 1666464484
transform -1 0 29164 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B
timestamp 1666464484
transform -1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__B
timestamp 1666464484
transform -1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A2
timestamp 1666464484
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__C1
timestamp 1666464484
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 1666464484
transform 1 0 8832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__B
timestamp 1666464484
transform -1 0 9568 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A1_N
timestamp 1666464484
transform 1 0 7176 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A2_N
timestamp 1666464484
transform -1 0 5520 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__B1
timestamp 1666464484
transform -1 0 5336 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A
timestamp 1666464484
transform 1 0 10856 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__B
timestamp 1666464484
transform -1 0 7912 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__C
timestamp 1666464484
transform 1 0 9200 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1666464484
transform -1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A
timestamp 1666464484
transform -1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__B
timestamp 1666464484
transform 1 0 10856 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A1
timestamp 1666464484
transform 1 0 5888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B2
timestamp 1666464484
transform 1 0 9752 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1666464484
transform -1 0 14168 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__B
timestamp 1666464484
transform 1 0 11040 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 1666464484
transform -1 0 12604 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__B1
timestamp 1666464484
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__C1
timestamp 1666464484
transform 1 0 28980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A
timestamp 1666464484
transform 1 0 18400 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A1
timestamp 1666464484
transform 1 0 14536 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A2
timestamp 1666464484
transform 1 0 11960 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__B1
timestamp 1666464484
transform 1 0 14904 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__B
timestamp 1666464484
transform 1 0 10304 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__C
timestamp 1666464484
transform 1 0 12328 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1666464484
transform -1 0 18400 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A1
timestamp 1666464484
transform 1 0 7360 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B1
timestamp 1666464484
transform 1 0 9384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__C1
timestamp 1666464484
transform 1 0 11040 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A
timestamp 1666464484
transform 1 0 12512 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B
timestamp 1666464484
transform -1 0 13800 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A1
timestamp 1666464484
transform -1 0 28888 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__C1
timestamp 1666464484
transform -1 0 27324 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1666464484
transform 1 0 28244 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B
timestamp 1666464484
transform -1 0 26680 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__C
timestamp 1666464484
transform -1 0 27232 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A1
timestamp 1666464484
transform 1 0 16928 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B1
timestamp 1666464484
transform 1 0 17664 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__C1
timestamp 1666464484
transform 1 0 12328 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A2
timestamp 1666464484
transform -1 0 6992 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__C1
timestamp 1666464484
transform -1 0 7912 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A1
timestamp 1666464484
transform 1 0 12880 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A2
timestamp 1666464484
transform 1 0 9936 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B1
timestamp 1666464484
transform 1 0 15456 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__C1
timestamp 1666464484
transform 1 0 10856 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1666464484
transform 1 0 11960 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1666464484
transform 1 0 15088 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1666464484
transform 1 0 9384 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B
timestamp 1666464484
transform -1 0 8464 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1666464484
transform -1 0 7544 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__B
timestamp 1666464484
transform -1 0 8096 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__C
timestamp 1666464484
transform -1 0 9384 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1666464484
transform 1 0 13248 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B
timestamp 1666464484
transform -1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1666464484
transform -1 0 17296 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__C
timestamp 1666464484
transform -1 0 18400 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1666464484
transform 1 0 11408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A1
timestamp 1666464484
transform 1 0 6624 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A1
timestamp 1666464484
transform 1 0 28796 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A2
timestamp 1666464484
transform -1 0 27784 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B1
timestamp 1666464484
transform 1 0 11040 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__C1
timestamp 1666464484
transform 1 0 10304 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A1
timestamp 1666464484
transform 1 0 7176 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__C1
timestamp 1666464484
transform -1 0 8464 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A1
timestamp 1666464484
transform 1 0 30176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__C1
timestamp 1666464484
transform 1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1666464484
transform 1 0 29532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 1666464484
transform -1 0 30544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1666464484
transform 1 0 14628 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B
timestamp 1666464484
transform 1 0 17664 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1666464484
transform -1 0 6992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B
timestamp 1666464484
transform 1 0 6992 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A1
timestamp 1666464484
transform -1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A2
timestamp 1666464484
transform -1 0 19688 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B1
timestamp 1666464484
transform -1 0 18952 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A1
timestamp 1666464484
transform 1 0 27324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1666464484
transform -1 0 24748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1666464484
transform 1 0 15088 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B
timestamp 1666464484
transform -1 0 17848 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1666464484
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B
timestamp 1666464484
transform -1 0 9936 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1666464484
transform 1 0 10488 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B
timestamp 1666464484
transform 1 0 13064 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B
timestamp 1666464484
transform -1 0 17848 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__C
timestamp 1666464484
transform 1 0 13432 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__D
timestamp 1666464484
transform 1 0 14720 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1666464484
transform 1 0 7912 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B
timestamp 1666464484
transform -1 0 7728 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__C
timestamp 1666464484
transform 1 0 9476 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__D
timestamp 1666464484
transform 1 0 8832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A2
timestamp 1666464484
transform -1 0 6440 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A3
timestamp 1666464484
transform -1 0 6992 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B1
timestamp 1666464484
transform -1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1666464484
transform 1 0 11776 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A2
timestamp 1666464484
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B1
timestamp 1666464484
transform 1 0 24748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1666464484
transform -1 0 30084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__C
timestamp 1666464484
transform -1 0 30636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1666464484
transform -1 0 28520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B
timestamp 1666464484
transform -1 0 28060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__C_N
timestamp 1666464484
transform -1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A
timestamp 1666464484
transform -1 0 14996 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B
timestamp 1666464484
transform -1 0 11960 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A2
timestamp 1666464484
transform -1 0 28520 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A3
timestamp 1666464484
transform -1 0 28980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A4
timestamp 1666464484
transform -1 0 27324 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A
timestamp 1666464484
transform -1 0 7912 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B
timestamp 1666464484
transform 1 0 10304 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__D
timestamp 1666464484
transform -1 0 8096 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B
timestamp 1666464484
transform -1 0 5888 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__C_N
timestamp 1666464484
transform -1 0 9568 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A2
timestamp 1666464484
transform -1 0 23000 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A3
timestamp 1666464484
transform -1 0 23184 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B
timestamp 1666464484
transform 1 0 8464 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__C
timestamp 1666464484
transform 1 0 5704 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1666464484
transform 1 0 11040 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B
timestamp 1666464484
transform -1 0 12144 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A
timestamp 1666464484
transform -1 0 14444 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B
timestamp 1666464484
transform 1 0 13432 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A2
timestamp 1666464484
transform -1 0 6992 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B1
timestamp 1666464484
transform 1 0 5888 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__C1
timestamp 1666464484
transform 1 0 6256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1666464484
transform -1 0 20976 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1666464484
transform -1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__C
timestamp 1666464484
transform 1 0 11776 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A
timestamp 1666464484
transform 1 0 18584 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B
timestamp 1666464484
transform 1 0 13064 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 1666464484
transform 1 0 14996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 1666464484
transform 1 0 13984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__C
timestamp 1666464484
transform -1 0 9568 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1666464484
transform 1 0 29716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__C
timestamp 1666464484
transform 1 0 27324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1666464484
transform -1 0 10120 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B
timestamp 1666464484
transform -1 0 7544 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A_N
timestamp 1666464484
transform -1 0 29900 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1666464484
transform -1 0 30728 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__C
timestamp 1666464484
transform -1 0 30636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__D
timestamp 1666464484
transform -1 0 31188 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 1666464484
transform -1 0 18952 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B1
timestamp 1666464484
transform -1 0 5888 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1666464484
transform 1 0 13984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B
timestamp 1666464484
transform -1 0 17480 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A2
timestamp 1666464484
transform 1 0 7176 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B1
timestamp 1666464484
transform -1 0 5336 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__C1
timestamp 1666464484
transform -1 0 9292 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__D1
timestamp 1666464484
transform -1 0 8464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A2
timestamp 1666464484
transform -1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A1
timestamp 1666464484
transform -1 0 5888 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B1_N
timestamp 1666464484
transform -1 0 4416 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A1
timestamp 1666464484
transform 1 0 10488 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A2
timestamp 1666464484
transform 1 0 9752 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1666464484
transform 1 0 19780 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B
timestamp 1666464484
transform 1 0 16376 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__C
timestamp 1666464484
transform 1 0 15640 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1666464484
transform 1 0 8464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A0
timestamp 1666464484
transform 1 0 21988 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A1
timestamp 1666464484
transform -1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B1
timestamp 1666464484
transform 1 0 5888 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A1
timestamp 1666464484
transform 1 0 7912 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A
timestamp 1666464484
transform 1 0 11040 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1666464484
transform 1 0 6256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B
timestamp 1666464484
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__C
timestamp 1666464484
transform -1 0 7912 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1666464484
transform -1 0 4784 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B
timestamp 1666464484
transform -1 0 4968 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__C
timestamp 1666464484
transform -1 0 4416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__D
timestamp 1666464484
transform -1 0 5520 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1666464484
transform -1 0 22172 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2
timestamp 1666464484
transform 1 0 20608 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A3
timestamp 1666464484
transform -1 0 20976 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A4
timestamp 1666464484
transform -1 0 20424 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A2
timestamp 1666464484
transform 1 0 19596 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A3
timestamp 1666464484
transform 1 0 13156 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B1
timestamp 1666464484
transform 1 0 17020 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A2
timestamp 1666464484
transform -1 0 19228 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A1_N
timestamp 1666464484
transform -1 0 29900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A2_N
timestamp 1666464484
transform -1 0 29532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B1
timestamp 1666464484
transform -1 0 5336 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1666464484
transform 1 0 16468 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B
timestamp 1666464484
transform -1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1
timestamp 1666464484
transform -1 0 4968 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2
timestamp 1666464484
transform -1 0 4784 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1_N
timestamp 1666464484
transform -1 0 4232 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1
timestamp 1666464484
transform 1 0 17204 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1
timestamp 1666464484
transform -1 0 18676 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B2
timestamp 1666464484
transform -1 0 23368 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B1
timestamp 1666464484
transform 1 0 14536 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__C1
timestamp 1666464484
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A1
timestamp 1666464484
transform 1 0 11408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2
timestamp 1666464484
transform 1 0 11960 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B1
timestamp 1666464484
transform 1 0 12512 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1666464484
transform 1 0 15180 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B
timestamp 1666464484
transform 1 0 13616 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1666464484
transform 1 0 6808 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__C
timestamp 1666464484
transform -1 0 5336 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1666464484
transform 1 0 26128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A1
timestamp 1666464484
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A3
timestamp 1666464484
transform -1 0 30452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B1
timestamp 1666464484
transform 1 0 29900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__C1
timestamp 1666464484
transform 1 0 27692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1666464484
transform -1 0 30544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B
timestamp 1666464484
transform -1 0 30452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1666464484
transform 1 0 25300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B
timestamp 1666464484
transform 1 0 26496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A
timestamp 1666464484
transform 1 0 24748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1666464484
transform 1 0 8464 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__B
timestamp 1666464484
transform 1 0 10212 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B
timestamp 1666464484
transform -1 0 4232 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__C
timestamp 1666464484
transform -1 0 4968 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__D
timestamp 1666464484
transform -1 0 4784 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A1_N
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B1
timestamp 1666464484
transform 1 0 29440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A
timestamp 1666464484
transform -1 0 29900 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B
timestamp 1666464484
transform -1 0 31188 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1666464484
transform 1 0 27600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B
timestamp 1666464484
transform 1 0 26680 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B
timestamp 1666464484
transform -1 0 13064 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A
timestamp 1666464484
transform 1 0 14536 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B
timestamp 1666464484
transform 1 0 15640 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__C
timestamp 1666464484
transform -1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A2_N
timestamp 1666464484
transform -1 0 30176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B2
timestamp 1666464484
transform -1 0 30728 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1666464484
transform -1 0 6992 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B
timestamp 1666464484
transform -1 0 8096 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A1
timestamp 1666464484
transform -1 0 28060 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A2
timestamp 1666464484
transform 1 0 30452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B1
timestamp 1666464484
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B2
timestamp 1666464484
transform 1 0 27140 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A1
timestamp 1666464484
transform 1 0 30268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B2
timestamp 1666464484
transform -1 0 29900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A1
timestamp 1666464484
transform -1 0 28980 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A2
timestamp 1666464484
transform 1 0 28980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A3
timestamp 1666464484
transform 1 0 28244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1
timestamp 1666464484
transform 1 0 27324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B2
timestamp 1666464484
transform -1 0 26680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A1
timestamp 1666464484
transform 1 0 12972 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A2
timestamp 1666464484
transform -1 0 7544 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A3
timestamp 1666464484
transform -1 0 8096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1666464484
transform -1 0 6992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A2_N
timestamp 1666464484
transform 1 0 7728 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__B1
timestamp 1666464484
transform -1 0 9384 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A2
timestamp 1666464484
transform -1 0 30084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B1
timestamp 1666464484
transform -1 0 31096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A2_N
timestamp 1666464484
transform -1 0 7544 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B2
timestamp 1666464484
transform -1 0 6808 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__C1
timestamp 1666464484
transform 1 0 17848 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1666464484
transform -1 0 5520 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A2
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A3
timestamp 1666464484
transform 1 0 18124 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__B1
timestamp 1666464484
transform 1 0 14628 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A1
timestamp 1666464484
transform 1 0 15640 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__C_N
timestamp 1666464484
transform -1 0 15640 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1
timestamp 1666464484
transform 1 0 12144 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2
timestamp 1666464484
transform 1 0 21160 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A3
timestamp 1666464484
transform 1 0 21896 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1666464484
transform 1 0 25668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B
timestamp 1666464484
transform 1 0 29072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__C
timestamp 1666464484
transform 1 0 28888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__D_N
timestamp 1666464484
transform 1 0 24564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2
timestamp 1666464484
transform 1 0 11040 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A3
timestamp 1666464484
transform 1 0 9936 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B1
timestamp 1666464484
transform 1 0 10580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1666464484
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1666464484
transform 1 0 8464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A2
timestamp 1666464484
transform -1 0 30544 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A3
timestamp 1666464484
transform 1 0 5336 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A4
timestamp 1666464484
transform -1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A1
timestamp 1666464484
transform -1 0 29348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A2
timestamp 1666464484
transform -1 0 5520 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A0
timestamp 1666464484
transform -1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A1
timestamp 1666464484
transform 1 0 28704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B1
timestamp 1666464484
transform -1 0 29532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B1
timestamp 1666464484
transform -1 0 30268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B2
timestamp 1666464484
transform -1 0 30912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1666464484
transform -1 0 7544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B
timestamp 1666464484
transform -1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A1
timestamp 1666464484
transform -1 0 21988 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__B1
timestamp 1666464484
transform -1 0 28704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__C1
timestamp 1666464484
transform -1 0 28520 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A1
timestamp 1666464484
transform -1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A2
timestamp 1666464484
transform 1 0 14260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B1
timestamp 1666464484
transform 1 0 12512 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B1
timestamp 1666464484
transform 1 0 9016 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__C1
timestamp 1666464484
transform -1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__C
timestamp 1666464484
transform 1 0 7912 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A2
timestamp 1666464484
transform -1 0 6992 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1666464484
transform 1 0 9660 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B
timestamp 1666464484
transform -1 0 12788 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__C
timestamp 1666464484
transform 1 0 11316 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A1
timestamp 1666464484
transform 1 0 13432 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A2
timestamp 1666464484
transform -1 0 10120 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B1
timestamp 1666464484
transform -1 0 8464 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1666464484
transform 1 0 7912 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B
timestamp 1666464484
transform 1 0 7176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1
timestamp 1666464484
transform -1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A2
timestamp 1666464484
transform -1 0 4232 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1
timestamp 1666464484
transform -1 0 4968 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B
timestamp 1666464484
transform -1 0 15364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1666464484
transform -1 0 16744 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B
timestamp 1666464484
transform -1 0 16192 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__C
timestamp 1666464484
transform -1 0 13248 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A2
timestamp 1666464484
transform 1 0 9108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A1
timestamp 1666464484
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A2
timestamp 1666464484
transform -1 0 21160 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A3
timestamp 1666464484
transform -1 0 20608 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1666464484
transform -1 0 30084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__B
timestamp 1666464484
transform -1 0 30636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__C
timestamp 1666464484
transform -1 0 30452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A2
timestamp 1666464484
transform -1 0 13248 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A1
timestamp 1666464484
transform -1 0 11316 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__B1
timestamp 1666464484
transform 1 0 10488 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A3
timestamp 1666464484
transform -1 0 16744 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__B1
timestamp 1666464484
transform 1 0 16192 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A
timestamp 1666464484
transform -1 0 6808 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__C
timestamp 1666464484
transform -1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__D_N
timestamp 1666464484
transform 1 0 7360 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1666464484
transform -1 0 7360 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A2
timestamp 1666464484
transform -1 0 6440 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1666464484
transform 1 0 11408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B
timestamp 1666464484
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A1
timestamp 1666464484
transform 1 0 11960 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A2
timestamp 1666464484
transform 1 0 12328 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B1
timestamp 1666464484
transform -1 0 15088 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__C1
timestamp 1666464484
transform -1 0 13064 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B
timestamp 1666464484
transform -1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A1
timestamp 1666464484
transform -1 0 11868 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2
timestamp 1666464484
transform 1 0 10212 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A3
timestamp 1666464484
transform -1 0 8280 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B1
timestamp 1666464484
transform -1 0 12512 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__B
timestamp 1666464484
transform 1 0 12512 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__C
timestamp 1666464484
transform 1 0 13984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A2
timestamp 1666464484
transform 1 0 13432 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B1
timestamp 1666464484
transform -1 0 11592 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A1
timestamp 1666464484
transform 1 0 13616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B1
timestamp 1666464484
transform -1 0 17296 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B
timestamp 1666464484
transform -1 0 11592 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1666464484
transform -1 0 15272 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__B
timestamp 1666464484
transform -1 0 16192 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B
timestamp 1666464484
transform 1 0 12420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A2
timestamp 1666464484
transform 1 0 28520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A3
timestamp 1666464484
transform 1 0 28796 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B1
timestamp 1666464484
transform -1 0 27600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A2
timestamp 1666464484
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__C
timestamp 1666464484
transform 1 0 10488 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__C
timestamp 1666464484
transform 1 0 6256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__D
timestamp 1666464484
transform 1 0 7912 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A2
timestamp 1666464484
transform 1 0 12696 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A
timestamp 1666464484
transform 1 0 10488 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1666464484
transform -1 0 29900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1666464484
transform 1 0 17112 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1666464484
transform -1 0 7912 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1666464484
transform 1 0 8832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1666464484
transform 1 0 13800 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 1666464484
transform 1 0 10304 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1666464484
transform 1 0 15640 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1666464484
transform 1 0 16836 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1666464484
transform -1 0 14536 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1666464484
transform 1 0 15732 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1666464484
transform 1 0 15272 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1666464484
transform 1 0 26496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1666464484
transform -1 0 9936 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1666464484
transform 1 0 25576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1666464484
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1666464484
transform 1 0 27968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1666464484
transform -1 0 30728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A
timestamp 1666464484
transform 1 0 27416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1666464484
transform 1 0 28244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A
timestamp 1666464484
transform 1 0 30360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1666464484
transform 1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1666464484
transform 1 0 26496 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1666464484
transform -1 0 10580 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A
timestamp 1666464484
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1666464484
transform -1 0 6992 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A
timestamp 1666464484
transform -1 0 5888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1666464484
transform -1 0 7544 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1666464484
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1666464484
transform 1 0 5888 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1666464484
transform 1 0 9752 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1666464484
transform -1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A
timestamp 1666464484
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1666464484
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1666464484
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1666464484
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1666464484
transform -1 0 8464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1666464484
transform 1 0 22448 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1666464484
transform 1 0 23092 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1666464484
transform -1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1666464484
transform 1 0 22448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1666464484
transform 1 0 28796 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1666464484
transform 1 0 21804 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1666464484
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1666464484
transform 1 0 21988 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1666464484
transform 1 0 29716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1666464484
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1666464484
transform 1 0 18216 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1666464484
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1666464484
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1666464484
transform -1 0 19688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1666464484
transform -1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A
timestamp 1666464484
transform 1 0 16928 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1666464484
transform 1 0 11960 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1666464484
transform 1 0 14352 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1666464484
transform 1 0 28796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1666464484
transform -1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1666464484
transform -1 0 24472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A
timestamp 1666464484
transform -1 0 23828 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1666464484
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A
timestamp 1666464484
transform 1 0 22816 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A
timestamp 1666464484
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A
timestamp 1666464484
transform 1 0 9292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1666464484
transform 1 0 23828 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1666464484
transform 1 0 23092 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1666464484
transform -1 0 25024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A
timestamp 1666464484
transform 1 0 25944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__CLK
timestamp 1666464484
transform 1 0 9936 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__CLK
timestamp 1666464484
transform -1 0 22172 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__CLK
timestamp 1666464484
transform -1 0 27876 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__CLK
timestamp 1666464484
transform 1 0 9384 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__CLK
timestamp 1666464484
transform -1 0 6808 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__CLK
timestamp 1666464484
transform 1 0 10856 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__CLK
timestamp 1666464484
transform -1 0 25484 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__CLK
timestamp 1666464484
transform 1 0 27140 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__CLK
timestamp 1666464484
transform 1 0 28244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__CLK
timestamp 1666464484
transform 1 0 28244 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__CLK
timestamp 1666464484
transform -1 0 31372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__CLK
timestamp 1666464484
transform -1 0 31372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__CLK
timestamp 1666464484
transform 1 0 8648 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__CLK
timestamp 1666464484
transform 1 0 29072 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__CLK
timestamp 1666464484
transform -1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__CLK
timestamp 1666464484
transform 1 0 23736 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__CLK
timestamp 1666464484
transform 1 0 23920 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__CLK
timestamp 1666464484
transform 1 0 29072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout12_A
timestamp 1666464484
transform -1 0 26588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout13_A
timestamp 1666464484
transform -1 0 28704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 29992 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 27876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1666464484
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1666464484
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 1666464484
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_329
timestamp 1666464484
transform 1 0 31372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1666464484
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1666464484
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1666464484
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1666464484
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1666464484
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1666464484
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_329
timestamp 1666464484
transform 1 0 31372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1666464484
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1666464484
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_317
timestamp 1666464484
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_329
timestamp 1666464484
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_305
timestamp 1666464484
transform 1 0 29164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1666464484
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_314
timestamp 1666464484
transform 1 0 29992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_320
timestamp 1666464484
transform 1 0 30544 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_329
timestamp 1666464484
transform 1 0 31372 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_301
timestamp 1666464484
transform 1 0 28796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_315
timestamp 1666464484
transform 1 0 30084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_327
timestamp 1666464484
transform 1 0 31188 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_291
timestamp 1666464484
transform 1 0 27876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_297
timestamp 1666464484
transform 1 0 28428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_303
timestamp 1666464484
transform 1 0 28980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_309
timestamp 1666464484
transform 1 0 29532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_317
timestamp 1666464484
transform 1 0 30268 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_320
timestamp 1666464484
transform 1 0 30544 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_326
timestamp 1666464484
transform 1 0 31096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_330
timestamp 1666464484
transform 1 0 31464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_8
timestamp 1666464484
transform 1 0 1840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1666464484
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_285
timestamp 1666464484
transform 1 0 27324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1666464484
transform 1 0 27600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_294
timestamp 1666464484
transform 1 0 28152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_300
timestamp 1666464484
transform 1 0 28704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666464484
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_313
timestamp 1666464484
transform 1 0 29900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_319
timestamp 1666464484
transform 1 0 30452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_325
timestamp 1666464484
transform 1 0 31004 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_329
timestamp 1666464484
transform 1 0 31372 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1666464484
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_287
timestamp 1666464484
transform 1 0 27508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_290
timestamp 1666464484
transform 1 0 27784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_296
timestamp 1666464484
transform 1 0 28336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_302
timestamp 1666464484
transform 1 0 28888 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_310
timestamp 1666464484
transform 1 0 29624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_313
timestamp 1666464484
transform 1 0 29900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_319
timestamp 1666464484
transform 1 0 30452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_325
timestamp 1666464484
transform 1 0 31004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_329
timestamp 1666464484
transform 1 0 31372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_8
timestamp 1666464484
transform 1 0 1840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1666464484
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_268
timestamp 1666464484
transform 1 0 25760 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_274
timestamp 1666464484
transform 1 0 26312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1666464484
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_286
timestamp 1666464484
transform 1 0 27416 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_296
timestamp 1666464484
transform 1 0 28336 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_302
timestamp 1666464484
transform 1 0 28888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1666464484
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1666464484
transform 1 0 30084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_327
timestamp 1666464484
transform 1 0 31188 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_257
timestamp 1666464484
transform 1 0 24748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_260
timestamp 1666464484
transform 1 0 25024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_266
timestamp 1666464484
transform 1 0 25576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_272
timestamp 1666464484
transform 1 0 26128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1666464484
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_287
timestamp 1666464484
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_290
timestamp 1666464484
transform 1 0 27784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_294
timestamp 1666464484
transform 1 0 28152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_297
timestamp 1666464484
transform 1 0 28428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_303
timestamp 1666464484
transform 1 0 28980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_309
timestamp 1666464484
transform 1 0 29532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_315
timestamp 1666464484
transform 1 0 30084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_321
timestamp 1666464484
transform 1 0 30636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_325
timestamp 1666464484
transform 1 0 31004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_329
timestamp 1666464484
transform 1 0 31372 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_259
timestamp 1666464484
transform 1 0 24932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1666464484
transform 1 0 26036 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_285
timestamp 1666464484
transform 1 0 27324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_291
timestamp 1666464484
transform 1 0 27876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_297
timestamp 1666464484
transform 1 0 28428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1666464484
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_313
timestamp 1666464484
transform 1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_317
timestamp 1666464484
transform 1 0 30268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_320
timestamp 1666464484
transform 1 0 30544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_326
timestamp 1666464484
transform 1 0 31096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_330
timestamp 1666464484
transform 1 0 31464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_8
timestamp 1666464484
transform 1 0 1840 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_20
timestamp 1666464484
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1666464484
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1666464484
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp 1666464484
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_234
timestamp 1666464484
transform 1 0 22632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_238
timestamp 1666464484
transform 1 0 23000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_241
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_247
timestamp 1666464484
transform 1 0 23828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_251
timestamp 1666464484
transform 1 0 24196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_254
timestamp 1666464484
transform 1 0 24472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_260
timestamp 1666464484
transform 1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_264
timestamp 1666464484
transform 1 0 25392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_267
timestamp 1666464484
transform 1 0 25668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_275
timestamp 1666464484
transform 1 0 26404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1666464484
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_285
timestamp 1666464484
transform 1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_291
timestamp 1666464484
transform 1 0 27876 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_297
timestamp 1666464484
transform 1 0 28428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_300
timestamp 1666464484
transform 1 0 28704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_304
timestamp 1666464484
transform 1 0 29072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_307
timestamp 1666464484
transform 1 0 29348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1666464484
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_319
timestamp 1666464484
transform 1 0 30452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_325
timestamp 1666464484
transform 1 0 31004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_329
timestamp 1666464484
transform 1 0 31372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_8
timestamp 1666464484
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1666464484
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_227
timestamp 1666464484
transform 1 0 21988 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_231
timestamp 1666464484
transform 1 0 22356 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1666464484
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_240
timestamp 1666464484
transform 1 0 23184 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1666464484
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_259
timestamp 1666464484
transform 1 0 24932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_273
timestamp 1666464484
transform 1 0 26220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_279
timestamp 1666464484
transform 1 0 26772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_285
timestamp 1666464484
transform 1 0 27324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_288
timestamp 1666464484
transform 1 0 27600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_294
timestamp 1666464484
transform 1 0 28152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_300
timestamp 1666464484
transform 1 0 28704 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1666464484
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_315
timestamp 1666464484
transform 1 0 30084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1666464484
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_324
timestamp 1666464484
transform 1 0 30912 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_330
timestamp 1666464484
transform 1 0 31464 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_213
timestamp 1666464484
transform 1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1666464484
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_229
timestamp 1666464484
transform 1 0 22172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_235
timestamp 1666464484
transform 1 0 22724 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_241
timestamp 1666464484
transform 1 0 23276 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_259
timestamp 1666464484
transform 1 0 24932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_265
timestamp 1666464484
transform 1 0 25484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_271
timestamp 1666464484
transform 1 0 26036 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1666464484
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_287
timestamp 1666464484
transform 1 0 27508 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_295
timestamp 1666464484
transform 1 0 28244 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_298
timestamp 1666464484
transform 1 0 28520 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_302
timestamp 1666464484
transform 1 0 28888 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_305
timestamp 1666464484
transform 1 0 29164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_311
timestamp 1666464484
transform 1 0 29716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_317
timestamp 1666464484
transform 1 0 30268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_325
timestamp 1666464484
transform 1 0 31004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_211
timestamp 1666464484
transform 1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1666464484
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_225
timestamp 1666464484
transform 1 0 21804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_232
timestamp 1666464484
transform 1 0 22448 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_238
timestamp 1666464484
transform 1 0 23000 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_244
timestamp 1666464484
transform 1 0 23552 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1666464484
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_257
timestamp 1666464484
transform 1 0 24748 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_267
timestamp 1666464484
transform 1 0 25668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_275
timestamp 1666464484
transform 1 0 26404 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_278
timestamp 1666464484
transform 1 0 26680 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_284
timestamp 1666464484
transform 1 0 27232 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_287
timestamp 1666464484
transform 1 0 27508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_293
timestamp 1666464484
transform 1 0 28060 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_299
timestamp 1666464484
transform 1 0 28612 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_302
timestamp 1666464484
transform 1 0 28888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_313
timestamp 1666464484
transform 1 0 29900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_319
timestamp 1666464484
transform 1 0 30452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_325
timestamp 1666464484
transform 1 0 31004 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_329
timestamp 1666464484
transform 1 0 31372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_8
timestamp 1666464484
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1666464484
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1666464484
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1666464484
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1666464484
transform 1 0 19412 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_202
timestamp 1666464484
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1666464484
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_216
timestamp 1666464484
transform 1 0 20976 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1666464484
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1666464484
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1666464484
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_250
timestamp 1666464484
transform 1 0 24104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_256
timestamp 1666464484
transform 1 0 24656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_262
timestamp 1666464484
transform 1 0 25208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_265
timestamp 1666464484
transform 1 0 25484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1666464484
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_285
timestamp 1666464484
transform 1 0 27324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_291
timestamp 1666464484
transform 1 0 27876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_297
timestamp 1666464484
transform 1 0 28428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1666464484
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_309
timestamp 1666464484
transform 1 0 29532 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_315
timestamp 1666464484
transform 1 0 30084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_321
timestamp 1666464484
transform 1 0 30636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_327
timestamp 1666464484
transform 1 0 31188 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1666464484
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1666464484
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1666464484
transform 1 0 19964 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1666464484
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1666464484
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_231
timestamp 1666464484
transform 1 0 22356 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1666464484
transform 1 0 23000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_257
timestamp 1666464484
transform 1 0 24748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_263
timestamp 1666464484
transform 1 0 25300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1666464484
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1666464484
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_281
timestamp 1666464484
transform 1 0 26956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_287
timestamp 1666464484
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_299
timestamp 1666464484
transform 1 0 28612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1666464484
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_313
timestamp 1666464484
transform 1 0 29900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_319
timestamp 1666464484
transform 1 0 30452 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_325
timestamp 1666464484
transform 1 0 31004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_329
timestamp 1666464484
transform 1 0 31372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1666464484
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1666464484
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1666464484
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_177
timestamp 1666464484
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1666464484
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1666464484
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1666464484
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_202
timestamp 1666464484
transform 1 0 19688 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1666464484
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1666464484
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_232
timestamp 1666464484
transform 1 0 22448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1666464484
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_246
timestamp 1666464484
transform 1 0 23736 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_253
timestamp 1666464484
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1666464484
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_264
timestamp 1666464484
transform 1 0 25392 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_268
timestamp 1666464484
transform 1 0 25760 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1666464484
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_285
timestamp 1666464484
transform 1 0 27324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_291
timestamp 1666464484
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_297
timestamp 1666464484
transform 1 0 28428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_303
timestamp 1666464484
transform 1 0 28980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_309
timestamp 1666464484
transform 1 0 29532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_315
timestamp 1666464484
transform 1 0 30084 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_321
timestamp 1666464484
transform 1 0 30636 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_325
timestamp 1666464484
transform 1 0 31004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_329
timestamp 1666464484
transform 1 0 31372 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_171
timestamp 1666464484
transform 1 0 16836 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1666464484
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1666464484
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1666464484
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_232
timestamp 1666464484
transform 1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_240
timestamp 1666464484
transform 1 0 23184 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1666464484
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1666464484
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1666464484
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_279
timestamp 1666464484
transform 1 0 26772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_285
timestamp 1666464484
transform 1 0 27324 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1666464484
transform 1 0 27876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_297
timestamp 1666464484
transform 1 0 28428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1666464484
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_313
timestamp 1666464484
transform 1 0 29900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_319
timestamp 1666464484
transform 1 0 30452 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_325
timestamp 1666464484
transform 1 0 31004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_329
timestamp 1666464484
transform 1 0 31372 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1666464484
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_182
timestamp 1666464484
transform 1 0 17848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1666464484
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_198
timestamp 1666464484
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1666464484
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1666464484
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1666464484
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_258
timestamp 1666464484
transform 1 0 24840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_263
timestamp 1666464484
transform 1 0 25300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_270
timestamp 1666464484
transform 1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1666464484
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1666464484
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_292
timestamp 1666464484
transform 1 0 27968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_298
timestamp 1666464484
transform 1 0 28520 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_304
timestamp 1666464484
transform 1 0 29072 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_310
timestamp 1666464484
transform 1 0 29624 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 1666464484
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_322
timestamp 1666464484
transform 1 0 30728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_155
timestamp 1666464484
transform 1 0 15364 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1666464484
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_169
timestamp 1666464484
transform 1 0 16652 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1666464484
transform 1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_183
timestamp 1666464484
transform 1 0 17940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1666464484
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 23460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1666464484
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1666464484
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_263
timestamp 1666464484
transform 1 0 25300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1666464484
transform 1 0 26036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_279
timestamp 1666464484
transform 1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1666464484
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_293
timestamp 1666464484
transform 1 0 28060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_300
timestamp 1666464484
transform 1 0 28704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1666464484
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_315
timestamp 1666464484
transform 1 0 30084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_322
timestamp 1666464484
transform 1 0 30728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_329
timestamp 1666464484
transform 1 0 31372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_8
timestamp 1666464484
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_20
timestamp 1666464484
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_32
timestamp 1666464484
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1666464484
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1666464484
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_139
timestamp 1666464484
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1666464484
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1666464484
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_152
timestamp 1666464484
transform 1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1666464484
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1666464484
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1666464484
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_189
timestamp 1666464484
transform 1 0 18492 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_213
timestamp 1666464484
transform 1 0 20700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1666464484
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1666464484
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1666464484
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_267
timestamp 1666464484
transform 1 0 25668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1666464484
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1666464484
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_300
timestamp 1666464484
transform 1 0 28704 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_307
timestamp 1666464484
transform 1 0 29348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_311
timestamp 1666464484
transform 1 0 29716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_315
timestamp 1666464484
transform 1 0 30084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_322
timestamp 1666464484
transform 1 0 30728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_329
timestamp 1666464484
transform 1 0 31372 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_129
timestamp 1666464484
transform 1 0 12972 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_132
timestamp 1666464484
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1666464484
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1666464484
transform 1 0 14720 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_155
timestamp 1666464484
transform 1 0 15364 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1666464484
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1666464484
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_183
timestamp 1666464484
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1666464484
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1666464484
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_244
timestamp 1666464484
transform 1 0 23552 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1666464484
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1666464484
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_273
timestamp 1666464484
transform 1 0 26220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_282
timestamp 1666464484
transform 1 0 27048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_290
timestamp 1666464484
transform 1 0 27784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_297
timestamp 1666464484
transform 1 0 28428 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1666464484
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1666464484
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_318
timestamp 1666464484
transform 1 0 30360 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_322
timestamp 1666464484
transform 1 0 30728 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_329
timestamp 1666464484
transform 1 0 31372 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1666464484
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_120
timestamp 1666464484
transform 1 0 12144 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_130
timestamp 1666464484
transform 1 0 13064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_141
timestamp 1666464484
transform 1 0 14076 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_148
timestamp 1666464484
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_156
timestamp 1666464484
transform 1 0 15456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_173
timestamp 1666464484
transform 1 0 17020 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1666464484
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1666464484
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1666464484
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_247
timestamp 1666464484
transform 1 0 23828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_271
timestamp 1666464484
transform 1 0 26036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1666464484
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_288
timestamp 1666464484
transform 1 0 27600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1666464484
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_304
timestamp 1666464484
transform 1 0 29072 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_311
timestamp 1666464484
transform 1 0 29716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1666464484
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_325
timestamp 1666464484
transform 1 0 31004 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_8
timestamp 1666464484
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1666464484
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_112
timestamp 1666464484
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 1666464484
transform 1 0 11960 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1666464484
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1666464484
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1666464484
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_150
timestamp 1666464484
transform 1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1666464484
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1666464484
transform 1 0 16744 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1666464484
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1666464484
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_243
timestamp 1666464484
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1666464484
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_275
timestamp 1666464484
transform 1 0 26404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_285
timestamp 1666464484
transform 1 0 27324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_294
timestamp 1666464484
transform 1 0 28152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1666464484
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666464484
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_315
timestamp 1666464484
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_323
timestamp 1666464484
transform 1 0 30820 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_329
timestamp 1666464484
transform 1 0 31372 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_101
timestamp 1666464484
transform 1 0 10396 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_104
timestamp 1666464484
transform 1 0 10672 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1666464484
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_128
timestamp 1666464484
transform 1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1666464484
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_143
timestamp 1666464484
transform 1 0 14260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1666464484
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_175
timestamp 1666464484
transform 1 0 17204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_188
timestamp 1666464484
transform 1 0 18400 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_212
timestamp 1666464484
transform 1 0 20608 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1666464484
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1666464484
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_271
timestamp 1666464484
transform 1 0 26036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1666464484
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 1666464484
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1666464484
transform 1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_307
timestamp 1666464484
transform 1 0 29348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1666464484
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_323
timestamp 1666464484
transform 1 0 30820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_8
timestamp 1666464484
transform 1 0 1840 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_20
timestamp 1666464484
transform 1 0 2944 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1666464484
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_103
timestamp 1666464484
transform 1 0 10580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_116
timestamp 1666464484
transform 1 0 11776 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1666464484
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1666464484
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1666464484
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1666464484
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_158
timestamp 1666464484
transform 1 0 15640 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1666464484
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1666464484
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1666464484
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_243
timestamp 1666464484
transform 1 0 23460 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1666464484
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_263
timestamp 1666464484
transform 1 0 25300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_274
timestamp 1666464484
transform 1 0 26312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_285
timestamp 1666464484
transform 1 0 27324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1666464484
transform 1 0 28244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1666464484
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_316
timestamp 1666464484
transform 1 0 30176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_324
timestamp 1666464484
transform 1 0 30912 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_330
timestamp 1666464484
transform 1 0 31464 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_91
timestamp 1666464484
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1666464484
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1666464484
transform 1 0 10580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1666464484
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1666464484
transform 1 0 11960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1666464484
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1666464484
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1666464484
transform 1 0 14352 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_154
timestamp 1666464484
transform 1 0 15272 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_175
timestamp 1666464484
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_189
timestamp 1666464484
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1666464484
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1666464484
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_248
timestamp 1666464484
transform 1 0 23920 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_272
timestamp 1666464484
transform 1 0 26128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1666464484
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1666464484
transform 1 0 27784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_301
timestamp 1666464484
transform 1 0 28796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_310
timestamp 1666464484
transform 1 0 29624 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_319
timestamp 1666464484
transform 1 0 30452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_328
timestamp 1666464484
transform 1 0 31280 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1666464484
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1666464484
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_96
timestamp 1666464484
transform 1 0 9936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_102
timestamp 1666464484
transform 1 0 10488 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_116
timestamp 1666464484
transform 1 0 11776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1666464484
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1666464484
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1666464484
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1666464484
transform 1 0 14812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1666464484
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1666464484
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_207
timestamp 1666464484
transform 1 0 20148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_232
timestamp 1666464484
transform 1 0 22448 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_263
timestamp 1666464484
transform 1 0 25300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_274
timestamp 1666464484
transform 1 0 26312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1666464484
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_296
timestamp 1666464484
transform 1 0 28336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1666464484
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_317
timestamp 1666464484
transform 1 0 30268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_326
timestamp 1666464484
transform 1 0 31096 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_330
timestamp 1666464484
transform 1 0 31464 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1666464484
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1666464484
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1666464484
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1666464484
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_77
timestamp 1666464484
transform 1 0 8188 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_80
timestamp 1666464484
transform 1 0 8464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_86
timestamp 1666464484
transform 1 0 9016 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_92
timestamp 1666464484
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 1666464484
transform 1 0 10120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_104
timestamp 1666464484
transform 1 0 10672 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1666464484
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1666464484
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1666464484
transform 1 0 12420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1666464484
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_138
timestamp 1666464484
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1666464484
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_156
timestamp 1666464484
transform 1 0 15456 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1666464484
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_175
timestamp 1666464484
transform 1 0 17204 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_183
timestamp 1666464484
transform 1 0 17940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_197
timestamp 1666464484
transform 1 0 19228 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1666464484
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1666464484
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_271
timestamp 1666464484
transform 1 0 26036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1666464484
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_290
timestamp 1666464484
transform 1 0 27784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1666464484
transform 1 0 28796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_312
timestamp 1666464484
transform 1 0 29808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_322
timestamp 1666464484
transform 1 0 30728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_329
timestamp 1666464484
transform 1 0 31372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_8
timestamp 1666464484
transform 1 0 1840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1666464484
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_70
timestamp 1666464484
transform 1 0 7544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_76
timestamp 1666464484
transform 1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1666464484
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1666464484
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_103
timestamp 1666464484
transform 1 0 10580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1666464484
transform 1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1666464484
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_130
timestamp 1666464484
transform 1 0 13064 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1666464484
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_147
timestamp 1666464484
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_162
timestamp 1666464484
transform 1 0 16008 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1666464484
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 1666464484
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1666464484
transform 1 0 19596 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_228
timestamp 1666464484
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_241
timestamp 1666464484
transform 1 0 23276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_275
timestamp 1666464484
transform 1 0 26404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_287
timestamp 1666464484
transform 1 0 27508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_298
timestamp 1666464484
transform 1 0 28520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1666464484
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_318
timestamp 1666464484
transform 1 0 30360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_328
timestamp 1666464484
transform 1 0 31280 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_61
timestamp 1666464484
transform 1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_67
timestamp 1666464484
transform 1 0 7268 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_73
timestamp 1666464484
transform 1 0 7820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1666464484
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1666464484
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_91
timestamp 1666464484
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_97
timestamp 1666464484
transform 1 0 10028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1666464484
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1666464484
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1666464484
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_121
timestamp 1666464484
transform 1 0 12236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_129
timestamp 1666464484
transform 1 0 12972 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1666464484
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_155
timestamp 1666464484
transform 1 0 15364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1666464484
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_185
timestamp 1666464484
transform 1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1666464484
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1666464484
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1666464484
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_251
timestamp 1666464484
transform 1 0 24196 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_291
timestamp 1666464484
transform 1 0 27876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1666464484
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_314
timestamp 1666464484
transform 1 0 29992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_325
timestamp 1666464484
transform 1 0 31004 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1666464484
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_64
timestamp 1666464484
transform 1 0 6992 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1666464484
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_76
timestamp 1666464484
transform 1 0 8096 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1666464484
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1666464484
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp 1666464484
transform 1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_98
timestamp 1666464484
transform 1 0 10120 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1666464484
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1666464484
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1666464484
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1666464484
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_160
timestamp 1666464484
transform 1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_171
timestamp 1666464484
transform 1 0 16836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_182
timestamp 1666464484
transform 1 0 17848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1666464484
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_202
timestamp 1666464484
transform 1 0 19688 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_229
timestamp 1666464484
transform 1 0 22172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1666464484
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_276
timestamp 1666464484
transform 1 0 26496 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666464484
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666464484
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_318
timestamp 1666464484
transform 1 0 30360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_329
timestamp 1666464484
transform 1 0 31372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1666464484
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_44
timestamp 1666464484
transform 1 0 5152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_48
timestamp 1666464484
transform 1 0 5520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1666464484
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1666464484
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_64
timestamp 1666464484
transform 1 0 6992 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_70
timestamp 1666464484
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_76
timestamp 1666464484
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1666464484
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_88
timestamp 1666464484
transform 1 0 9200 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_95
timestamp 1666464484
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_102
timestamp 1666464484
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1666464484
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1666464484
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_126
timestamp 1666464484
transform 1 0 12696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1666464484
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1666464484
transform 1 0 14352 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1666464484
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1666464484
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1666464484
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_185
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_197
timestamp 1666464484
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1666464484
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_248
timestamp 1666464484
transform 1 0 23920 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1666464484
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1666464484
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_315
timestamp 1666464484
transform 1 0 30084 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_326
timestamp 1666464484
transform 1 0 31096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_330
timestamp 1666464484
transform 1 0 31464 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_46
timestamp 1666464484
transform 1 0 5336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_52
timestamp 1666464484
transform 1 0 5888 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1666464484
transform 1 0 6440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_64
timestamp 1666464484
transform 1 0 6992 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1666464484
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_76
timestamp 1666464484
transform 1 0 8096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1666464484
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_89
timestamp 1666464484
transform 1 0 9292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1666464484
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1666464484
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_111
timestamp 1666464484
transform 1 0 11316 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_120
timestamp 1666464484
transform 1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1666464484
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1666464484
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1666464484
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_159
timestamp 1666464484
transform 1 0 15732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1666464484
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_182
timestamp 1666464484
transform 1 0 17848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1666464484
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1666464484
transform 1 0 19596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1666464484
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666464484
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666464484
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_319
timestamp 1666464484
transform 1 0 30452 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_329
timestamp 1666464484
transform 1 0 31372 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1666464484
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1666464484
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_32
timestamp 1666464484
transform 1 0 4048 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_42
timestamp 1666464484
transform 1 0 4968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_48
timestamp 1666464484
transform 1 0 5520 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1666464484
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_61
timestamp 1666464484
transform 1 0 6716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_64
timestamp 1666464484
transform 1 0 6992 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_70
timestamp 1666464484
transform 1 0 7544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_76
timestamp 1666464484
transform 1 0 8096 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1666464484
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_88
timestamp 1666464484
transform 1 0 9200 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_95
timestamp 1666464484
transform 1 0 9844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_102
timestamp 1666464484
transform 1 0 10488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1666464484
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1666464484
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1666464484
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1666464484
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_155
timestamp 1666464484
transform 1 0 15364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1666464484
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1666464484
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_195
timestamp 1666464484
transform 1 0 19044 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_248
timestamp 1666464484
transform 1 0 23920 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_256
timestamp 1666464484
transform 1 0 24656 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1666464484
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_303
timestamp 1666464484
transform 1 0 28980 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_315
timestamp 1666464484
transform 1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_327
timestamp 1666464484
transform 1 0 31188 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_34
timestamp 1666464484
transform 1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_40
timestamp 1666464484
transform 1 0 4784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_46
timestamp 1666464484
transform 1 0 5336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_52
timestamp 1666464484
transform 1 0 5888 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1666464484
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_64
timestamp 1666464484
transform 1 0 6992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1666464484
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_76
timestamp 1666464484
transform 1 0 8096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1666464484
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1666464484
transform 1 0 9476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_95
timestamp 1666464484
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_102
timestamp 1666464484
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1666464484
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1666464484
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1666464484
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1666464484
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_148
timestamp 1666464484
transform 1 0 14720 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1666464484
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_170
timestamp 1666464484
transform 1 0 16744 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_182
timestamp 1666464484
transform 1 0 17848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1666464484
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_276
timestamp 1666464484
transform 1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_296
timestamp 1666464484
transform 1 0 28336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1666464484
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_319
timestamp 1666464484
transform 1 0 30452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_329
timestamp 1666464484
transform 1 0 31372 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_33
timestamp 1666464484
transform 1 0 4140 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_36
timestamp 1666464484
transform 1 0 4416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_42
timestamp 1666464484
transform 1 0 4968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_48
timestamp 1666464484
transform 1 0 5520 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1666464484
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_63
timestamp 1666464484
transform 1 0 6900 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_66
timestamp 1666464484
transform 1 0 7176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_72
timestamp 1666464484
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_78
timestamp 1666464484
transform 1 0 8280 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1666464484
transform 1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1666464484
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_96
timestamp 1666464484
transform 1 0 9936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_103
timestamp 1666464484
transform 1 0 10580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1666464484
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1666464484
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_127
timestamp 1666464484
transform 1 0 12788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_136
timestamp 1666464484
transform 1 0 13616 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1666464484
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1666464484
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1666464484
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_173
timestamp 1666464484
transform 1 0 17020 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1666464484
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_233
timestamp 1666464484
transform 1 0 22540 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_250
timestamp 1666464484
transform 1 0 24104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1666464484
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1666464484
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1666464484
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_318
timestamp 1666464484
transform 1 0 30360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_329
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_8
timestamp 1666464484
transform 1 0 1840 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_20
timestamp 1666464484
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_34
timestamp 1666464484
transform 1 0 4232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_40
timestamp 1666464484
transform 1 0 4784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_46
timestamp 1666464484
transform 1 0 5336 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_52
timestamp 1666464484
transform 1 0 5888 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_58
timestamp 1666464484
transform 1 0 6440 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_64
timestamp 1666464484
transform 1 0 6992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_70
timestamp 1666464484
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_76
timestamp 1666464484
transform 1 0 8096 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1666464484
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_89
timestamp 1666464484
transform 1 0 9292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_95
timestamp 1666464484
transform 1 0 9844 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_101
timestamp 1666464484
transform 1 0 10396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1666464484
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_114
timestamp 1666464484
transform 1 0 11592 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_129
timestamp 1666464484
transform 1 0 12972 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1666464484
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1666464484
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_160
timestamp 1666464484
transform 1 0 15824 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1666464484
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_182
timestamp 1666464484
transform 1 0 17848 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1666464484
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_203
timestamp 1666464484
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_212
timestamp 1666464484
transform 1 0 20608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1666464484
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_275
timestamp 1666464484
transform 1 0 26404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_292
timestamp 1666464484
transform 1 0 27968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1666464484
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_319
timestamp 1666464484
transform 1 0 30452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_329
timestamp 1666464484
transform 1 0 31372 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1666464484
transform 1 0 1840 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_20
timestamp 1666464484
transform 1 0 2944 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_32
timestamp 1666464484
transform 1 0 4048 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_36
timestamp 1666464484
transform 1 0 4416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_42
timestamp 1666464484
transform 1 0 4968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_48
timestamp 1666464484
transform 1 0 5520 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1666464484
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1666464484
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_68
timestamp 1666464484
transform 1 0 7360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_74
timestamp 1666464484
transform 1 0 7912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_80
timestamp 1666464484
transform 1 0 8464 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_86
timestamp 1666464484
transform 1 0 9016 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_92
timestamp 1666464484
transform 1 0 9568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_98
timestamp 1666464484
transform 1 0 10120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_104
timestamp 1666464484
transform 1 0 10672 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1666464484
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1666464484
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1666464484
transform 1 0 12420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_130
timestamp 1666464484
transform 1 0 13064 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_138
timestamp 1666464484
transform 1 0 13800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_147
timestamp 1666464484
transform 1 0 14628 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_156
timestamp 1666464484
transform 1 0 15456 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1666464484
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_182
timestamp 1666464484
transform 1 0 17848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1666464484
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_263
timestamp 1666464484
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1666464484
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_305
timestamp 1666464484
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_317
timestamp 1666464484
transform 1 0 30268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_329
timestamp 1666464484
transform 1 0 31372 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1666464484
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1666464484
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_46
timestamp 1666464484
transform 1 0 5336 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_52
timestamp 1666464484
transform 1 0 5888 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_58
timestamp 1666464484
transform 1 0 6440 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_64
timestamp 1666464484
transform 1 0 6992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_70
timestamp 1666464484
transform 1 0 7544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_76
timestamp 1666464484
transform 1 0 8096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1666464484
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_93
timestamp 1666464484
transform 1 0 9660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1666464484
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_105
timestamp 1666464484
transform 1 0 10764 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_111
timestamp 1666464484
transform 1 0 11316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_117
timestamp 1666464484
transform 1 0 11868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1666464484
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_131
timestamp 1666464484
transform 1 0 13156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1666464484
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1666464484
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_162
timestamp 1666464484
transform 1 0 16008 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1666464484
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1666464484
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1666464484
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_226
timestamp 1666464484
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1666464484
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_276
timestamp 1666464484
transform 1 0 26496 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_300
timestamp 1666464484
transform 1 0 28704 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1666464484
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_319
timestamp 1666464484
transform 1 0 30452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_329
timestamp 1666464484
transform 1 0 31372 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_42
timestamp 1666464484
transform 1 0 4968 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_48
timestamp 1666464484
transform 1 0 5520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1666464484
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1666464484
transform 1 0 6808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_68
timestamp 1666464484
transform 1 0 7360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_74
timestamp 1666464484
transform 1 0 7912 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1666464484
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_86
timestamp 1666464484
transform 1 0 9016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_92
timestamp 1666464484
transform 1 0 9568 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_98
timestamp 1666464484
transform 1 0 10120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_104
timestamp 1666464484
transform 1 0 10672 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1666464484
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_117
timestamp 1666464484
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_120
timestamp 1666464484
transform 1 0 12144 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1666464484
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_133
timestamp 1666464484
transform 1 0 13340 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_140
timestamp 1666464484
transform 1 0 13984 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_148
timestamp 1666464484
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_157
timestamp 1666464484
transform 1 0 15548 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1666464484
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1666464484
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_188
timestamp 1666464484
transform 1 0 18400 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_199
timestamp 1666464484
transform 1 0 19412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_210
timestamp 1666464484
transform 1 0 20424 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_235
timestamp 1666464484
transform 1 0 22724 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_262
timestamp 1666464484
transform 1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1666464484
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_291
timestamp 1666464484
transform 1 0 27876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_303
timestamp 1666464484
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_315
timestamp 1666464484
transform 1 0 30084 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_326
timestamp 1666464484
transform 1 0 31096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_330
timestamp 1666464484
transform 1 0 31464 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_8
timestamp 1666464484
transform 1 0 1840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1666464484
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_46
timestamp 1666464484
transform 1 0 5336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_52
timestamp 1666464484
transform 1 0 5888 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1666464484
transform 1 0 6440 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_64
timestamp 1666464484
transform 1 0 6992 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_70
timestamp 1666464484
transform 1 0 7544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_76
timestamp 1666464484
transform 1 0 8096 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1666464484
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1666464484
transform 1 0 9292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_95
timestamp 1666464484
transform 1 0 9844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1666464484
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1666464484
transform 1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_113
timestamp 1666464484
transform 1 0 11500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_119
timestamp 1666464484
transform 1 0 12052 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1666464484
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_131
timestamp 1666464484
transform 1 0 13156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1666464484
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_150
timestamp 1666464484
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_157
timestamp 1666464484
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_166
timestamp 1666464484
transform 1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1666464484
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_184
timestamp 1666464484
transform 1 0 18032 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1666464484
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_203
timestamp 1666464484
transform 1 0 19780 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_214
timestamp 1666464484
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_226
timestamp 1666464484
transform 1 0 21896 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1666464484
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_276
timestamp 1666464484
transform 1 0 26496 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_288
timestamp 1666464484
transform 1 0 27600 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_300
timestamp 1666464484
transform 1 0 28704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1666464484
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_318
timestamp 1666464484
transform 1 0 30360 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_329
timestamp 1666464484
transform 1 0 31372 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_45
timestamp 1666464484
transform 1 0 5244 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_48
timestamp 1666464484
transform 1 0 5520 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1666464484
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_62
timestamp 1666464484
transform 1 0 6808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_68
timestamp 1666464484
transform 1 0 7360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_74
timestamp 1666464484
transform 1 0 7912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_80
timestamp 1666464484
transform 1 0 8464 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_86
timestamp 1666464484
transform 1 0 9016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_92
timestamp 1666464484
transform 1 0 9568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_98
timestamp 1666464484
transform 1 0 10120 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_104
timestamp 1666464484
transform 1 0 10672 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1666464484
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_121
timestamp 1666464484
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_127
timestamp 1666464484
transform 1 0 12788 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_133
timestamp 1666464484
transform 1 0 13340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_139
timestamp 1666464484
transform 1 0 13892 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_145
timestamp 1666464484
transform 1 0 14444 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_152
timestamp 1666464484
transform 1 0 15088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_159
timestamp 1666464484
transform 1 0 15732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1666464484
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_175
timestamp 1666464484
transform 1 0 17204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_190
timestamp 1666464484
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_200
timestamp 1666464484
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1666464484
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1666464484
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1666464484
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1666464484
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_291
timestamp 1666464484
transform 1 0 27876 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_302
timestamp 1666464484
transform 1 0 28888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_313
timestamp 1666464484
transform 1 0 29900 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_323
timestamp 1666464484
transform 1 0 30820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1666464484
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1666464484
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_49
timestamp 1666464484
transform 1 0 5612 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_52
timestamp 1666464484
transform 1 0 5888 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_58
timestamp 1666464484
transform 1 0 6440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_64
timestamp 1666464484
transform 1 0 6992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_70
timestamp 1666464484
transform 1 0 7544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_76
timestamp 1666464484
transform 1 0 8096 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1666464484
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_90
timestamp 1666464484
transform 1 0 9384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_96
timestamp 1666464484
transform 1 0 9936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1666464484
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_108
timestamp 1666464484
transform 1 0 11040 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1666464484
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1666464484
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1666464484
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_132
timestamp 1666464484
transform 1 0 13248 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1666464484
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_149
timestamp 1666464484
transform 1 0 14812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_155
timestamp 1666464484
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_162
timestamp 1666464484
transform 1 0 16008 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_169
timestamp 1666464484
transform 1 0 16652 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_185
timestamp 1666464484
transform 1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_220
timestamp 1666464484
transform 1 0 21344 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_231
timestamp 1666464484
transform 1 0 22356 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1666464484
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_264
timestamp 1666464484
transform 1 0 25392 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_276
timestamp 1666464484
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1666464484
transform 1 0 27600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_299
timestamp 1666464484
transform 1 0 28612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1666464484
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_317
timestamp 1666464484
transform 1 0 30268 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_326
timestamp 1666464484
transform 1 0 31096 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_330
timestamp 1666464484
transform 1 0 31464 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_62
timestamp 1666464484
transform 1 0 6808 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_68
timestamp 1666464484
transform 1 0 7360 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_74
timestamp 1666464484
transform 1 0 7912 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_80
timestamp 1666464484
transform 1 0 8464 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1666464484
transform 1 0 9016 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_92
timestamp 1666464484
transform 1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_98
timestamp 1666464484
transform 1 0 10120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_104
timestamp 1666464484
transform 1 0 10672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1666464484
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1666464484
transform 1 0 11960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1666464484
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_130
timestamp 1666464484
transform 1 0 13064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1666464484
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_142
timestamp 1666464484
transform 1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_148
timestamp 1666464484
transform 1 0 14720 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_154
timestamp 1666464484
transform 1 0 15272 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_160
timestamp 1666464484
transform 1 0 15824 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_178
timestamp 1666464484
transform 1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_186
timestamp 1666464484
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_194
timestamp 1666464484
transform 1 0 18952 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_203
timestamp 1666464484
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_212
timestamp 1666464484
transform 1 0 20608 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1666464484
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_229
timestamp 1666464484
transform 1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_240
timestamp 1666464484
transform 1 0 23184 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_254
timestamp 1666464484
transform 1 0 24472 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_266
timestamp 1666464484
transform 1 0 25576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1666464484
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_290
timestamp 1666464484
transform 1 0 27784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1666464484
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_311
timestamp 1666464484
transform 1 0 29716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_320
timestamp 1666464484
transform 1 0 30544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_329
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_58
timestamp 1666464484
transform 1 0 6440 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_64
timestamp 1666464484
transform 1 0 6992 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_70
timestamp 1666464484
transform 1 0 7544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_76
timestamp 1666464484
transform 1 0 8096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1666464484
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_90
timestamp 1666464484
transform 1 0 9384 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_96
timestamp 1666464484
transform 1 0 9936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_102
timestamp 1666464484
transform 1 0 10488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_108
timestamp 1666464484
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_114
timestamp 1666464484
transform 1 0 11592 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_120
timestamp 1666464484
transform 1 0 12144 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_126
timestamp 1666464484
transform 1 0 12696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_132
timestamp 1666464484
transform 1 0 13248 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1666464484
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_147
timestamp 1666464484
transform 1 0 14628 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_157
timestamp 1666464484
transform 1 0 15548 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_160
timestamp 1666464484
transform 1 0 15824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_166
timestamp 1666464484
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_172
timestamp 1666464484
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1666464484
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_186
timestamp 1666464484
transform 1 0 18216 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_205
timestamp 1666464484
transform 1 0 19964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_214
timestamp 1666464484
transform 1 0 20792 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_223
timestamp 1666464484
transform 1 0 21620 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_229
timestamp 1666464484
transform 1 0 22172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1666464484
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1666464484
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_263
timestamp 1666464484
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_274
timestamp 1666464484
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1666464484
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_296
timestamp 1666464484
transform 1 0 28336 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1666464484
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_316
timestamp 1666464484
transform 1 0 30176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_324
timestamp 1666464484
transform 1 0 30912 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_330
timestamp 1666464484
transform 1 0 31464 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1666464484
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1666464484
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1666464484
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1666464484
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_65
timestamp 1666464484
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_68
timestamp 1666464484
transform 1 0 7360 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_74
timestamp 1666464484
transform 1 0 7912 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_80
timestamp 1666464484
transform 1 0 8464 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_86
timestamp 1666464484
transform 1 0 9016 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1666464484
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_98
timestamp 1666464484
transform 1 0 10120 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_104
timestamp 1666464484
transform 1 0 10672 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1666464484
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_119
timestamp 1666464484
transform 1 0 12052 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1666464484
transform 1 0 12328 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_128
timestamp 1666464484
transform 1 0 12880 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_134
timestamp 1666464484
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_140
timestamp 1666464484
transform 1 0 13984 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_146
timestamp 1666464484
transform 1 0 14536 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_155
timestamp 1666464484
transform 1 0 15364 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_163
timestamp 1666464484
transform 1 0 16100 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1666464484
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_177
timestamp 1666464484
transform 1 0 17388 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_183
timestamp 1666464484
transform 1 0 17940 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_190
timestamp 1666464484
transform 1 0 18584 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_197
timestamp 1666464484
transform 1 0 19228 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1666464484
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1666464484
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_232
timestamp 1666464484
transform 1 0 22448 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1666464484
transform 1 0 23460 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_254
timestamp 1666464484
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_265
timestamp 1666464484
transform 1 0 25484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1666464484
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_290
timestamp 1666464484
transform 1 0 27784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_300
timestamp 1666464484
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_309
timestamp 1666464484
transform 1 0 29532 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_317
timestamp 1666464484
transform 1 0 30268 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_329
timestamp 1666464484
transform 1 0 31372 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_8
timestamp 1666464484
transform 1 0 1840 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1666464484
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_70
timestamp 1666464484
transform 1 0 7544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_76
timestamp 1666464484
transform 1 0 8096 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1666464484
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_90
timestamp 1666464484
transform 1 0 9384 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_96
timestamp 1666464484
transform 1 0 9936 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_102
timestamp 1666464484
transform 1 0 10488 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_108
timestamp 1666464484
transform 1 0 11040 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_114
timestamp 1666464484
transform 1 0 11592 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_120
timestamp 1666464484
transform 1 0 12144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_126
timestamp 1666464484
transform 1 0 12696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_132
timestamp 1666464484
transform 1 0 13248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1666464484
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_149
timestamp 1666464484
transform 1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_155
timestamp 1666464484
transform 1 0 15364 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_161
timestamp 1666464484
transform 1 0 15916 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_169
timestamp 1666464484
transform 1 0 16652 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_175
timestamp 1666464484
transform 1 0 17204 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_181
timestamp 1666464484
transform 1 0 17756 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_187
timestamp 1666464484
transform 1 0 18308 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1666464484
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_205
timestamp 1666464484
transform 1 0 19964 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_213
timestamp 1666464484
transform 1 0 20700 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_230
timestamp 1666464484
transform 1 0 22264 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_239
timestamp 1666464484
transform 1 0 23092 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1666464484
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_262
timestamp 1666464484
transform 1 0 25208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_273
timestamp 1666464484
transform 1 0 26220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_283
timestamp 1666464484
transform 1 0 27140 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_292
timestamp 1666464484
transform 1 0 27968 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_314
timestamp 1666464484
transform 1 0 29992 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_321
timestamp 1666464484
transform 1 0 30636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_329
timestamp 1666464484
transform 1 0 31372 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_74
timestamp 1666464484
transform 1 0 7912 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_80
timestamp 1666464484
transform 1 0 8464 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_86
timestamp 1666464484
transform 1 0 9016 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_92
timestamp 1666464484
transform 1 0 9568 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_98
timestamp 1666464484
transform 1 0 10120 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_104
timestamp 1666464484
transform 1 0 10672 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1666464484
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_118
timestamp 1666464484
transform 1 0 11960 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_124
timestamp 1666464484
transform 1 0 12512 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_130
timestamp 1666464484
transform 1 0 13064 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_136
timestamp 1666464484
transform 1 0 13616 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_142
timestamp 1666464484
transform 1 0 14168 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_148
timestamp 1666464484
transform 1 0 14720 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1666464484
transform 1 0 15272 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_160
timestamp 1666464484
transform 1 0 15824 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1666464484
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_173
timestamp 1666464484
transform 1 0 17020 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_179
timestamp 1666464484
transform 1 0 17572 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_185
timestamp 1666464484
transform 1 0 18124 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_191
timestamp 1666464484
transform 1 0 18676 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_197
timestamp 1666464484
transform 1 0 19228 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_203
timestamp 1666464484
transform 1 0 19780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_207
timestamp 1666464484
transform 1 0 20148 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_214
timestamp 1666464484
transform 1 0 20792 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1666464484
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1666464484
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_246
timestamp 1666464484
transform 1 0 23736 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_252
timestamp 1666464484
transform 1 0 24288 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_260
timestamp 1666464484
transform 1 0 25024 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_271
timestamp 1666464484
transform 1 0 26036 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1666464484
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_288
timestamp 1666464484
transform 1 0 27600 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_296
timestamp 1666464484
transform 1 0 28336 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_303
timestamp 1666464484
transform 1 0 28980 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_310
timestamp 1666464484
transform 1 0 29624 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_317
timestamp 1666464484
transform 1 0 30268 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1666464484
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_90
timestamp 1666464484
transform 1 0 9384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_96
timestamp 1666464484
transform 1 0 9936 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_102
timestamp 1666464484
transform 1 0 10488 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_108
timestamp 1666464484
transform 1 0 11040 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_114
timestamp 1666464484
transform 1 0 11592 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_120
timestamp 1666464484
transform 1 0 12144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_126
timestamp 1666464484
transform 1 0 12696 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_132
timestamp 1666464484
transform 1 0 13248 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1666464484
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1666464484
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_150
timestamp 1666464484
transform 1 0 14904 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_156
timestamp 1666464484
transform 1 0 15456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_162
timestamp 1666464484
transform 1 0 16008 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1666464484
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_174
timestamp 1666464484
transform 1 0 17112 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_180
timestamp 1666464484
transform 1 0 17664 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1666464484
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1666464484
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_201
timestamp 1666464484
transform 1 0 19596 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_209
timestamp 1666464484
transform 1 0 20332 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1666464484
transform 1 0 20700 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_217
timestamp 1666464484
transform 1 0 21068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_224
timestamp 1666464484
transform 1 0 21712 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_232
timestamp 1666464484
transform 1 0 22448 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_241
timestamp 1666464484
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1666464484
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_263
timestamp 1666464484
transform 1 0 25300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_272
timestamp 1666464484
transform 1 0 26128 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_281
timestamp 1666464484
transform 1 0 26956 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_296
timestamp 1666464484
transform 1 0 28336 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1666464484
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_314
timestamp 1666464484
transform 1 0 29992 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_325
timestamp 1666464484
transform 1 0 31004 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_329
timestamp 1666464484
transform 1 0 31372 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_8
timestamp 1666464484
transform 1 0 1840 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_20
timestamp 1666464484
transform 1 0 2944 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_32
timestamp 1666464484
transform 1 0 4048 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_44
timestamp 1666464484
transform 1 0 5152 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_86
timestamp 1666464484
transform 1 0 9016 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_92
timestamp 1666464484
transform 1 0 9568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_98
timestamp 1666464484
transform 1 0 10120 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_104
timestamp 1666464484
transform 1 0 10672 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1666464484
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1666464484
transform 1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_124
timestamp 1666464484
transform 1 0 12512 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_130
timestamp 1666464484
transform 1 0 13064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1666464484
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_142
timestamp 1666464484
transform 1 0 14168 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_148
timestamp 1666464484
transform 1 0 14720 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_154
timestamp 1666464484
transform 1 0 15272 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_160
timestamp 1666464484
transform 1 0 15824 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1666464484
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1666464484
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_176
timestamp 1666464484
transform 1 0 17296 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_182
timestamp 1666464484
transform 1 0 17848 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_188
timestamp 1666464484
transform 1 0 18400 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_194
timestamp 1666464484
transform 1 0 18952 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_200
timestamp 1666464484
transform 1 0 19504 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_203
timestamp 1666464484
transform 1 0 19780 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_209
timestamp 1666464484
transform 1 0 20332 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_212
timestamp 1666464484
transform 1 0 20608 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_218
timestamp 1666464484
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_229
timestamp 1666464484
transform 1 0 22172 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_233
timestamp 1666464484
transform 1 0 22540 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_241
timestamp 1666464484
transform 1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_250
timestamp 1666464484
transform 1 0 24104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_259
timestamp 1666464484
transform 1 0 24932 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_268
timestamp 1666464484
transform 1 0 25760 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1666464484
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_286
timestamp 1666464484
transform 1 0 27416 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_300
timestamp 1666464484
transform 1 0 28704 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_307
timestamp 1666464484
transform 1 0 29348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_314
timestamp 1666464484
transform 1 0 29992 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_321
timestamp 1666464484
transform 1 0 30636 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_93
timestamp 1666464484
transform 1 0 9660 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_96
timestamp 1666464484
transform 1 0 9936 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_102
timestamp 1666464484
transform 1 0 10488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_108
timestamp 1666464484
transform 1 0 11040 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_114
timestamp 1666464484
transform 1 0 11592 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_120
timestamp 1666464484
transform 1 0 12144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_126
timestamp 1666464484
transform 1 0 12696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_132
timestamp 1666464484
transform 1 0 13248 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1666464484
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1666464484
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_152
timestamp 1666464484
transform 1 0 15088 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_158
timestamp 1666464484
transform 1 0 15640 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_164
timestamp 1666464484
transform 1 0 16192 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_170
timestamp 1666464484
transform 1 0 16744 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_176
timestamp 1666464484
transform 1 0 17296 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_182
timestamp 1666464484
transform 1 0 17848 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_188
timestamp 1666464484
transform 1 0 18400 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_202
timestamp 1666464484
transform 1 0 19688 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1666464484
transform 1 0 20424 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_216
timestamp 1666464484
transform 1 0 20976 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_224
timestamp 1666464484
transform 1 0 21712 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_227
timestamp 1666464484
transform 1 0 21988 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_231
timestamp 1666464484
transform 1 0 22356 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_235
timestamp 1666464484
transform 1 0 22724 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_242
timestamp 1666464484
transform 1 0 23368 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1666464484
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_260
timestamp 1666464484
transform 1 0 25024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_269
timestamp 1666464484
transform 1 0 25852 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_284
timestamp 1666464484
transform 1 0 27232 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1666464484
transform 1 0 27876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_297
timestamp 1666464484
transform 1 0 28428 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1666464484
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_316
timestamp 1666464484
transform 1 0 30176 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_322
timestamp 1666464484
transform 1 0 30728 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_329
timestamp 1666464484
transform 1 0 31372 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_8
timestamp 1666464484
transform 1 0 1840 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_20
timestamp 1666464484
transform 1 0 2944 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_32
timestamp 1666464484
transform 1 0 4048 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_44
timestamp 1666464484
transform 1 0 5152 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_101
timestamp 1666464484
transform 1 0 10396 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_104
timestamp 1666464484
transform 1 0 10672 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1666464484
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1666464484
transform 1 0 11960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_124
timestamp 1666464484
transform 1 0 12512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_130
timestamp 1666464484
transform 1 0 13064 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1666464484
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_142
timestamp 1666464484
transform 1 0 14168 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_148
timestamp 1666464484
transform 1 0 14720 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_154
timestamp 1666464484
transform 1 0 15272 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_160
timestamp 1666464484
transform 1 0 15824 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1666464484
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_175
timestamp 1666464484
transform 1 0 17204 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_178
timestamp 1666464484
transform 1 0 17480 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_184
timestamp 1666464484
transform 1 0 18032 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_190
timestamp 1666464484
transform 1 0 18584 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_196
timestamp 1666464484
transform 1 0 19136 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_204
timestamp 1666464484
transform 1 0 19872 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_214
timestamp 1666464484
transform 1 0 20792 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1666464484
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_229
timestamp 1666464484
transform 1 0 22172 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_235
timestamp 1666464484
transform 1 0 22724 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_238
timestamp 1666464484
transform 1 0 23000 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_242
timestamp 1666464484
transform 1 0 23368 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_246
timestamp 1666464484
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_253
timestamp 1666464484
transform 1 0 24380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_257
timestamp 1666464484
transform 1 0 24748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_262
timestamp 1666464484
transform 1 0 25208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_269
timestamp 1666464484
transform 1 0 25852 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1666464484
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_285
timestamp 1666464484
transform 1 0 27324 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_291
timestamp 1666464484
transform 1 0 27876 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_297
timestamp 1666464484
transform 1 0 28428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_303
timestamp 1666464484
transform 1 0 28980 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_311
timestamp 1666464484
transform 1 0 29716 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_315
timestamp 1666464484
transform 1 0 30084 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_322
timestamp 1666464484
transform 1 0 30728 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_8
timestamp 1666464484
transform 1 0 1840 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_20
timestamp 1666464484
transform 1 0 2944 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_114
timestamp 1666464484
transform 1 0 11592 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_120
timestamp 1666464484
transform 1 0 12144 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_126
timestamp 1666464484
transform 1 0 12696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_132
timestamp 1666464484
transform 1 0 13248 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1666464484
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_146
timestamp 1666464484
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_152
timestamp 1666464484
transform 1 0 15088 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_158
timestamp 1666464484
transform 1 0 15640 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_164
timestamp 1666464484
transform 1 0 16192 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp 1666464484
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_176
timestamp 1666464484
transform 1 0 17296 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_182
timestamp 1666464484
transform 1 0 17848 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_188
timestamp 1666464484
transform 1 0 18400 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1666464484
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_205
timestamp 1666464484
transform 1 0 19964 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_213
timestamp 1666464484
transform 1 0 20700 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_219
timestamp 1666464484
transform 1 0 21252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_225
timestamp 1666464484
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_228
timestamp 1666464484
transform 1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_234
timestamp 1666464484
transform 1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_240
timestamp 1666464484
transform 1 0 23184 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1666464484
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_258
timestamp 1666464484
transform 1 0 24840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_265
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_272
timestamp 1666464484
transform 1 0 26128 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_278
timestamp 1666464484
transform 1 0 26680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_284
timestamp 1666464484
transform 1 0 27232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_290
timestamp 1666464484
transform 1 0 27784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_296
timestamp 1666464484
transform 1 0 28336 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_302
timestamp 1666464484
transform 1 0 28888 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_313
timestamp 1666464484
transform 1 0 29900 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_317
timestamp 1666464484
transform 1 0 30268 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_329
timestamp 1666464484
transform 1 0 31372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_8
timestamp 1666464484
transform 1 0 1840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_22
timestamp 1666464484
transform 1 0 3128 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_29
timestamp 1666464484
transform 1 0 3772 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_37
timestamp 1666464484
transform 1 0 4508 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_41
timestamp 1666464484
transform 1 0 4876 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_49
timestamp 1666464484
transform 1 0 5612 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1666464484
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_80
timestamp 1666464484
transform 1 0 8464 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_85
timestamp 1666464484
transform 1 0 8924 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_89
timestamp 1666464484
transform 1 0 9292 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_119
timestamp 1666464484
transform 1 0 12052 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_132
timestamp 1666464484
transform 1 0 13248 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_138
timestamp 1666464484
transform 1 0 13800 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_141
timestamp 1666464484
transform 1 0 14076 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_145
timestamp 1666464484
transform 1 0 14444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_151
timestamp 1666464484
transform 1 0 14996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_158
timestamp 1666464484
transform 1 0 15640 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1666464484
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_174
timestamp 1666464484
transform 1 0 17112 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_182
timestamp 1666464484
transform 1 0 17848 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_188
timestamp 1666464484
transform 1 0 18400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_194
timestamp 1666464484
transform 1 0 18952 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_197
timestamp 1666464484
transform 1 0 19228 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_202
timestamp 1666464484
transform 1 0 19688 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_206
timestamp 1666464484
transform 1 0 20056 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_210
timestamp 1666464484
transform 1 0 20424 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_216
timestamp 1666464484
transform 1 0 20976 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1666464484
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_229
timestamp 1666464484
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_236
timestamp 1666464484
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_242
timestamp 1666464484
transform 1 0 23368 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_249
timestamp 1666464484
transform 1 0 24012 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_253
timestamp 1666464484
transform 1 0 24380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_257
timestamp 1666464484
transform 1 0 24748 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_265
timestamp 1666464484
transform 1 0 25484 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_271
timestamp 1666464484
transform 1 0 26036 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1666464484
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666464484
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_288
timestamp 1666464484
transform 1 0 27600 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_298
timestamp 1666464484
transform 1 0 28520 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_304
timestamp 1666464484
transform 1 0 29072 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_309
timestamp 1666464484
transform 1 0 29532 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_314
timestamp 1666464484
transform 1 0 29992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_320
timestamp 1666464484
transform 1 0 30544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_327
timestamp 1666464484
transform 1 0 31188 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 31832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 31832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 31832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 31832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 31832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 31832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 31832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 31832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 31832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 31832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 31832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 31832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 31832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 31832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 31832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 31832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 31832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 31832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 31832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 31832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 31832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 31832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 31832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 31832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 31832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 31832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 31832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 31832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 31832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 31832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 31832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 31832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 31832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 31832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 31832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 31832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 31832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 31832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 31832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 31832 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 31832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 31832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 31832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 31832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 31832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 31832 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 31832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 31832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 31832 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 31832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 31832 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 31832 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 31832 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 31832 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 8832 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 24288 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 29440 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _0438_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23736 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0439_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22816 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0440_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0441_
timestamp 1666464484
transform 1 0 22448 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0442_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24104 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0443_
timestamp 1666464484
transform 1 0 27784 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0444_
timestamp 1666464484
transform -1 0 16008 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0445_
timestamp 1666464484
transform -1 0 15548 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0446_
timestamp 1666464484
transform 1 0 19872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0447_
timestamp 1666464484
transform -1 0 15088 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0448_
timestamp 1666464484
transform 1 0 15916 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0449_
timestamp 1666464484
transform -1 0 13340 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0450_
timestamp 1666464484
transform 1 0 18308 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0451_
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0452_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0453_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17296 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0454_
timestamp 1666464484
transform 1 0 25208 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _0455_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0456_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18584 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0457_
timestamp 1666464484
transform -1 0 22540 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0458_
timestamp 1666464484
transform 1 0 24564 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0459_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0460_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16928 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0461_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19964 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0462_
timestamp 1666464484
transform 1 0 12880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0463_
timestamp 1666464484
transform -1 0 20792 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0464_
timestamp 1666464484
transform -1 0 17480 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0465_
timestamp 1666464484
transform -1 0 14904 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0466_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0468_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26680 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0469_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19872 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0470_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0471_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28888 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0472_
timestamp 1666464484
transform -1 0 28336 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0473_
timestamp 1666464484
transform -1 0 26128 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0474_
timestamp 1666464484
transform 1 0 28060 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0475_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1666464484
transform -1 0 25024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0477_
timestamp 1666464484
transform -1 0 25760 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0478_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25668 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0479_
timestamp 1666464484
transform 1 0 29716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _0480_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0481_
timestamp 1666464484
transform -1 0 27968 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0482_
timestamp 1666464484
transform -1 0 26772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0483_
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0484_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0485_
timestamp 1666464484
transform -1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0486_
timestamp 1666464484
transform -1 0 25208 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0487_
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0488_
timestamp 1666464484
transform 1 0 28888 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _0489_
timestamp 1666464484
transform -1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0490_
timestamp 1666464484
transform 1 0 25208 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0491_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0492_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29992 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0493_
timestamp 1666464484
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0494_
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0495_
timestamp 1666464484
transform -1 0 27416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0496_
timestamp 1666464484
transform -1 0 28796 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0497_
timestamp 1666464484
transform -1 0 27784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0498_
timestamp 1666464484
transform -1 0 30176 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0499_
timestamp 1666464484
transform -1 0 28060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0500_
timestamp 1666464484
transform -1 0 31372 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0501_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0502_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0503_
timestamp 1666464484
transform -1 0 27048 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1666464484
transform -1 0 26128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1666464484
transform 1 0 28980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0506_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19228 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0507_
timestamp 1666464484
transform 1 0 10488 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0508_
timestamp 1666464484
transform 1 0 18492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1666464484
transform 1 0 26404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0510_
timestamp 1666464484
transform -1 0 26220 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0511_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23552 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _0512_
timestamp 1666464484
transform -1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _0513_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _0514_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23644 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0515_
timestamp 1666464484
transform -1 0 18400 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0516_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20240 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0517_
timestamp 1666464484
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0518_
timestamp 1666464484
transform 1 0 14996 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0519_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15732 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0520_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0521_
timestamp 1666464484
transform 1 0 15088 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0522_
timestamp 1666464484
transform -1 0 30084 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0523_
timestamp 1666464484
transform -1 0 12972 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0524_
timestamp 1666464484
transform 1 0 13064 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0525_
timestamp 1666464484
transform 1 0 23184 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0526_
timestamp 1666464484
transform 1 0 26404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1666464484
transform -1 0 23736 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0528_
timestamp 1666464484
transform -1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0529_
timestamp 1666464484
transform 1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0530_
timestamp 1666464484
transform -1 0 11224 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0531_
timestamp 1666464484
transform 1 0 13432 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1666464484
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0533_
timestamp 1666464484
transform 1 0 16100 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0534_
timestamp 1666464484
transform -1 0 19780 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0535_
timestamp 1666464484
transform -1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0536_
timestamp 1666464484
transform 1 0 16100 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0537_
timestamp 1666464484
transform -1 0 16376 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0538_
timestamp 1666464484
transform -1 0 13800 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0539_
timestamp 1666464484
transform 1 0 14904 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0540_
timestamp 1666464484
transform 1 0 15272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0541_
timestamp 1666464484
transform -1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0542_
timestamp 1666464484
transform -1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _0543_
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0544_
timestamp 1666464484
transform 1 0 12972 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0545_
timestamp 1666464484
transform -1 0 17848 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1666464484
transform -1 0 9844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0547_
timestamp 1666464484
transform -1 0 14720 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1666464484
transform -1 0 10488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0549_
timestamp 1666464484
transform 1 0 17572 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0550_
timestamp 1666464484
transform -1 0 16376 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0551_
timestamp 1666464484
transform -1 0 14720 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1666464484
transform -1 0 13064 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0553_
timestamp 1666464484
transform 1 0 16100 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0554_
timestamp 1666464484
transform 1 0 13984 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0555_
timestamp 1666464484
transform -1 0 20608 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0556_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21528 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0557_
timestamp 1666464484
transform -1 0 15364 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0558_
timestamp 1666464484
transform -1 0 21068 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0559_
timestamp 1666464484
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0560_
timestamp 1666464484
transform 1 0 26404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0561_
timestamp 1666464484
transform 1 0 12144 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1666464484
transform 1 0 12788 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0563_
timestamp 1666464484
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0564_
timestamp 1666464484
transform 1 0 11684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0565_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17940 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0566_
timestamp 1666464484
transform -1 0 18124 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0567_
timestamp 1666464484
transform 1 0 17480 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1666464484
transform 1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0569_
timestamp 1666464484
transform -1 0 21528 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1666464484
transform -1 0 19688 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0571_
timestamp 1666464484
transform 1 0 15548 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0572_
timestamp 1666464484
transform -1 0 19688 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0573_
timestamp 1666464484
transform -1 0 24104 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0574_
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0575_
timestamp 1666464484
transform 1 0 17204 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0576_
timestamp 1666464484
transform -1 0 14904 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0577_
timestamp 1666464484
transform -1 0 18952 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0578_
timestamp 1666464484
transform -1 0 15180 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0579_
timestamp 1666464484
transform 1 0 14076 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1666464484
transform 1 0 24196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0581_
timestamp 1666464484
transform -1 0 31372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0582_
timestamp 1666464484
transform -1 0 19228 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0583_
timestamp 1666464484
transform -1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0584_
timestamp 1666464484
transform -1 0 24840 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0585_
timestamp 1666464484
transform -1 0 22448 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0586_
timestamp 1666464484
transform 1 0 22816 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0587_
timestamp 1666464484
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0588_
timestamp 1666464484
transform 1 0 28428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0589_
timestamp 1666464484
transform -1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0590_
timestamp 1666464484
transform 1 0 18308 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0591_
timestamp 1666464484
transform -1 0 19320 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0592_
timestamp 1666464484
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0593_
timestamp 1666464484
transform -1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0594_
timestamp 1666464484
transform 1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0595_
timestamp 1666464484
transform -1 0 25208 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0596_
timestamp 1666464484
transform -1 0 21528 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _0597_
timestamp 1666464484
transform -1 0 14260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0598_
timestamp 1666464484
transform 1 0 17848 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0599_
timestamp 1666464484
transform -1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0600_
timestamp 1666464484
transform 1 0 17388 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0601_
timestamp 1666464484
transform -1 0 15272 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0602_
timestamp 1666464484
transform 1 0 17296 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0603_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1666464484
transform -1 0 14076 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0605_
timestamp 1666464484
transform 1 0 18308 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0606_
timestamp 1666464484
transform -1 0 16928 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0607_
timestamp 1666464484
transform 1 0 14536 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0608_
timestamp 1666464484
transform -1 0 21528 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1666464484
transform -1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1666464484
transform -1 0 18952 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0611_
timestamp 1666464484
transform 1 0 17572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1666464484
transform 1 0 19412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0613_
timestamp 1666464484
transform -1 0 15732 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _0614_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14720 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0615_
timestamp 1666464484
transform 1 0 19412 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1666464484
transform -1 0 12420 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0617_
timestamp 1666464484
transform -1 0 16744 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0618_
timestamp 1666464484
transform 1 0 13248 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0619_
timestamp 1666464484
transform -1 0 20148 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0620_
timestamp 1666464484
transform -1 0 13800 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0621_
timestamp 1666464484
transform 1 0 14168 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0622_
timestamp 1666464484
transform 1 0 18308 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0623_
timestamp 1666464484
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0624_
timestamp 1666464484
transform -1 0 13064 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0625_
timestamp 1666464484
transform 1 0 20976 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0626_
timestamp 1666464484
transform -1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0627_
timestamp 1666464484
transform 1 0 13892 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0628_
timestamp 1666464484
transform -1 0 17940 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0629_
timestamp 1666464484
transform 1 0 14352 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0630_
timestamp 1666464484
transform -1 0 17940 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1666464484
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0632_
timestamp 1666464484
transform -1 0 15456 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1666464484
transform -1 0 13064 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0634_
timestamp 1666464484
transform -1 0 21252 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1666464484
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0636_
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0637_
timestamp 1666464484
transform 1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0638_
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0639_
timestamp 1666464484
transform 1 0 16100 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0640_
timestamp 1666464484
transform -1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0641_
timestamp 1666464484
transform 1 0 13064 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1666464484
transform -1 0 21712 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0643_
timestamp 1666464484
transform 1 0 25668 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0644_
timestamp 1666464484
transform -1 0 16376 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0645_
timestamp 1666464484
transform -1 0 26312 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0646_
timestamp 1666464484
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0647_
timestamp 1666464484
transform -1 0 29624 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0648_
timestamp 1666464484
transform 1 0 11500 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1666464484
transform 1 0 12144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0650_
timestamp 1666464484
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0651_
timestamp 1666464484
transform 1 0 29072 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0652_
timestamp 1666464484
transform 1 0 28336 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0653_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30636 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0654_
timestamp 1666464484
transform -1 0 28704 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0655_
timestamp 1666464484
transform -1 0 28704 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0656_
timestamp 1666464484
transform 1 0 29348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0657_
timestamp 1666464484
transform -1 0 27416 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0658_
timestamp 1666464484
transform 1 0 29256 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0659_
timestamp 1666464484
transform -1 0 27140 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1666464484
transform -1 0 30268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1666464484
transform 1 0 26220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _0662_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0663_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29164 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0664_
timestamp 1666464484
transform 1 0 19596 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _0665_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23460 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0666_
timestamp 1666464484
transform 1 0 27140 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0667_
timestamp 1666464484
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0668_
timestamp 1666464484
transform -1 0 27600 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0669_
timestamp 1666464484
transform -1 0 24840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  _0670_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__nor3_4  _0671_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27968 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__a211oi_1  _0672_
timestamp 1666464484
transform -1 0 20332 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0673_
timestamp 1666464484
transform -1 0 30452 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0674_
timestamp 1666464484
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0675_
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 1666464484
transform 1 0 28704 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0677_
timestamp 1666464484
transform -1 0 27692 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0678_
timestamp 1666464484
transform -1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0679_
timestamp 1666464484
transform 1 0 30912 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0680_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26312 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0681_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0682_
timestamp 1666464484
transform 1 0 22080 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 1666464484
transform 1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0684_
timestamp 1666464484
transform 1 0 29716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_2  _0685_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__a211oi_1  _0686_
timestamp 1666464484
transform -1 0 29716 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0687_
timestamp 1666464484
transform -1 0 31004 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0688_
timestamp 1666464484
transform -1 0 30360 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0689_
timestamp 1666464484
transform 1 0 18952 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1666464484
transform 1 0 11592 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0691_
timestamp 1666464484
transform 1 0 18952 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0692_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27324 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0693_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24104 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0694_
timestamp 1666464484
transform 1 0 22448 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0695_
timestamp 1666464484
transform 1 0 24840 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1666464484
transform 1 0 30084 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0697_
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0698_
timestamp 1666464484
transform -1 0 24472 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0699_
timestamp 1666464484
transform -1 0 12788 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0700_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30452 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1666464484
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0702_
timestamp 1666464484
transform -1 0 25300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0703_
timestamp 1666464484
transform -1 0 31280 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0704_
timestamp 1666464484
transform -1 0 28980 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0705_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27692 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0706_
timestamp 1666464484
transform -1 0 27784 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0707_
timestamp 1666464484
transform 1 0 24472 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0708_
timestamp 1666464484
transform 1 0 26128 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _0709_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0710_
timestamp 1666464484
transform 1 0 27968 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0711_
timestamp 1666464484
transform -1 0 30360 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _0712_
timestamp 1666464484
transform -1 0 22816 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0713_
timestamp 1666464484
transform -1 0 31096 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0714_
timestamp 1666464484
transform -1 0 12420 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0715_
timestamp 1666464484
transform -1 0 24380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0716_
timestamp 1666464484
transform 1 0 29716 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0717_
timestamp 1666464484
transform -1 0 20608 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0718_
timestamp 1666464484
transform 1 0 18124 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0719_
timestamp 1666464484
transform 1 0 24840 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0720_
timestamp 1666464484
transform 1 0 14168 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0721_
timestamp 1666464484
transform 1 0 26772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0722_
timestamp 1666464484
transform -1 0 29164 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0723_
timestamp 1666464484
transform -1 0 30452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1666464484
transform -1 0 21712 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0725_
timestamp 1666464484
transform -1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0726_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29532 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0727_
timestamp 1666464484
transform -1 0 22264 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0728_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0729_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27600 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0730_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29532 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0731_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0732_
timestamp 1666464484
transform -1 0 26588 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0733_
timestamp 1666464484
transform 1 0 19320 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0734_
timestamp 1666464484
transform 1 0 15732 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1666464484
transform -1 0 19044 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0736_
timestamp 1666464484
transform 1 0 17112 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0737_
timestamp 1666464484
transform 1 0 10856 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 1666464484
transform 1 0 19780 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0739_
timestamp 1666464484
transform -1 0 14352 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0740_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18216 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0741_
timestamp 1666464484
transform 1 0 21160 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0742_
timestamp 1666464484
transform -1 0 22724 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1666464484
transform 1 0 10948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0744_
timestamp 1666464484
transform 1 0 14996 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0745_
timestamp 1666464484
transform -1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1666464484
transform 1 0 21988 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0747_
timestamp 1666464484
transform 1 0 15732 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1666464484
transform 1 0 9568 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0749_
timestamp 1666464484
transform -1 0 15824 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0750_
timestamp 1666464484
transform -1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0751_
timestamp 1666464484
transform 1 0 30728 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0752_
timestamp 1666464484
transform 1 0 21712 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0753_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0754_
timestamp 1666464484
transform -1 0 19412 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0755_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19228 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0756_
timestamp 1666464484
transform 1 0 15088 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0757_
timestamp 1666464484
transform -1 0 30452 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 1666464484
transform 1 0 16376 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _0759_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31372 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0760_
timestamp 1666464484
transform 1 0 17112 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0761_
timestamp 1666464484
transform -1 0 16836 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0762_
timestamp 1666464484
transform 1 0 16928 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0763_
timestamp 1666464484
transform -1 0 20792 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0764_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0765_
timestamp 1666464484
transform -1 0 18952 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0766_
timestamp 1666464484
transform 1 0 18308 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0767_
timestamp 1666464484
transform -1 0 18952 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0768_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22080 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0769_
timestamp 1666464484
transform -1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0770_
timestamp 1666464484
transform -1 0 18952 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0771_
timestamp 1666464484
transform -1 0 17848 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _0772_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0773_
timestamp 1666464484
transform 1 0 14720 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1666464484
transform -1 0 30176 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0775_
timestamp 1666464484
transform 1 0 17020 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0776_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31372 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0777_
timestamp 1666464484
transform 1 0 16744 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0778_
timestamp 1666464484
transform 1 0 22264 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0779_
timestamp 1666464484
transform 1 0 25392 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1666464484
transform 1 0 26312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0781_
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0782_
timestamp 1666464484
transform 1 0 30636 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1666464484
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0784_
timestamp 1666464484
transform -1 0 25484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0785_
timestamp 1666464484
transform 1 0 11316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0786_
timestamp 1666464484
transform 1 0 30820 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0787_
timestamp 1666464484
transform 1 0 25300 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0788_
timestamp 1666464484
transform 1 0 29992 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0789_
timestamp 1666464484
transform 1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1666464484
transform 1 0 26404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0791_
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0792_
timestamp 1666464484
transform 1 0 28060 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0793_
timestamp 1666464484
transform 1 0 10948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0794_
timestamp 1666464484
transform 1 0 11684 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0795_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0796_
timestamp 1666464484
transform 1 0 29716 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1666464484
transform 1 0 27876 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0798_
timestamp 1666464484
transform -1 0 27324 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0799_
timestamp 1666464484
transform -1 0 21528 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _0800_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12972 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0801_
timestamp 1666464484
transform 1 0 27140 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0802_
timestamp 1666464484
transform -1 0 31280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _0803_
timestamp 1666464484
transform 1 0 28428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0804_
timestamp 1666464484
transform -1 0 23920 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0805_
timestamp 1666464484
transform -1 0 30820 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0806_
timestamp 1666464484
transform 1 0 17296 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0807_
timestamp 1666464484
transform -1 0 16376 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0808_
timestamp 1666464484
transform -1 0 26220 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0809_
timestamp 1666464484
transform 1 0 24840 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _0810_
timestamp 1666464484
transform 1 0 21160 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0811_
timestamp 1666464484
transform 1 0 24196 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _0812_
timestamp 1666464484
transform 1 0 13156 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0813_
timestamp 1666464484
transform -1 0 16836 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0814_
timestamp 1666464484
transform 1 0 14720 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _0815_
timestamp 1666464484
transform -1 0 27968 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _0816_
timestamp 1666464484
transform -1 0 30084 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1666464484
transform 1 0 22448 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0818_
timestamp 1666464484
transform 1 0 18308 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0819_
timestamp 1666464484
transform -1 0 29256 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0820_
timestamp 1666464484
transform 1 0 22448 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _0821_
timestamp 1666464484
transform -1 0 15364 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0822_
timestamp 1666464484
transform 1 0 30452 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0823_
timestamp 1666464484
transform 1 0 12420 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0824_
timestamp 1666464484
transform 1 0 21988 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0825_
timestamp 1666464484
transform -1 0 16376 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0826_
timestamp 1666464484
transform -1 0 13800 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _0827_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28704 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0828_
timestamp 1666464484
transform -1 0 17848 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 1666464484
transform 1 0 12604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0830_
timestamp 1666464484
transform -1 0 23184 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0831_
timestamp 1666464484
transform -1 0 17848 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1666464484
transform 1 0 10212 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0833_
timestamp 1666464484
transform 1 0 13892 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0834_
timestamp 1666464484
transform -1 0 12696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0835_
timestamp 1666464484
transform 1 0 14444 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0836_
timestamp 1666464484
transform 1 0 13432 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0837_
timestamp 1666464484
transform -1 0 10580 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0838_
timestamp 1666464484
transform -1 0 31372 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0839_
timestamp 1666464484
transform 1 0 20884 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0840_
timestamp 1666464484
transform 1 0 22632 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0841_
timestamp 1666464484
transform 1 0 15732 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0842_
timestamp 1666464484
transform -1 0 18952 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_2  _0843_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21896 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0844_
timestamp 1666464484
transform 1 0 30820 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1666464484
transform -1 0 19964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0846_
timestamp 1666464484
transform -1 0 23828 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0847_
timestamp 1666464484
transform 1 0 13248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _0848_
timestamp 1666464484
transform -1 0 23736 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0849_
timestamp 1666464484
transform 1 0 27968 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0850_
timestamp 1666464484
transform -1 0 30912 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0851_
timestamp 1666464484
transform -1 0 25300 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0852_
timestamp 1666464484
transform 1 0 24380 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0853_
timestamp 1666464484
transform -1 0 21344 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0854_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _0855_
timestamp 1666464484
transform 1 0 12144 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0856_
timestamp 1666464484
transform -1 0 27784 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0857_
timestamp 1666464484
transform 1 0 23644 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0858_
timestamp 1666464484
transform 1 0 25852 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0859_
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0860_
timestamp 1666464484
transform 1 0 26496 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1666464484
transform -1 0 23368 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0862_
timestamp 1666464484
transform 1 0 15548 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _0863_
timestamp 1666464484
transform 1 0 28336 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _0864_
timestamp 1666464484
transform -1 0 24472 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0865_
timestamp 1666464484
transform -1 0 26036 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0866_
timestamp 1666464484
transform 1 0 29348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0867_
timestamp 1666464484
transform -1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _0868_
timestamp 1666464484
transform -1 0 25300 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0869_
timestamp 1666464484
transform -1 0 23460 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0870_
timestamp 1666464484
transform -1 0 28796 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0871_
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0872_
timestamp 1666464484
transform -1 0 27876 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0873_
timestamp 1666464484
transform -1 0 27876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0874_
timestamp 1666464484
transform -1 0 30820 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0875_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30268 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1666464484
transform 1 0 18676 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1666464484
transform 1 0 30360 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1666464484
transform -1 0 28980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1666464484
transform 1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1666464484
transform 1 0 26956 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1666464484
transform 1 0 20792 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1666464484
transform 1 0 17940 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1666464484
transform 1 0 23460 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1666464484
transform 1 0 15456 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1666464484
transform 1 0 20516 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0886_
timestamp 1666464484
transform 1 0 30176 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1666464484
transform -1 0 29992 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1666464484
transform -1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1666464484
transform -1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1666464484
transform 1 0 27784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1666464484
transform 1 0 30728 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1666464484
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1666464484
transform -1 0 28704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1666464484
transform -1 0 30360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1666464484
transform -1 0 29348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1666464484
transform -1 0 26772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0897_
timestamp 1666464484
transform -1 0 15824 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1666464484
transform 1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1666464484
transform 1 0 11960 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1666464484
transform 1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1666464484
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1666464484
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1666464484
transform 1 0 10212 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1666464484
transform 1 0 12788 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1666464484
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1666464484
transform 1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1666464484
transform 1 0 11960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0908_
timestamp 1666464484
transform 1 0 27140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1666464484
transform 1 0 11500 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1666464484
transform 1 0 12144 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1666464484
transform 1 0 22172 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1666464484
transform -1 0 23552 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1666464484
transform 1 0 29716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1666464484
transform 1 0 22632 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1666464484
transform -1 0 29716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1666464484
transform 1 0 21528 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1666464484
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1666464484
transform -1 0 21160 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0919_
timestamp 1666464484
transform -1 0 29256 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1666464484
transform 1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1666464484
transform 1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1666464484
transform -1 0 19044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1666464484
transform 1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1666464484
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1666464484
transform 1 0 19688 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1666464484
transform 1 0 17020 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1666464484
transform 1 0 11684 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1666464484
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0930_
timestamp 1666464484
transform -1 0 28244 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1666464484
transform 1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1666464484
transform -1 0 24380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1666464484
transform -1 0 23644 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1666464484
transform 1 0 22724 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1666464484
transform 1 0 22080 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1666464484
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1666464484
transform 1 0 11500 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1666464484
transform 1 0 23552 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1666464484
transform -1 0 23092 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1666464484
transform -1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1666464484
transform -1 0 25944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _0942_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25116 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0943_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21896 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1666464484
transform 1 0 22264 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0945_
timestamp 1666464484
transform 1 0 24564 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0946_
timestamp 1666464484
transform 1 0 26864 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0947_
timestamp 1666464484
transform 1 0 24564 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1666464484
transform 1 0 22264 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0949_
timestamp 1666464484
transform 1 0 23276 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1666464484
transform -1 0 24104 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0951_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23184 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0952_
timestamp 1666464484
transform -1 0 26404 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0953_
timestamp 1666464484
transform -1 0 26496 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1666464484
transform -1 0 26404 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1666464484
transform 1 0 27140 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0956_
timestamp 1666464484
transform -1 0 26680 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1666464484
transform 1 0 26956 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0958_
timestamp 1666464484
transform 1 0 27140 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0959_
timestamp 1666464484
transform -1 0 26588 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0960_
timestamp 1666464484
transform -1 0 26680 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0961_
timestamp 1666464484
transform -1 0 26588 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0962_
timestamp 1666464484
transform -1 0 23920 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0963_
timestamp 1666464484
transform 1 0 21988 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0964_
timestamp 1666464484
transform -1 0 21436 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0965_
timestamp 1666464484
transform 1 0 19412 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0966_
timestamp 1666464484
transform 1 0 19964 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0967_
timestamp 1666464484
transform -1 0 23736 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0968_
timestamp 1666464484
transform 1 0 19964 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0969_
timestamp 1666464484
transform 1 0 20056 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0970_
timestamp 1666464484
transform 1 0 19596 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0971_
timestamp 1666464484
transform -1 0 21528 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0972_
timestamp 1666464484
transform -1 0 22448 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0973_
timestamp 1666464484
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0974_
timestamp 1666464484
transform 1 0 24196 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0975_
timestamp 1666464484
transform 1 0 20608 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0976_
timestamp 1666464484
transform 1 0 21988 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0977_
timestamp 1666464484
transform 1 0 21620 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0978_
timestamp 1666464484
transform 1 0 21988 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0979_
timestamp 1666464484
transform 1 0 24564 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0980_
timestamp 1666464484
transform 1 0 24196 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0981_
timestamp 1666464484
transform 1 0 19688 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0982_
timestamp 1666464484
transform -1 0 21252 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0983_
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0984_
timestamp 1666464484
transform -1 0 18952 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0985_
timestamp 1666464484
transform -1 0 20240 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0986_
timestamp 1666464484
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0987_
timestamp 1666464484
transform -1 0 23460 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0988_
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0989_
timestamp 1666464484
transform 1 0 18768 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0990_
timestamp 1666464484
transform -1 0 20700 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0991_
timestamp 1666464484
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0992_
timestamp 1666464484
transform -1 0 18952 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0993_
timestamp 1666464484
transform -1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0994_
timestamp 1666464484
transform -1 0 23828 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0995_
timestamp 1666464484
transform 1 0 24288 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0996_
timestamp 1666464484
transform 1 0 21620 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0997_
timestamp 1666464484
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0998_
timestamp 1666464484
transform 1 0 19596 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0999_
timestamp 1666464484
transform -1 0 26404 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1000_
timestamp 1666464484
transform -1 0 23920 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1001_
timestamp 1666464484
transform 1 0 22264 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1002_
timestamp 1666464484
transform 1 0 24564 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1666464484
transform -1 0 30636 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1666464484
transform -1 0 30636 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1666464484
transform -1 0 29992 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1077_
timestamp 1666464484
transform -1 0 30176 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1666464484
transform -1 0 29348 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout8
timestamp 1666464484
transform 1 0 16836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout9
timestamp 1666464484
transform -1 0 18492 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout10
timestamp 1666464484
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout11
timestamp 1666464484
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1666464484
transform -1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1666464484
transform -1 0 30912 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 1666464484
transform 1 0 28704 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout15
timestamp 1666464484
transform -1 0 26588 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform 1 0 30452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 31096 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1666464484
transform 1 0 31004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform 1 0 31004 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform 1 0 31004 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform 1 0 31004 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_17
timestamp 1666464484
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_18
timestamp 1666464484
transform 1 0 31096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_19
timestamp 1666464484
transform 1 0 31096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_20
timestamp 1666464484
transform 1 0 31096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_21
timestamp 1666464484
transform 1 0 29808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_22
timestamp 1666464484
transform 1 0 31096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_23
timestamp 1666464484
transform 1 0 30452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_24
timestamp 1666464484
transform 1 0 31096 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_25
timestamp 1666464484
transform 1 0 29716 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_26
timestamp 1666464484
transform 1 0 31096 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_27
timestamp 1666464484
transform 1 0 31096 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_28
timestamp 1666464484
transform 1 0 30452 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_29
timestamp 1666464484
transform 1 0 29808 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_30
timestamp 1666464484
transform 1 0 30360 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_31
timestamp 1666464484
transform -1 0 29992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_32
timestamp 1666464484
transform -1 0 26404 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33
timestamp 1666464484
transform -1 0 22816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform -1 0 19688 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform -1 0 15640 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform -1 0 12052 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform -1 0 8464 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform -1 0 4876 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform -1 0 1840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform -1 0 1840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform -1 0 1840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform -1 0 1840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform -1 0 1840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform -1 0 1840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform -1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform -1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform -1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform 1 0 31096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform 1 0 31096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform 1 0 31096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform 1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform 1 0 31096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform 1 0 31096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform 1 0 30452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform 1 0 29808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform 1 0 31096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform 1 0 31096 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform -1 0 31188 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform -1 0 27600 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform -1 0 24012 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform -1 0 20424 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform -1 0 17112 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 13248 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 9660 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform -1 0 6072 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform -1 0 2484 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform -1 0 3128 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform -1 0 1840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform -1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform -1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_77
timestamp 1666464484
transform -1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_78
timestamp 1666464484
transform -1 0 1840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_79
timestamp 1666464484
transform -1 0 1840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_80
timestamp 1666464484
transform -1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_81
timestamp 1666464484
transform -1 0 1840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_82
timestamp 1666464484
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_83
timestamp 1666464484
transform -1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_84
timestamp 1666464484
transform -1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_85
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_86
timestamp 1666464484
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
<< labels >>
flabel metal3 s 32206 2456 33006 2576 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 32206 22856 33006 22976 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 32206 24896 33006 25016 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 32206 26936 33006 27056 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 32206 28976 33006 29096 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 32206 31016 33006 31136 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 32034 34350 32090 35150 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 28446 34350 28502 35150 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 24858 34350 24914 35150 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 21270 34350 21326 35150 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 17682 34350 17738 35150 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 32206 4496 33006 4616 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 14094 34350 14150 35150 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 10506 34350 10562 35150 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 6918 34350 6974 35150 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 3330 34350 3386 35150 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 31696 800 31816 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 32206 6536 33006 6656 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 32206 8576 33006 8696 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 32206 10616 33006 10736 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 32206 12656 33006 12776 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 32206 14696 33006 14816 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 32206 16736 33006 16856 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 32206 18776 33006 18896 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 32206 20816 33006 20936 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 32206 3816 33006 3936 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 32206 24216 33006 24336 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 32206 26256 33006 26376 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 32206 28296 33006 28416 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 32206 30336 33006 30456 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 32206 32376 33006 32496 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 29642 34350 29698 35150 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 26054 34350 26110 35150 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 22466 34350 22522 35150 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 18878 34350 18934 35150 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 15290 34350 15346 35150 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 32206 5856 33006 5976 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 11702 34350 11758 35150 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 8114 34350 8170 35150 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 4526 34350 4582 35150 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 938 34350 994 35150 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 30064 800 30184 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 32206 7896 33006 8016 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 32206 9936 33006 10056 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 32206 11976 33006 12096 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 32206 14016 33006 14136 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 32206 16056 33006 16176 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 32206 18096 33006 18216 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 32206 20136 33006 20256 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 32206 22176 33006 22296 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 32206 3136 33006 3256 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 32206 23536 33006 23656 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 32206 25576 33006 25696 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 32206 27616 33006 27736 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 32206 29656 33006 29776 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 32206 31696 33006 31816 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 30838 34350 30894 35150 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 27250 34350 27306 35150 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 23662 34350 23718 35150 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 20074 34350 20130 35150 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 16486 34350 16542 35150 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 32206 5176 33006 5296 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 12898 34350 12954 35150 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 9310 34350 9366 35150 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 5722 34350 5778 35150 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 2134 34350 2190 35150 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 32206 7216 33006 7336 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 32206 9256 33006 9376 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 32206 11296 33006 11416 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 32206 13336 33006 13456 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 32206 15376 33006 15496 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 32206 17416 33006 17536 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 32206 19456 33006 19576 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 32206 21496 33006 21616 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4785 2128 5105 32688 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 12467 2128 12787 32688 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 20149 2128 20469 32688 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 27831 2128 28151 32688 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 8626 2128 8946 32688 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 16308 2128 16628 32688 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 23990 2128 24310 32688 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 31672 2128 31992 32688 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 16468 32096 16468 32096 0 vccd1
rlabel via1 16548 32640 16548 32640 0 vssd1
rlabel metal2 19642 28288 19642 28288 0 _0000_
rlabel metal2 30406 28441 30406 28441 0 _0001_
rlabel metal1 24019 25262 24019 25262 0 _0002_
rlabel metal2 13662 25619 13662 25619 0 _0003_
rlabel metal1 27784 30770 27784 30770 0 _0004_
rlabel metal1 22264 30362 22264 30362 0 _0005_
rlabel metal2 18354 27353 18354 27353 0 _0006_
rlabel metal1 23959 24854 23959 24854 0 _0007_
rlabel metal2 22126 22440 22126 22440 0 _0008_
rlabel metal2 20654 29427 20654 29427 0 _0009_
rlabel metal2 25346 22389 25346 22389 0 _0010_
rlabel via3 24771 18020 24771 18020 0 _0011_
rlabel metal1 22954 11696 22954 11696 0 _0012_
rlabel metal1 28060 13498 28060 13498 0 _0013_
rlabel metal1 30682 15062 30682 15062 0 _0014_
rlabel metal1 27324 12954 27324 12954 0 _0015_
rlabel metal2 28566 15147 28566 15147 0 _0016_
rlabel metal1 30130 14926 30130 14926 0 _0017_
rlabel metal3 25783 16524 25783 16524 0 _0018_
rlabel metal2 25254 20771 25254 20771 0 _0019_
rlabel via2 9706 20315 9706 20315 0 _0020_
rlabel metal2 12098 21981 12098 21981 0 _0021_
rlabel metal1 19727 21930 19727 21930 0 _0022_
rlabel metal4 13340 21828 13340 21828 0 _0023_
rlabel metal1 13202 18768 13202 18768 0 _0024_
rlabel metal3 15525 11764 15525 11764 0 _0025_
rlabel metal2 17434 11900 17434 11900 0 _0026_
rlabel metal1 21627 19754 21627 19754 0 _0027_
rlabel metal1 20187 19414 20187 19414 0 _0028_
rlabel metal2 12098 19533 12098 19533 0 _0029_
rlabel metal2 21022 16269 21022 16269 0 _0030_
rlabel via2 14122 18309 14122 18309 0 _0031_
rlabel metal1 23782 10166 23782 10166 0 _0032_
rlabel metal1 22954 10710 22954 10710 0 _0033_
rlabel metal2 29854 13566 29854 13566 0 _0034_
rlabel metal1 22724 10778 22724 10778 0 _0035_
rlabel metal1 25162 13906 25162 13906 0 _0036_
rlabel metal1 23322 15606 23322 15606 0 _0037_
rlabel metal2 20010 11764 20010 11764 0 _0038_
rlabel metal2 21022 11560 21022 11560 0 _0039_
rlabel metal1 17940 12750 17940 12750 0 _0040_
rlabel metal2 16974 13753 16974 13753 0 _0041_
rlabel metal1 18262 11662 18262 11662 0 _0042_
rlabel metal1 15410 14314 15410 14314 0 _0043_
rlabel metal1 16399 14042 16399 14042 0 _0044_
rlabel metal1 20838 11254 20838 11254 0 _0045_
rlabel metal1 14766 16150 14766 16150 0 _0046_
rlabel metal1 18032 13158 18032 13158 0 _0047_
rlabel metal1 17240 17136 17240 17136 0 _0048_
rlabel metal1 14766 14858 14766 14858 0 _0049_
rlabel via2 13478 17595 13478 17595 0 _0050_
rlabel metal2 21482 13379 21482 13379 0 _0051_
rlabel metal2 23506 12614 23506 12614 0 _0052_
rlabel metal2 23230 15708 23230 15708 0 _0053_
rlabel metal1 22303 15402 22303 15402 0 _0054_
rlabel metal1 22671 16150 22671 16150 0 _0055_
rlabel metal2 13478 15215 13478 15215 0 _0056_
rlabel metal1 24334 12342 24334 12342 0 _0057_
rlabel metal2 22954 14552 22954 14552 0 _0058_
rlabel metal1 23835 19414 23835 19414 0 _0059_
rlabel metal1 25852 12954 25852 12954 0 _0060_
rlabel metal1 27830 30260 27830 30260 0 _0061_
rlabel metal1 22494 30736 22494 30736 0 _0062_
rlabel via2 23230 30005 23230 30005 0 _0063_
rlabel metal3 16031 27540 16031 27540 0 _0064_
rlabel metal2 13294 24531 13294 24531 0 _0065_
rlabel metal2 15042 27676 15042 27676 0 _0066_
rlabel metal1 27002 27404 27002 27404 0 _0067_
rlabel metal1 13294 24922 13294 24922 0 _0068_
rlabel metal1 16376 24310 16376 24310 0 _0069_
rlabel metal1 8004 27846 8004 27846 0 _0070_
rlabel metal1 6946 24786 6946 24786 0 _0071_
rlabel metal1 9200 28594 9200 28594 0 _0072_
rlabel metal4 14076 9644 14076 9644 0 _0073_
rlabel metal1 18860 27574 18860 27574 0 _0074_
rlabel metal3 14329 12308 14329 12308 0 _0075_
rlabel metal1 12144 24242 12144 24242 0 _0076_
rlabel metal2 17434 21743 17434 21743 0 _0077_
rlabel metal1 9315 25942 9315 25942 0 _0078_
rlabel metal1 17434 27030 17434 27030 0 _0079_
rlabel metal2 16790 25041 16790 25041 0 _0080_
rlabel metal1 14168 24718 14168 24718 0 _0081_
rlabel metal1 21114 25840 21114 25840 0 _0082_
rlabel metal1 14963 24786 14963 24786 0 _0083_
rlabel metal1 28336 29002 28336 29002 0 _0084_
rlabel metal2 2714 18275 2714 18275 0 _0085_
rlabel metal1 11500 29138 11500 29138 0 _0086_
rlabel metal2 31878 17238 31878 17238 0 _0087_
rlabel metal2 27554 26860 27554 26860 0 _0088_
rlabel metal2 30682 21743 30682 21743 0 _0089_
rlabel metal2 14122 24684 14122 24684 0 _0090_
rlabel metal2 29670 17340 29670 17340 0 _0091_
rlabel metal1 28934 19278 28934 19278 0 _0092_
rlabel metal1 28060 4726 28060 4726 0 _0093_
rlabel metal1 28428 19414 28428 19414 0 _0094_
rlabel metal1 29808 19142 29808 19142 0 _0095_
rlabel metal3 16123 7956 16123 7956 0 _0096_
rlabel metal1 30958 24174 30958 24174 0 _0097_
rlabel metal1 29900 19278 29900 19278 0 _0098_
rlabel metal2 27646 14416 27646 14416 0 _0099_
rlabel metal1 25622 13804 25622 13804 0 _0100_
rlabel metal1 27186 13328 27186 13328 0 _0101_
rlabel metal1 28750 18190 28750 18190 0 _0102_
rlabel metal2 27830 14212 27830 14212 0 _0103_
rlabel metal1 30682 17578 30682 17578 0 _0104_
rlabel metal2 26818 14960 26818 14960 0 _0105_
rlabel via1 26810 14314 26810 14314 0 _0106_
rlabel metal1 25990 12206 25990 12206 0 _0107_
rlabel metal1 8142 21386 8142 21386 0 _0108_
rlabel metal1 14536 20910 14536 20910 0 _0109_
rlabel metal1 13294 19414 13294 19414 0 _0110_
rlabel metal2 19182 19431 19182 19431 0 _0111_
rlabel metal1 25530 15912 25530 15912 0 _0112_
rlabel metal1 24564 14382 24564 14382 0 _0113_
rlabel metal2 15410 14348 15410 14348 0 _0114_
rlabel metal2 16100 17476 16100 17476 0 _0115_
rlabel metal2 28106 16099 28106 16099 0 _0116_
rlabel metal1 18216 15878 18216 15878 0 _0117_
rlabel metal1 16330 18190 16330 18190 0 _0118_
rlabel metal2 18262 11900 18262 11900 0 _0119_
rlabel metal1 15686 16218 15686 16218 0 _0120_
rlabel metal1 15640 16422 15640 16422 0 _0121_
rlabel metal1 17158 17204 17158 17204 0 _0122_
rlabel metal1 17199 17306 17199 17306 0 _0123_
rlabel via2 10534 16949 10534 16949 0 _0124_
rlabel via3 13317 19380 13317 19380 0 _0125_
rlabel metal1 18630 19924 18630 19924 0 _0126_
rlabel metal2 13754 18836 13754 18836 0 _0127_
rlabel via2 17802 11883 17802 11883 0 _0128_
rlabel metal1 11730 19822 11730 19822 0 _0129_
rlabel metal2 11178 19448 11178 19448 0 _0130_
rlabel metal2 14950 23596 14950 23596 0 _0131_
rlabel metal1 9936 20842 9936 20842 0 _0132_
rlabel metal1 18400 21658 18400 21658 0 _0133_
rlabel metal1 16739 15674 16739 15674 0 _0134_
rlabel metal1 13900 18258 13900 18258 0 _0135_
rlabel metal1 19412 17646 19412 17646 0 _0136_
rlabel metal1 15226 25194 15226 25194 0 _0137_
rlabel metal1 13524 21590 13524 21590 0 _0138_
rlabel metal1 13428 20910 13428 20910 0 _0139_
rlabel metal1 13754 20808 13754 20808 0 _0140_
rlabel metal1 13938 21114 13938 21114 0 _0141_
rlabel metal1 14030 22712 14030 22712 0 _0142_
rlabel metal1 20286 23018 20286 23018 0 _0143_
rlabel metal2 10626 21284 10626 21284 0 _0144_
rlabel metal2 14490 23392 14490 23392 0 _0145_
rlabel metal1 14528 21930 14528 21930 0 _0146_
rlabel metal2 14306 22882 14306 22882 0 _0147_
rlabel metal2 20700 25228 20700 25228 0 _0148_
rlabel metal1 19458 23188 19458 23188 0 _0149_
rlabel metal1 20240 25398 20240 25398 0 _0150_
rlabel metal1 15410 22678 15410 22678 0 _0151_
rlabel metal1 23322 10472 23322 10472 0 _0152_
rlabel metal2 17066 18887 17066 18887 0 _0153_
rlabel metal2 12834 18428 12834 18428 0 _0154_
rlabel metal1 16882 19312 16882 19312 0 _0155_
rlabel metal2 13570 19618 13570 19618 0 _0156_
rlabel metal1 20194 16966 20194 16966 0 _0157_
rlabel metal1 23874 16490 23874 16490 0 _0158_
rlabel metal2 23966 17034 23966 17034 0 _0159_
rlabel metal1 20286 17306 20286 17306 0 _0160_
rlabel metal1 16606 18802 16606 18802 0 _0161_
rlabel metal1 24196 10438 24196 10438 0 _0162_
rlabel metal1 23230 18870 23230 18870 0 _0163_
rlabel metal1 14766 19414 14766 19414 0 _0164_
rlabel metal1 18446 19788 18446 19788 0 _0165_
rlabel metal1 14536 18938 14536 18938 0 _0166_
rlabel metal1 18814 20400 18814 20400 0 _0167_
rlabel metal2 30498 18547 30498 18547 0 _0168_
rlabel metal1 31004 18394 31004 18394 0 _0169_
rlabel metal1 21160 11866 21160 11866 0 _0170_
rlabel viali 15959 13294 15959 13294 0 _0171_
rlabel metal1 20286 10608 20286 10608 0 _0172_
rlabel metal1 15502 13872 15502 13872 0 _0173_
rlabel metal2 14674 14586 14674 14586 0 _0174_
rlabel metal1 14858 14042 14858 14042 0 _0175_
rlabel metal2 21482 14756 21482 14756 0 _0176_
rlabel metal1 14536 16082 14536 16082 0 _0177_
rlabel metal1 17940 12410 17940 12410 0 _0178_
rlabel metal1 16422 14416 16422 14416 0 _0179_
rlabel metal2 17342 14722 17342 14722 0 _0180_
rlabel metal1 13846 14960 13846 14960 0 _0181_
rlabel metal1 20240 13702 20240 13702 0 _0182_
rlabel metal1 14904 15674 14904 15674 0 _0183_
rlabel metal2 18262 13430 18262 13430 0 _0184_
rlabel metal1 16284 12342 16284 12342 0 _0185_
rlabel metal1 19458 11764 19458 11764 0 _0186_
rlabel metal2 16514 14858 16514 14858 0 _0187_
rlabel metal1 15226 15674 15226 15674 0 _0188_
rlabel metal1 19734 17612 19734 17612 0 _0189_
rlabel metal2 16238 16252 16238 16252 0 _0190_
rlabel via2 13386 15861 13386 15861 0 _0191_
rlabel metal1 15778 14416 15778 14416 0 _0192_
rlabel metal1 17959 18156 17959 18156 0 _0193_
rlabel metal1 20378 16150 20378 16150 0 _0194_
rlabel metal1 21252 16082 21252 16082 0 _0195_
rlabel metal1 16422 13464 16422 13464 0 _0196_
rlabel metal2 14306 15062 14306 15062 0 _0197_
rlabel metal1 15226 17816 15226 17816 0 _0198_
rlabel metal2 13478 11735 13478 11735 0 _0199_
rlabel metal1 15356 18394 15356 18394 0 _0200_
rlabel metal1 13938 17646 13938 17646 0 _0201_
rlabel metal1 15870 14552 15870 14552 0 _0202_
rlabel metal2 12282 16235 12282 16235 0 _0203_
rlabel via2 20930 10795 20930 10795 0 _0204_
rlabel metal1 13524 16966 13524 16966 0 _0205_
rlabel via1 13302 17238 13302 17238 0 _0206_
rlabel metal2 21482 11373 21482 11373 0 _0207_
rlabel metal2 21482 16082 21482 16082 0 _0208_
rlabel metal2 21574 13260 21574 13260 0 _0209_
rlabel viali 11727 16558 11727 16558 0 _0210_
rlabel via2 29210 17051 29210 17051 0 _0211_
rlabel via2 14582 17867 14582 17867 0 _0212_
rlabel metal3 23230 34340 23230 34340 0 _0213_
rlabel metal1 31326 23766 31326 23766 0 _0214_
rlabel metal2 30682 25755 30682 25755 0 _0215_
rlabel metal2 28198 28407 28198 28407 0 _0216_
rlabel metal2 29762 27404 29762 27404 0 _0217_
rlabel metal2 21482 29529 21482 29529 0 _0218_
rlabel metal1 29256 26010 29256 26010 0 _0219_
rlabel metal1 26634 28628 26634 28628 0 _0220_
rlabel via1 27187 26350 27187 26350 0 _0221_
rlabel metal1 26818 22066 26818 22066 0 _0222_
rlabel metal2 9522 28458 9522 28458 0 _0223_
rlabel metal1 5980 24038 5980 24038 0 _0224_
rlabel metal1 8556 28526 8556 28526 0 _0225_
rlabel metal1 12374 23800 12374 23800 0 _0226_
rlabel metal2 7130 23188 7130 23188 0 _0227_
rlabel metal1 14858 24140 14858 24140 0 _0228_
rlabel metal1 24610 31994 24610 31994 0 _0229_
rlabel metal1 6348 28390 6348 28390 0 _0230_
rlabel metal1 5060 24786 5060 24786 0 _0231_
rlabel metal1 29900 27387 29900 27387 0 _0232_
rlabel metal1 29670 24378 29670 24378 0 _0233_
rlabel metal1 30866 26248 30866 26248 0 _0234_
rlabel metal2 30958 25415 30958 25415 0 _0235_
rlabel metal1 29210 29274 29210 29274 0 _0236_
rlabel metal2 8234 13709 8234 13709 0 _0237_
rlabel metal1 31004 27030 31004 27030 0 _0238_
rlabel metal1 25438 29614 25438 29614 0 _0239_
rlabel metal1 26082 25738 26082 25738 0 _0240_
rlabel metal2 6302 26248 6302 26248 0 _0241_
rlabel metal2 25806 30260 25806 30260 0 _0242_
rlabel metal1 27600 31926 27600 31926 0 _0243_
rlabel metal1 24748 26962 24748 26962 0 _0244_
rlabel metal2 8418 27744 8418 27744 0 _0245_
rlabel metal1 29026 27030 29026 27030 0 _0246_
rlabel metal2 30958 16473 30958 16473 0 _0247_
rlabel metal4 6532 11276 6532 11276 0 _0248_
rlabel metal1 16008 31450 16008 31450 0 _0249_
rlabel via3 5451 9588 5451 9588 0 _0250_
rlabel metal2 9798 25466 9798 25466 0 _0251_
rlabel metal1 29854 23086 29854 23086 0 _0252_
rlabel metal2 8234 27200 8234 27200 0 _0253_
rlabel via2 21390 26197 21390 26197 0 _0254_
rlabel metal3 22724 33388 22724 33388 0 _0255_
rlabel via2 17158 30651 17158 30651 0 _0256_
rlabel metal2 12190 6085 12190 6085 0 _0257_
rlabel metal2 12742 23052 12742 23052 0 _0258_
rlabel metal1 18354 33490 18354 33490 0 _0259_
rlabel metal1 30452 24786 30452 24786 0 _0260_
rlabel via2 30866 26333 30866 26333 0 _0261_
rlabel metal1 27462 17068 27462 17068 0 _0262_
rlabel metal1 29716 15402 29716 15402 0 _0263_
rlabel via2 8050 27387 8050 27387 0 _0264_
rlabel metal2 7406 11752 7406 11752 0 _0265_
rlabel metal2 11592 20060 11592 20060 0 _0266_
rlabel metal1 25944 30226 25944 30226 0 _0267_
rlabel metal1 5382 21862 5382 21862 0 _0268_
rlabel via2 30038 23715 30038 23715 0 _0269_
rlabel metal3 21252 33932 21252 33932 0 _0270_
rlabel metal2 22494 23052 22494 23052 0 _0271_
rlabel metal1 29900 22610 29900 22610 0 _0272_
rlabel via1 9614 23171 9614 23171 0 _0273_
rlabel metal3 12581 8364 12581 8364 0 _0274_
rlabel metal2 25254 28560 25254 28560 0 _0275_
rlabel metal1 13294 29818 13294 29818 0 _0276_
rlabel metal3 21781 19516 21781 19516 0 _0277_
rlabel metal1 24932 28050 24932 28050 0 _0278_
rlabel metal1 27406 25296 27406 25296 0 _0279_
rlabel metal1 5658 27370 5658 27370 0 _0280_
rlabel metal2 27462 18921 27462 18921 0 _0281_
rlabel metal3 21436 26928 21436 26928 0 _0282_
rlabel metal1 24978 23256 24978 23256 0 _0283_
rlabel metal1 18076 29546 18076 29546 0 _0284_
rlabel metal2 10350 9282 10350 9282 0 _0285_
rlabel metal2 30314 22270 30314 22270 0 _0286_
rlabel metal2 13478 22253 13478 22253 0 _0287_
rlabel metal1 28060 23290 28060 23290 0 _0288_
rlabel metal1 26680 25466 26680 25466 0 _0289_
rlabel metal1 29348 23834 29348 23834 0 _0290_
rlabel metal1 26128 30702 26128 30702 0 _0291_
rlabel metal1 24334 30669 24334 30669 0 _0292_
rlabel metal2 18446 21386 18446 21386 0 _0293_
rlabel metal1 22724 24718 22724 24718 0 _0294_
rlabel metal1 17848 22474 17848 22474 0 _0295_
rlabel metal1 11224 21658 11224 21658 0 _0296_
rlabel metal1 21068 24582 21068 24582 0 _0297_
rlabel metal1 14628 21658 14628 21658 0 _0298_
rlabel metal1 18538 22032 18538 22032 0 _0299_
rlabel metal1 17920 23596 17920 23596 0 _0300_
rlabel metal1 5244 21590 5244 21590 0 _0301_
rlabel metal1 11592 22746 11592 22746 0 _0302_
rlabel metal2 22218 27982 22218 27982 0 _0303_
rlabel metal1 20700 27914 20700 27914 0 _0304_
rlabel metal1 15732 22542 15732 22542 0 _0305_
rlabel metal1 16606 23120 16606 23120 0 _0306_
rlabel metal1 10902 22134 10902 22134 0 _0307_
rlabel via2 4738 21981 4738 21981 0 _0308_
rlabel metal1 12052 21862 12052 21862 0 _0309_
rlabel metal2 29670 22576 29670 22576 0 _0310_
rlabel metal1 21022 24684 21022 24684 0 _0311_
rlabel metal1 19733 23732 19733 23732 0 _0312_
rlabel via1 19923 23720 19923 23720 0 _0313_
rlabel metal2 17434 22066 17434 22066 0 _0314_
rlabel via2 16422 26333 16422 26333 0 _0315_
rlabel metal1 30360 21862 30360 21862 0 _0316_
rlabel metal1 17480 22066 17480 22066 0 _0317_
rlabel metal2 17802 21777 17802 21777 0 _0318_
rlabel metal1 16836 21930 16836 21930 0 _0319_
rlabel metal1 16836 23086 16836 23086 0 _0320_
rlabel metal1 18446 22576 18446 22576 0 _0321_
rlabel metal1 18308 22610 18308 22610 0 _0322_
rlabel metal1 18354 22474 18354 22474 0 _0323_
rlabel metal2 18906 23120 18906 23120 0 _0324_
rlabel metal1 18354 25466 18354 25466 0 _0325_
rlabel metal1 18768 25126 18768 25126 0 _0326_
rlabel metal1 19182 25976 19182 25976 0 _0327_
rlabel metal2 18630 27285 18630 27285 0 _0328_
rlabel metal2 17342 23783 17342 23783 0 _0329_
rlabel metal2 25254 31127 25254 31127 0 _0330_
rlabel metal2 9614 32241 9614 32241 0 _0331_
rlabel metal1 15088 24378 15088 24378 0 _0332_
rlabel metal1 29716 27642 29716 27642 0 _0333_
rlabel metal1 22287 27302 22287 27302 0 _0334_
rlabel metal1 30774 25160 30774 25160 0 _0335_
rlabel via2 17158 25483 17158 25483 0 _0336_
rlabel metal1 24526 30770 24526 30770 0 _0337_
rlabel metal2 27554 25823 27554 25823 0 _0338_
rlabel metal1 27370 19210 27370 19210 0 _0339_
rlabel via3 10925 20740 10925 20740 0 _0340_
rlabel metal1 8602 21930 8602 21930 0 _0341_
rlabel metal1 26358 12274 26358 12274 0 _0342_
rlabel via2 12558 20893 12558 20893 0 _0343_
rlabel metal3 18055 34068 18055 34068 0 _0344_
rlabel metal1 31464 24038 31464 24038 0 _0345_
rlabel metal4 17204 18836 17204 18836 0 _0346_
rlabel metal2 32614 24412 32614 24412 0 _0347_
rlabel metal1 12880 31110 12880 31110 0 _0348_
rlabel metal2 31188 21046 31188 21046 0 _0349_
rlabel metal4 15916 14658 15916 14658 0 _0350_
rlabel metal4 16100 16116 16100 16116 0 _0351_
rlabel metal2 11270 20485 11270 20485 0 _0352_
rlabel metal2 20654 9282 20654 9282 0 _0353_
rlabel metal2 30222 19142 30222 19142 0 _0354_
rlabel metal2 29762 20111 29762 20111 0 _0355_
rlabel metal2 28244 22372 28244 22372 0 _0356_
rlabel metal2 26726 17697 26726 17697 0 _0357_
rlabel metal2 22954 27200 22954 27200 0 _0358_
rlabel metal1 12512 21114 12512 21114 0 _0359_
rlabel metal1 26496 24582 26496 24582 0 _0360_
rlabel metal2 25346 25228 25346 25228 0 _0361_
rlabel metal1 27406 23562 27406 23562 0 _0362_
rlabel metal1 24058 27438 24058 27438 0 _0363_
rlabel metal2 30774 27064 30774 27064 0 _0364_
rlabel metal1 15962 23732 15962 23732 0 _0365_
rlabel metal1 16376 23494 16376 23494 0 _0366_
rlabel metal1 21666 25228 21666 25228 0 _0367_
rlabel metal1 21850 25228 21850 25228 0 _0368_
rlabel metal2 21206 25823 21206 25823 0 _0369_
rlabel metal2 29900 20740 29900 20740 0 _0370_
rlabel metal2 28842 21505 28842 21505 0 _0371_
rlabel metal1 15042 20332 15042 20332 0 _0372_
rlabel metal2 15318 20621 15318 20621 0 _0373_
rlabel metal2 28750 22372 28750 22372 0 _0374_
rlabel metal1 29762 21318 29762 21318 0 _0375_
rlabel metal2 23506 20162 23506 20162 0 _0376_
rlabel metal1 19504 18870 19504 18870 0 _0377_
rlabel metal1 25484 20774 25484 20774 0 _0378_
rlabel metal1 25484 20978 25484 20978 0 _0379_
rlabel metal2 12650 21913 12650 21913 0 _0380_
rlabel metal2 30498 20077 30498 20077 0 _0381_
rlabel metal1 13248 22066 13248 22066 0 _0382_
rlabel metal1 19366 21114 19366 21114 0 _0383_
rlabel metal1 7452 20570 7452 20570 0 _0384_
rlabel via2 28382 32283 28382 32283 0 _0385_
rlabel via2 12834 23069 12834 23069 0 _0386_
rlabel metal1 17848 23154 17848 23154 0 _0387_
rlabel metal2 6670 28951 6670 28951 0 _0388_
rlabel metal1 23414 26350 23414 26350 0 _0389_
rlabel metal2 9614 23698 9614 23698 0 _0390_
rlabel metal1 11454 20570 11454 20570 0 _0391_
rlabel metal1 17112 32334 17112 32334 0 _0392_
rlabel metal3 18653 8636 18653 8636 0 _0393_
rlabel metal2 16146 31059 16146 31059 0 _0394_
rlabel metal2 21390 8092 21390 8092 0 _0395_
rlabel metal1 12788 27574 12788 27574 0 _0396_
rlabel metal1 31188 23154 31188 23154 0 _0397_
rlabel metal1 21942 25738 21942 25738 0 _0398_
rlabel metal1 23230 26384 23230 26384 0 _0399_
rlabel metal1 16652 20570 16652 20570 0 _0400_
rlabel metal1 21252 23018 21252 23018 0 _0401_
rlabel metal1 18446 23052 18446 23052 0 _0402_
rlabel via2 23690 29155 23690 29155 0 _0403_
rlabel metal1 22862 26350 22862 26350 0 _0404_
rlabel via3 12259 21692 12259 21692 0 _0405_
rlabel metal2 13294 21760 13294 21760 0 _0406_
rlabel via2 8234 22763 8234 22763 0 _0407_
rlabel metal2 30590 26452 30590 26452 0 _0408_
rlabel metal1 25806 27506 25806 27506 0 _0409_
rlabel metal1 18768 23120 18768 23120 0 _0410_
rlabel metal2 22034 26996 22034 26996 0 _0411_
rlabel metal1 19228 23086 19228 23086 0 _0412_
rlabel metal1 12650 21522 12650 21522 0 _0413_
rlabel via2 12558 21403 12558 21403 0 _0414_
rlabel metal1 27462 25840 27462 25840 0 _0415_
rlabel via1 26080 28050 26080 28050 0 _0416_
rlabel metal1 21298 28560 21298 28560 0 _0417_
rlabel metal2 26542 30277 26542 30277 0 _0418_
rlabel metal1 27324 25874 27324 25874 0 _0419_
rlabel metal2 23874 28730 23874 28730 0 _0420_
rlabel metal1 15502 24038 15502 24038 0 _0421_
rlabel metal4 24748 24548 24748 24548 0 _0422_
rlabel metal1 27870 26894 27870 26894 0 _0423_
rlabel metal1 25898 29274 25898 29274 0 _0424_
rlabel metal1 31326 24582 31326 24582 0 _0425_
rlabel metal2 23782 29920 23782 29920 0 _0426_
rlabel metal1 28555 26758 28555 26758 0 _0427_
rlabel metal2 28382 27506 28382 27506 0 _0428_
rlabel metal1 28106 27098 28106 27098 0 _0429_
rlabel metal1 27186 25908 27186 25908 0 _0430_
rlabel metal2 14306 10409 14306 10409 0 _0431_
rlabel metal1 30682 17714 30682 17714 0 _0432_
rlabel metal2 13386 30515 13386 30515 0 _0433_
rlabel metal1 12926 18734 12926 18734 0 _0434_
rlabel metal1 21344 10030 21344 10030 0 _0435_
rlabel metal2 16238 13090 16238 13090 0 _0436_
rlabel metal1 11224 17646 11224 17646 0 _0437_
rlabel metal1 30866 14382 30866 14382 0 io_in[8]
rlabel metal1 31280 13294 31280 13294 0 io_in[9]
rlabel metal1 30774 27846 30774 27846 0 io_out[10]
rlabel metal1 31280 28390 31280 28390 0 io_out[11]
rlabel metal2 31234 28339 31234 28339 0 io_out[12]
rlabel metal2 31234 29869 31234 29869 0 io_out[13]
rlabel metal2 31234 31841 31234 31841 0 io_out[14]
rlabel metal1 29026 30226 29026 30226 0 mod.thorkn_vgaclock.io_b
rlabel metal1 30222 30702 30222 30702 0 mod.thorkn_vgaclock.io_g
rlabel metal1 30406 29648 30406 29648 0 mod.thorkn_vgaclock.io_h_sync
rlabel metal2 29762 30532 29762 30532 0 mod.thorkn_vgaclock.io_r
rlabel metal2 30222 29750 30222 29750 0 mod.thorkn_vgaclock.io_v_sync
rlabel metal1 29026 9894 29026 9894 0 mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l39\[1\]
rlabel metal1 7820 22474 7820 22474 0 mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l45\[1\]
rlabel metal1 7544 20230 7544 20230 0 mod.thorkn_vgaclock.vga_content._zz_when_VgaContent_l51\[1\]
rlabel metal3 23368 13396 23368 13396 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[0\]
rlabel metal2 18906 14926 18906 14926 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[10\]
rlabel metal1 18998 12682 18998 12682 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[11\]
rlabel metal1 16917 16626 16917 16626 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[12\]
rlabel metal1 18078 16762 18078 16762 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[13\]
rlabel metal2 19734 16456 19734 16456 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[14\]
rlabel metal2 16974 15028 16974 15028 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[15\]
rlabel metal1 21068 16150 21068 16150 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[16\]
rlabel metal1 18584 13498 18584 13498 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[17\]
rlabel metal2 13018 17612 13018 17612 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[18\]
rlabel metal1 22494 14450 22494 14450 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[19\]
rlabel metal1 23966 13838 23966 13838 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[1\]
rlabel metal1 24058 15062 24058 15062 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[20\]
rlabel metal2 21666 14178 21666 14178 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[21\]
rlabel metal1 21344 15538 21344 15538 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[22\]
rlabel metal2 11638 16371 11638 16371 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[23\]
rlabel metal2 19918 18105 19918 18105 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[24\]
rlabel metal1 22310 12920 22310 12920 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[2\]
rlabel metal1 20378 10778 20378 10778 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[3\]
rlabel metal1 18768 13362 18768 13362 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[4\]
rlabel metal1 15088 14586 15088 14586 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[5\]
rlabel via2 14214 15963 14214 15963 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[6\]
rlabel metal1 19826 12886 19826 12886 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[7\]
rlabel metal1 20884 13226 20884 13226 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[8\]
rlabel metal2 14030 14280 14030 14280 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_valueNext\[9\]
rlabel metal1 22218 11594 22218 11594 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[0\]
rlabel metal1 15686 15368 15686 15368 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[10\]
rlabel metal2 17802 13804 17802 13804 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[11\]
rlabel metal1 18676 12206 18676 12206 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[12\]
rlabel metal1 19688 14246 19688 14246 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[13\]
rlabel metal1 14628 18054 14628 18054 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[14\]
rlabel metal1 13754 16456 13754 16456 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[15\]
rlabel metal1 21114 16048 21114 16048 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[16\]
rlabel metal1 21344 16762 21344 16762 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[17\]
rlabel metal1 17618 18224 17618 18224 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[18\]
rlabel metal1 20424 14246 20424 14246 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[19\]
rlabel metal1 24702 13906 24702 13906 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[1\]
rlabel metal1 24886 17578 24886 17578 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[20\]
rlabel metal1 25760 17646 25760 17646 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[21\]
rlabel metal2 26174 15980 26174 15980 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[22\]
rlabel metal2 17802 15827 17802 15827 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[23\]
rlabel metal1 12374 17714 12374 17714 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[24\]
rlabel metal1 24288 12750 24288 12750 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[2\]
rlabel metal2 24242 13532 24242 13532 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[3\]
rlabel via2 18538 13277 18538 13277 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[4\]
rlabel metal2 15134 13294 15134 13294 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[5\]
rlabel metal2 15686 13243 15686 13243 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[6\]
rlabel metal2 15410 15538 15410 15538 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[7\]
rlabel metal1 14950 16048 14950 16048 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[8\]
rlabel metal2 15226 15827 15226 15827 0 mod.thorkn_vgaclock.vga_content.clock_counters.c_counter_value\[9\]
rlabel metal1 26128 18666 26128 18666 0 mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext\[0\]
rlabel metal1 25668 15130 25668 15130 0 mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext\[1\]
rlabel metal3 14628 14620 14628 14620 0 mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext\[2\]
rlabel metal3 20700 19312 20700 19312 0 mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_valueNext\[3\]
rlabel metal2 12926 19822 12926 19822 0 mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value\[1\]
rlabel metal1 7452 19686 7452 19686 0 mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value\[2\]
rlabel metal2 9568 11764 9568 11764 0 mod.thorkn_vgaclock.vga_content.clock_counters.h_counter_value\[3\]
rlabel metal1 5888 21658 5888 21658 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes\[1\]
rlabel metal1 13064 21522 13064 21522 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes\[2\]
rlabel metal2 21022 21828 21022 21828 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes\[3\]
rlabel metal1 14260 20366 14260 20366 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes\[4\]
rlabel metal1 17158 25262 17158 25262 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_minutes\[5\]
rlabel metal2 19366 30651 19366 30651 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds\[1\]
rlabel metal1 23966 18870 23966 18870 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds\[2\]
rlabel metal2 12328 20740 12328 20740 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds\[3\]
rlabel metal1 10534 19788 10534 19788 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds\[4\]
rlabel metal2 14950 18547 14950 18547 0 mod.thorkn_vgaclock.vga_content.clock_counters.io_seconds\[5\]
rlabel metal1 17250 21114 17250 21114 0 mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext\[0\]
rlabel metal2 10442 20621 10442 20621 0 mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext\[1\]
rlabel metal3 13340 18904 13340 18904 0 mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext\[2\]
rlabel via3 17963 21964 17963 21964 0 mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext\[3\]
rlabel metal1 20427 20842 20427 20842 0 mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext\[4\]
rlabel metal1 22224 22202 22224 22202 0 mod.thorkn_vgaclock.vga_content.clock_counters.m_counter_valueNext\[5\]
rlabel metal1 19413 18802 19413 18802 0 mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext\[0\]
rlabel metal1 18630 18938 18630 18938 0 mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext\[1\]
rlabel via1 19921 19278 19921 19278 0 mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext\[2\]
rlabel metal2 21666 20162 21666 20162 0 mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext\[3\]
rlabel metal1 20700 17714 20700 17714 0 mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext\[4\]
rlabel metal1 22264 18326 22264 18326 0 mod.thorkn_vgaclock.vga_content.clock_counters.s_counter_valueNext\[5\]
rlabel metal1 24656 25942 24656 25942 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[0\]
rlabel metal1 22172 30634 22172 30634 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[1\]
rlabel metal1 22080 25330 22080 25330 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[2\]
rlabel metal2 21942 25313 21942 25313 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[3\]
rlabel metal4 20884 24752 20884 24752 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[4\]
rlabel metal1 23920 24242 23920 24242 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[5\]
rlabel metal1 22494 24242 22494 24242 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[6\]
rlabel metal2 22954 24514 22954 24514 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[7\]
rlabel metal1 24242 23018 24242 23018 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[8\]
rlabel via2 23506 23613 23506 23613 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_valueNext\[9\]
rlabel metal1 11914 26554 11914 26554 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[0\]
rlabel metal1 17710 24140 17710 24140 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[1\]
rlabel via1 29578 28050 29578 28050 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[2\]
rlabel metal2 7958 26146 7958 26146 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[3\]
rlabel metal1 7130 27302 7130 27302 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[4\]
rlabel metal1 12420 32198 12420 32198 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[5\]
rlabel metal1 13386 32198 13386 32198 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[6\]
rlabel metal2 9614 28866 9614 28866 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[7\]
rlabel metal1 25001 31314 25001 31314 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[8\]
rlabel metal1 9384 24786 9384 24786 0 mod.thorkn_vgaclock.vga_sync_gen.h_counter_value\[9\]
rlabel metal1 26229 22542 26229 22542 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[0\]
rlabel via3 26197 22100 26197 22100 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[1\]
rlabel metal2 31142 21233 31142 21233 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[2\]
rlabel metal1 27324 21590 27324 21590 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[3\]
rlabel metal1 29440 19278 29440 19278 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[4\]
rlabel metal2 27370 17034 27370 17034 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[5\]
rlabel metal2 28198 18530 28198 18530 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[6\]
rlabel metal1 28290 14042 28290 14042 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[7\]
rlabel metal1 29532 19210 29532 19210 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[8\]
rlabel metal3 25691 20740 25691 20740 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_valueNext\[9\]
rlabel metal1 26726 19822 26726 19822 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[0\]
rlabel metal2 5842 24718 5842 24718 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[1\]
rlabel metal1 25024 22950 25024 22950 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[2\]
rlabel metal1 28244 17238 28244 17238 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[3\]
rlabel metal2 14030 31008 14030 31008 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[4\]
rlabel metal2 29486 16864 29486 16864 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[5\]
rlabel metal1 27554 14416 27554 14416 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[6\]
rlabel metal2 24610 32946 24610 32946 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[7\]
rlabel metal2 4554 17901 4554 17901 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[8\]
rlabel metal1 5589 6834 5589 6834 0 mod.thorkn_vgaclock.vga_sync_gen.v_counter_value\[9\]
rlabel metal2 30498 14739 30498 14739 0 net1
rlabel metal2 12834 19737 12834 19737 0 net10
rlabel metal1 23092 13158 23092 13158 0 net11
rlabel metal2 26358 22848 26358 22848 0 net12
rlabel metal2 20746 10370 20746 10370 0 net13
rlabel metal3 17779 34612 17779 34612 0 net14
rlabel metal2 24058 13549 24058 13549 0 net15
rlabel via2 31326 3893 31326 3893 0 net16
rlabel metal2 31326 6001 31326 6001 0 net17
rlabel metal2 31326 8143 31326 8143 0 net18
rlabel via2 31326 10013 31326 10013 0 net19
rlabel metal1 30912 13498 30912 13498 0 net2
rlabel via2 31326 11747 31326 11747 0 net20
rlabel metal2 30038 13719 30038 13719 0 net21
rlabel metal2 31326 14467 31326 14467 0 net22
rlabel metal1 30774 13906 30774 13906 0 net23
rlabel metal1 31418 13906 31418 13906 0 net24
rlabel via2 29946 29597 29946 29597 0 net25
rlabel metal1 31464 30702 31464 30702 0 net26
rlabel metal1 31694 31110 31694 31110 0 net27
rlabel metal2 30682 29801 30682 29801 0 net28
rlabel metal2 30038 30889 30038 30889 0 net29
rlabel metal2 31050 28764 31050 28764 0 net3
rlabel metal2 30590 32215 30590 32215 0 net30
rlabel metal1 29716 32402 29716 32402 0 net31
rlabel metal1 26128 32402 26128 32402 0 net32
rlabel metal1 22540 32402 22540 32402 0 net33
rlabel metal1 19182 32402 19182 32402 0 net34
rlabel metal2 15410 33439 15410 33439 0 net35
rlabel metal2 11822 33439 11822 33439 0 net36
rlabel metal2 8234 33439 8234 33439 0 net37
rlabel metal2 4646 33439 4646 33439 0 net38
rlabel metal1 1288 32402 1288 32402 0 net39
rlabel metal1 30820 28526 30820 28526 0 net4
rlabel metal2 1610 32283 1610 32283 0 net40
rlabel metal3 1142 30124 1142 30124 0 net41
rlabel metal3 1142 27676 1142 27676 0 net42
rlabel metal3 1142 25228 1142 25228 0 net43
rlabel metal3 1142 22780 1142 22780 0 net44
rlabel metal3 1142 20332 1142 20332 0 net45
rlabel metal3 1142 17884 1142 17884 0 net46
rlabel metal3 1142 15436 1142 15436 0 net47
rlabel metal3 1142 12988 1142 12988 0 net48
rlabel metal3 1142 10540 1142 10540 0 net49
rlabel metal1 30728 29138 30728 29138 0 net5
rlabel metal3 1142 8092 1142 8092 0 net50
rlabel metal3 1142 5644 1142 5644 0 net51
rlabel metal3 1142 3196 1142 3196 0 net52
rlabel metal3 1050 748 1050 748 0 net53
rlabel via2 31326 3485 31326 3485 0 net54
rlabel metal2 31326 5457 31326 5457 0 net55
rlabel via2 31326 7259 31326 7259 0 net56
rlabel via2 31326 9333 31326 9333 0 net57
rlabel via2 31326 11339 31326 11339 0 net58
rlabel metal2 31372 12716 31372 12716 0 net59
rlabel metal1 31050 30260 31050 30260 0 net6
rlabel metal1 30728 13362 30728 13362 0 net60
rlabel metal1 29624 13838 29624 13838 0 net61
rlabel metal1 31372 14586 31372 14586 0 net62
rlabel metal3 31280 21692 31280 21692 0 net63
rlabel metal2 30958 33439 30958 33439 0 net64
rlabel metal1 27324 32402 27324 32402 0 net65
rlabel metal1 23736 32402 23736 32402 0 net66
rlabel metal1 20148 32402 20148 32402 0 net67
rlabel metal1 16790 32402 16790 32402 0 net68
rlabel metal2 13018 33439 13018 33439 0 net69
rlabel metal1 30452 31790 30452 31790 0 net7
rlabel metal2 9430 33439 9430 33439 0 net70
rlabel metal2 5842 33439 5842 33439 0 net71
rlabel metal2 2254 33439 2254 33439 0 net72
rlabel metal2 2898 32895 2898 32895 0 net73
rlabel metal3 1142 30940 1142 30940 0 net74
rlabel metal3 1142 28492 1142 28492 0 net75
rlabel metal3 1142 26044 1142 26044 0 net76
rlabel metal3 1142 23596 1142 23596 0 net77
rlabel metal3 1142 21148 1142 21148 0 net78
rlabel metal3 1142 18700 1142 18700 0 net79
rlabel metal2 23690 16490 23690 16490 0 net8
rlabel metal3 1142 16252 1142 16252 0 net80
rlabel metal3 1142 13804 1142 13804 0 net81
rlabel metal3 1142 11356 1142 11356 0 net82
rlabel metal3 1142 8908 1142 8908 0 net83
rlabel metal3 1142 6460 1142 6460 0 net84
rlabel metal3 1142 4012 1142 4012 0 net85
rlabel metal3 1142 1564 1142 1564 0 net86
rlabel metal2 20654 12313 20654 12313 0 net9
<< properties >>
string FIXED_BBOX 0 0 33006 35150
<< end >>
