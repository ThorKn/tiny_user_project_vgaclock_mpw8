magic
tech sky130A
magscale 1 2
timestamp 1672510421
<< viali >>
rect 1869 31433 1903 31467
rect 5181 31433 5215 31467
rect 9229 31433 9263 31467
rect 10241 31433 10275 31467
rect 11805 31433 11839 31467
rect 13461 31433 13495 31467
rect 14933 31433 14967 31467
rect 28181 31433 28215 31467
rect 12449 31365 12483 31399
rect 17776 31365 17810 31399
rect 21198 31365 21232 31399
rect 12679 31331 12713 31365
rect 2053 31297 2087 31331
rect 3985 31297 4019 31331
rect 5365 31297 5399 31331
rect 7113 31297 7147 31331
rect 8585 31297 8619 31331
rect 9413 31297 9447 31331
rect 10425 31297 10459 31331
rect 11161 31297 11195 31331
rect 11989 31297 12023 31331
rect 13277 31297 13311 31331
rect 13369 31297 13403 31331
rect 14473 31297 14507 31331
rect 16057 31297 16091 31331
rect 17049 31297 17083 31331
rect 17509 31297 17543 31331
rect 19625 31297 19659 31331
rect 23130 31297 23164 31331
rect 24860 31297 24894 31331
rect 26617 31297 26651 31331
rect 27169 31297 27203 31331
rect 27261 31297 27295 31331
rect 27445 31297 27479 31331
rect 27537 31297 27571 31331
rect 28365 31297 28399 31331
rect 2513 31229 2547 31263
rect 13737 31229 13771 31263
rect 16313 31229 16347 31263
rect 21465 31229 21499 31263
rect 23397 31229 23431 31263
rect 24593 31229 24627 31263
rect 14289 31161 14323 31195
rect 20085 31161 20119 31195
rect 22017 31161 22051 31195
rect 27721 31161 27755 31195
rect 3433 31093 3467 31127
rect 6009 31093 6043 31127
rect 6653 31093 6687 31127
rect 7941 31093 7975 31127
rect 10977 31093 11011 31127
rect 12633 31093 12667 31127
rect 12817 31093 12851 31127
rect 16865 31093 16899 31127
rect 18889 31093 18923 31127
rect 19441 31093 19475 31127
rect 23857 31093 23891 31127
rect 25973 31093 26007 31127
rect 26433 31093 26467 31127
rect 6193 30889 6227 30923
rect 9321 30889 9355 30923
rect 11621 30889 11655 30923
rect 11805 30889 11839 30923
rect 20637 30889 20671 30923
rect 7941 30821 7975 30855
rect 10149 30821 10183 30855
rect 17509 30821 17543 30855
rect 5181 30753 5215 30787
rect 12725 30753 12759 30787
rect 18889 30753 18923 30787
rect 21097 30753 21131 30787
rect 1593 30685 1627 30719
rect 4077 30685 4111 30719
rect 8401 30685 8435 30719
rect 9505 30685 9539 30719
rect 9965 30685 9999 30719
rect 12265 30685 12299 30719
rect 13185 30685 13219 30719
rect 13277 30685 13311 30719
rect 13461 30685 13495 30719
rect 13553 30685 13587 30719
rect 13737 30685 13771 30719
rect 14841 30685 14875 30719
rect 14933 30685 14967 30719
rect 15117 30685 15151 30719
rect 15209 30685 15243 30719
rect 17049 30685 17083 30719
rect 19993 30685 20027 30719
rect 20361 30685 20395 30719
rect 20453 30685 20487 30719
rect 23489 30685 23523 30719
rect 23765 30685 23799 30719
rect 25973 30685 26007 30719
rect 27813 30685 27847 30719
rect 11667 30651 11701 30685
rect 6837 30617 6871 30651
rect 10793 30617 10827 30651
rect 11437 30617 11471 30651
rect 16804 30617 16838 30651
rect 18644 30617 18678 30651
rect 20131 30617 20165 30651
rect 20269 30617 20303 30651
rect 21364 30617 21398 30651
rect 25706 30617 25740 30651
rect 27546 30617 27580 30651
rect 3433 30549 3467 30583
rect 4629 30549 4663 30583
rect 5733 30549 5767 30583
rect 7389 30549 7423 30583
rect 8585 30549 8619 30583
rect 10885 30549 10919 30583
rect 12357 30549 12391 30583
rect 12449 30549 12483 30583
rect 14657 30549 14691 30583
rect 15669 30549 15703 30583
rect 19441 30549 19475 30583
rect 22477 30549 22511 30583
rect 24593 30549 24627 30583
rect 26433 30549 26467 30583
rect 28273 30549 28307 30583
rect 6561 30345 6595 30379
rect 17141 30345 17175 30379
rect 25237 30345 25271 30379
rect 27169 30345 27203 30379
rect 5457 30277 5491 30311
rect 7113 30277 7147 30311
rect 8217 30277 8251 30311
rect 10793 30277 10827 30311
rect 10993 30277 11027 30311
rect 17627 30277 17661 30311
rect 19380 30277 19414 30311
rect 27445 30277 27479 30311
rect 27655 30277 27689 30311
rect 4353 30209 4387 30243
rect 9413 30209 9447 30243
rect 10241 30209 10275 30243
rect 12265 30209 12299 30243
rect 12357 30209 12391 30243
rect 12541 30209 12575 30243
rect 12633 30209 12667 30243
rect 13360 30209 13394 30243
rect 16057 30209 16091 30243
rect 17325 30209 17359 30243
rect 17417 30209 17451 30243
rect 17509 30209 17543 30243
rect 20085 30209 20119 30243
rect 20352 30209 20386 30243
rect 22284 30209 22318 30243
rect 24113 30209 24147 30243
rect 26249 30209 26283 30243
rect 27353 30209 27387 30243
rect 27537 30209 27571 30243
rect 6009 30141 6043 30175
rect 8953 30141 8987 30175
rect 13093 30141 13127 30175
rect 16313 30141 16347 30175
rect 17785 30141 17819 30175
rect 19625 30141 19659 30175
rect 22017 30141 22051 30175
rect 23857 30141 23891 30175
rect 26525 30141 26559 30175
rect 27813 30141 27847 30175
rect 7757 30073 7791 30107
rect 11161 30073 11195 30107
rect 14473 30073 14507 30107
rect 4905 30005 4939 30039
rect 9597 30005 9631 30039
rect 10149 30005 10183 30039
rect 10977 30005 11011 30039
rect 12081 30005 12115 30039
rect 14933 30005 14967 30039
rect 18245 30005 18279 30039
rect 21465 30005 21499 30039
rect 23397 30005 23431 30039
rect 28273 30005 28307 30039
rect 5733 29801 5767 29835
rect 7941 29801 7975 29835
rect 8493 29801 8527 29835
rect 9781 29801 9815 29835
rect 26433 29801 26467 29835
rect 9965 29733 9999 29767
rect 13737 29733 13771 29767
rect 14841 29733 14875 29767
rect 14933 29733 14967 29767
rect 17049 29733 17083 29767
rect 4721 29665 4755 29699
rect 11345 29665 11379 29699
rect 15669 29665 15703 29699
rect 17509 29665 17543 29699
rect 1593 29597 1627 29631
rect 7481 29597 7515 29631
rect 10425 29597 10459 29631
rect 10885 29597 10919 29631
rect 11529 29597 11563 29631
rect 11621 29597 11655 29631
rect 11805 29597 11839 29631
rect 11897 29597 11931 29631
rect 12357 29597 12391 29631
rect 14749 29597 14783 29631
rect 15025 29597 15059 29631
rect 17776 29597 17810 29631
rect 20269 29597 20303 29631
rect 20545 29597 20579 29631
rect 22118 29597 22152 29631
rect 22385 29597 22419 29631
rect 22845 29597 22879 29631
rect 23121 29597 23155 29631
rect 24593 29597 24627 29631
rect 24849 29597 24883 29631
rect 27813 29597 27847 29631
rect 6285 29529 6319 29563
rect 9597 29529 9631 29563
rect 12602 29529 12636 29563
rect 15936 29529 15970 29563
rect 27546 29529 27580 29563
rect 5273 29461 5307 29495
rect 6929 29461 6963 29495
rect 9807 29461 9841 29495
rect 10517 29461 10551 29495
rect 10609 29461 10643 29495
rect 15209 29461 15243 29495
rect 18889 29461 18923 29495
rect 21005 29461 21039 29495
rect 25973 29461 26007 29495
rect 28273 29461 28307 29495
rect 6745 29257 6779 29291
rect 7849 29257 7883 29291
rect 8493 29257 8527 29291
rect 27169 29257 27203 29291
rect 10793 29189 10827 29223
rect 10993 29189 11027 29223
rect 17417 29189 17451 29223
rect 17647 29189 17681 29223
rect 24102 29189 24136 29223
rect 27445 29189 27479 29223
rect 10149 29121 10183 29155
rect 12265 29121 12299 29155
rect 12430 29121 12464 29155
rect 12541 29121 12575 29155
rect 12633 29121 12667 29155
rect 13093 29121 13127 29155
rect 13360 29121 13394 29155
rect 15200 29121 15234 29155
rect 17141 29121 17175 29155
rect 17325 29121 17359 29155
rect 17509 29121 17543 29155
rect 18245 29121 18279 29155
rect 18512 29121 18546 29155
rect 21198 29121 21232 29155
rect 23130 29121 23164 29155
rect 27353 29121 27387 29155
rect 27537 29121 27571 29155
rect 27655 29121 27689 29155
rect 27813 29121 27847 29155
rect 7389 29053 7423 29087
rect 14933 29053 14967 29087
rect 17785 29053 17819 29087
rect 21465 29053 21499 29087
rect 23397 29053 23431 29087
rect 23857 29053 23891 29087
rect 25697 29053 25731 29087
rect 25973 29053 26007 29087
rect 6009 28985 6043 29019
rect 8953 28985 8987 29019
rect 11161 28985 11195 29019
rect 20085 28985 20119 29019
rect 22017 28985 22051 29019
rect 9505 28917 9539 28951
rect 10241 28917 10275 28951
rect 10977 28917 11011 28951
rect 12081 28917 12115 28951
rect 14473 28917 14507 28951
rect 16313 28917 16347 28951
rect 19625 28917 19659 28951
rect 25237 28917 25271 28951
rect 28365 28917 28399 28951
rect 6377 28713 6411 28747
rect 8585 28713 8619 28747
rect 10885 28713 10919 28747
rect 11621 28713 11655 28747
rect 11805 28713 11839 28747
rect 14657 28713 14691 28747
rect 6929 28645 6963 28679
rect 7389 28645 7423 28679
rect 7941 28645 7975 28679
rect 9689 28645 9723 28679
rect 17049 28645 17083 28679
rect 21005 28645 21039 28679
rect 15669 28577 15703 28611
rect 20453 28577 20487 28611
rect 23121 28577 23155 28611
rect 24593 28577 24627 28611
rect 1593 28509 1627 28543
rect 10149 28509 10183 28543
rect 12265 28509 12299 28543
rect 12541 28509 12575 28543
rect 12725 28509 12759 28543
rect 13369 28509 13403 28543
rect 13461 28509 13495 28543
rect 13645 28509 13679 28543
rect 13737 28509 13771 28543
rect 14841 28509 14875 28543
rect 14933 28509 14967 28543
rect 15117 28509 15151 28543
rect 15209 28509 15243 28543
rect 18633 28509 18667 28543
rect 18889 28509 18923 28543
rect 22385 28509 22419 28543
rect 22845 28509 22879 28543
rect 26433 28509 26467 28543
rect 10793 28441 10827 28475
rect 11437 28441 11471 28475
rect 11653 28441 11687 28475
rect 15936 28441 15970 28475
rect 22140 28441 22174 28475
rect 24838 28441 24872 28475
rect 26678 28441 26712 28475
rect 12357 28373 12391 28407
rect 13185 28373 13219 28407
rect 17509 28373 17543 28407
rect 19809 28373 19843 28407
rect 20177 28373 20211 28407
rect 20269 28373 20303 28407
rect 25973 28373 26007 28407
rect 27813 28373 27847 28407
rect 28365 28373 28399 28407
rect 7297 28169 7331 28203
rect 10057 28169 10091 28203
rect 10517 28169 10551 28203
rect 11069 28169 11103 28203
rect 13093 28169 13127 28203
rect 14473 28169 14507 28203
rect 18245 28169 18279 28203
rect 7757 28101 7791 28135
rect 8309 28101 8343 28135
rect 12173 28101 12207 28135
rect 12373 28101 12407 28135
rect 15200 28101 15234 28135
rect 17417 28101 17451 28135
rect 17508 28101 17542 28135
rect 19358 28101 19392 28135
rect 21198 28101 21232 28135
rect 25881 28101 25915 28135
rect 26065 28101 26099 28135
rect 13001 28033 13035 28067
rect 13921 28033 13955 28067
rect 14013 28033 14047 28067
rect 14164 28033 14198 28067
rect 14289 28033 14323 28067
rect 14933 28033 14967 28067
rect 17279 28033 17313 28067
rect 17601 28033 17635 28067
rect 17785 28033 17819 28067
rect 21465 28033 21499 28067
rect 23141 28033 23175 28067
rect 24113 28033 24147 28067
rect 27169 28033 27203 28067
rect 27353 28033 27387 28067
rect 27629 28033 27663 28067
rect 28181 28033 28215 28067
rect 28365 28033 28399 28067
rect 8953 27965 8987 27999
rect 13277 27965 13311 27999
rect 13461 27965 13495 27999
rect 17141 27965 17175 27999
rect 19625 27965 19659 27999
rect 23397 27965 23431 27999
rect 23857 27965 23891 27999
rect 25789 27965 25823 27999
rect 27537 27965 27571 27999
rect 25237 27897 25271 27931
rect 27445 27897 27479 27931
rect 1593 27829 1627 27863
rect 9413 27829 9447 27863
rect 12357 27829 12391 27863
rect 12541 27829 12575 27863
rect 16313 27829 16347 27863
rect 20085 27829 20119 27863
rect 22017 27829 22051 27863
rect 26341 27829 26375 27863
rect 28273 27829 28307 27863
rect 8493 27625 8527 27659
rect 10977 27625 11011 27659
rect 12173 27625 12207 27659
rect 13553 27625 13587 27659
rect 15669 27625 15703 27659
rect 25973 27625 26007 27659
rect 27813 27625 27847 27659
rect 9413 27557 9447 27591
rect 9965 27557 9999 27591
rect 11621 27557 11655 27591
rect 12909 27557 12943 27591
rect 15209 27557 15243 27591
rect 21097 27557 21131 27591
rect 10517 27421 10551 27455
rect 14657 27421 14691 27455
rect 14749 27421 14783 27455
rect 14933 27421 14967 27455
rect 15025 27421 15059 27455
rect 17049 27421 17083 27455
rect 18889 27421 18923 27455
rect 20177 27421 20211 27455
rect 20361 27421 20395 27455
rect 20637 27421 20671 27455
rect 22477 27421 22511 27455
rect 22937 27421 22971 27455
rect 23213 27421 23247 27455
rect 24593 27421 24627 27455
rect 26433 27421 26467 27455
rect 12725 27353 12759 27387
rect 13369 27353 13403 27387
rect 16804 27353 16838 27387
rect 18644 27353 18678 27387
rect 20269 27353 20303 27387
rect 20499 27353 20533 27387
rect 22232 27353 22266 27387
rect 24849 27353 24883 27387
rect 26678 27353 26712 27387
rect 8033 27285 8067 27319
rect 13569 27285 13603 27319
rect 13737 27285 13771 27319
rect 17509 27285 17543 27319
rect 19533 27285 19567 27319
rect 19993 27285 20027 27319
rect 28365 27285 28399 27319
rect 9505 27081 9539 27115
rect 9965 27081 9999 27115
rect 10609 27081 10643 27115
rect 11161 27081 11195 27115
rect 12173 27081 12207 27115
rect 14013 27081 14047 27115
rect 16313 27081 16347 27115
rect 17785 27081 17819 27115
rect 23857 27081 23891 27115
rect 25697 27081 25731 27115
rect 14165 27013 14199 27047
rect 14381 27013 14415 27047
rect 27169 27013 27203 27047
rect 12817 26945 12851 26979
rect 13461 26945 13495 26979
rect 14841 26945 14875 26979
rect 14933 26945 14967 26979
rect 15301 26945 15335 26979
rect 15853 26945 15887 26979
rect 16129 26945 16163 26979
rect 17312 26945 17346 26979
rect 17601 26945 17635 26979
rect 18245 26945 18279 26979
rect 18512 26945 18546 26979
rect 20352 26945 20386 26979
rect 22284 26945 22318 26979
rect 24981 26945 25015 26979
rect 25881 26945 25915 26979
rect 26157 26945 26191 26979
rect 27353 26945 27387 26979
rect 27629 26945 27663 26979
rect 28365 26945 28399 26979
rect 15117 26877 15151 26911
rect 17417 26877 17451 26911
rect 20085 26877 20119 26911
rect 22017 26877 22051 26911
rect 25237 26877 25271 26911
rect 25973 26877 26007 26911
rect 27445 26877 27479 26911
rect 15945 26809 15979 26843
rect 16037 26809 16071 26843
rect 17509 26809 17543 26843
rect 26065 26809 26099 26843
rect 27537 26809 27571 26843
rect 8953 26741 8987 26775
rect 13369 26741 13403 26775
rect 14197 26741 14231 26775
rect 19625 26741 19659 26775
rect 21465 26741 21499 26775
rect 23397 26741 23431 26775
rect 28181 26741 28215 26775
rect 10425 26537 10459 26571
rect 11437 26537 11471 26571
rect 12081 26537 12115 26571
rect 14841 26537 14875 26571
rect 16037 26537 16071 26571
rect 27813 26537 27847 26571
rect 28365 26537 28399 26571
rect 10977 26469 11011 26503
rect 15025 26469 15059 26503
rect 17049 26469 17083 26503
rect 18889 26469 18923 26503
rect 20913 26469 20947 26503
rect 23213 26469 23247 26503
rect 24593 26469 24627 26503
rect 12633 26401 12667 26435
rect 17509 26401 17543 26435
rect 19533 26401 19567 26435
rect 1593 26333 1627 26367
rect 9873 26333 9907 26367
rect 13093 26333 13127 26367
rect 15475 26333 15509 26367
rect 15577 26333 15611 26367
rect 15761 26333 15795 26367
rect 15853 26333 15887 26367
rect 16497 26333 16531 26367
rect 16589 26333 16623 26367
rect 16773 26333 16807 26367
rect 16865 26333 16899 26367
rect 19800 26333 19834 26367
rect 22753 26333 22787 26367
rect 23397 26333 23431 26367
rect 23489 26333 23523 26367
rect 23857 26333 23891 26367
rect 25973 26333 26007 26367
rect 26433 26333 26467 26367
rect 14657 26265 14691 26299
rect 14857 26265 14891 26299
rect 17776 26265 17810 26299
rect 22508 26265 22542 26299
rect 23581 26265 23615 26299
rect 23699 26265 23733 26299
rect 25728 26265 25762 26299
rect 26678 26265 26712 26299
rect 13737 26197 13771 26231
rect 21373 26197 21407 26231
rect 10425 25993 10459 26027
rect 13001 25993 13035 26027
rect 15945 25993 15979 26027
rect 25697 25993 25731 26027
rect 28273 25993 28307 26027
rect 15485 25925 15519 25959
rect 16113 25925 16147 25959
rect 16313 25925 16347 25959
rect 17233 25925 17267 25959
rect 18512 25925 18546 25959
rect 21198 25925 21232 25959
rect 24970 25925 25004 25959
rect 14657 25857 14691 25891
rect 15301 25857 15335 25891
rect 17417 25857 17451 25891
rect 17509 25857 17543 25891
rect 17693 25857 17727 25891
rect 17785 25857 17819 25891
rect 18245 25857 18279 25891
rect 21465 25857 21499 25891
rect 22273 25857 22307 25891
rect 25237 25857 25271 25891
rect 25881 25857 25915 25891
rect 26157 25857 26191 25891
rect 27353 25857 27387 25891
rect 27445 25857 27479 25891
rect 27629 25857 27663 25891
rect 27721 25857 27755 25891
rect 28181 25857 28215 25891
rect 28365 25857 28399 25891
rect 22017 25789 22051 25823
rect 26065 25789 26099 25823
rect 11161 25721 11195 25755
rect 14197 25721 14231 25755
rect 19625 25721 19659 25755
rect 23857 25721 23891 25755
rect 25973 25721 26007 25755
rect 27169 25721 27203 25755
rect 1593 25653 1627 25687
rect 11989 25653 12023 25687
rect 12541 25653 12575 25687
rect 13553 25653 13587 25687
rect 16129 25653 16163 25687
rect 20085 25653 20119 25687
rect 23397 25653 23431 25687
rect 12081 25449 12115 25483
rect 13093 25449 13127 25483
rect 16497 25449 16531 25483
rect 16681 25449 16715 25483
rect 18337 25449 18371 25483
rect 19441 25449 19475 25483
rect 26985 25449 27019 25483
rect 15761 25381 15795 25415
rect 17325 25381 17359 25415
rect 23489 25381 23523 25415
rect 17509 25245 17543 25279
rect 17601 25245 17635 25279
rect 17785 25245 17819 25279
rect 17877 25245 17911 25279
rect 18521 25245 18555 25279
rect 18613 25245 18647 25279
rect 18797 25245 18831 25279
rect 18889 25245 18923 25279
rect 20554 25245 20588 25279
rect 20821 25245 20855 25279
rect 22661 25245 22695 25279
rect 23305 25245 23339 25279
rect 23397 25245 23431 25279
rect 23581 25245 23615 25279
rect 25973 25245 26007 25279
rect 26433 25245 26467 25279
rect 26525 25245 26559 25279
rect 26709 25245 26743 25279
rect 26801 25245 26835 25279
rect 27629 25245 27663 25279
rect 27905 25245 27939 25279
rect 15945 25177 15979 25211
rect 16649 25177 16683 25211
rect 16865 25177 16899 25211
rect 22416 25177 22450 25211
rect 25706 25177 25740 25211
rect 13737 25109 13771 25143
rect 14749 25109 14783 25143
rect 15209 25109 15243 25143
rect 21281 25109 21315 25143
rect 23121 25109 23155 25143
rect 24593 25109 24627 25143
rect 27445 25109 27479 25143
rect 27813 25109 27847 25143
rect 18245 24905 18279 24939
rect 21465 24905 21499 24939
rect 26249 24905 26283 24939
rect 14013 24837 14047 24871
rect 16221 24837 16255 24871
rect 17477 24837 17511 24871
rect 17693 24837 17727 24871
rect 20330 24837 20364 24871
rect 27321 24837 27355 24871
rect 27537 24837 27571 24871
rect 13369 24769 13403 24803
rect 15025 24769 15059 24803
rect 18153 24769 18187 24803
rect 18613 24769 18647 24803
rect 19073 24769 19107 24803
rect 19257 24769 19291 24803
rect 19349 24769 19383 24803
rect 19533 24769 19567 24803
rect 19635 24769 19669 24803
rect 20085 24769 20119 24803
rect 23130 24769 23164 24803
rect 23397 24769 23431 24803
rect 24970 24769 25004 24803
rect 25237 24769 25271 24803
rect 25697 24769 25731 24803
rect 25789 24769 25823 24803
rect 25900 24769 25934 24803
rect 26065 24769 26099 24803
rect 27997 24769 28031 24803
rect 18429 24701 18463 24735
rect 14565 24633 14599 24667
rect 17325 24633 17359 24667
rect 15669 24565 15703 24599
rect 17509 24565 17543 24599
rect 22017 24565 22051 24599
rect 23857 24565 23891 24599
rect 27169 24565 27203 24599
rect 27353 24565 27387 24599
rect 27997 24565 28031 24599
rect 15393 24361 15427 24395
rect 17877 24361 17911 24395
rect 18705 24361 18739 24395
rect 19625 24361 19659 24395
rect 19809 24361 19843 24395
rect 23673 24361 23707 24395
rect 24593 24361 24627 24395
rect 26617 24361 26651 24395
rect 26801 24361 26835 24395
rect 17049 24293 17083 24327
rect 17693 24293 17727 24327
rect 18889 24293 18923 24327
rect 20269 24293 20303 24327
rect 22661 24293 22695 24327
rect 28089 24293 28123 24327
rect 14841 24225 14875 24259
rect 1593 24157 1627 24191
rect 15945 24157 15979 24191
rect 16497 24157 16531 24191
rect 20445 24157 20479 24191
rect 20537 24157 20571 24191
rect 20729 24157 20763 24191
rect 20821 24157 20855 24191
rect 21281 24157 21315 24191
rect 23121 24157 23155 24191
rect 23213 24157 23247 24191
rect 23397 24157 23431 24191
rect 23489 24157 23523 24191
rect 25973 24157 26007 24191
rect 27445 24157 27479 24191
rect 18035 24089 18069 24123
rect 18521 24089 18555 24123
rect 19441 24089 19475 24123
rect 21526 24089 21560 24123
rect 25706 24089 25740 24123
rect 26433 24089 26467 24123
rect 27261 24089 27295 24123
rect 28273 24089 28307 24123
rect 17851 24021 17885 24055
rect 18721 24021 18755 24055
rect 19651 24021 19685 24055
rect 26633 24021 26667 24055
rect 15209 23817 15243 23851
rect 17233 23817 17267 23851
rect 25697 23817 25731 23851
rect 17877 23749 17911 23783
rect 18429 23749 18463 23783
rect 18613 23749 18647 23783
rect 19317 23749 19351 23783
rect 19533 23749 19567 23783
rect 20085 23749 20119 23783
rect 24992 23749 25026 23783
rect 16221 23681 16255 23715
rect 19993 23681 20027 23715
rect 20269 23681 20303 23715
rect 20453 23681 20487 23715
rect 21097 23681 21131 23715
rect 21189 23681 21223 23715
rect 21358 23681 21392 23715
rect 21465 23681 21499 23715
rect 22273 23681 22307 23715
rect 25237 23681 25271 23715
rect 25881 23681 25915 23715
rect 26065 23681 26099 23715
rect 26617 23681 26651 23715
rect 27721 23681 27755 23715
rect 28365 23681 28399 23715
rect 15761 23613 15795 23647
rect 22017 23613 22051 23647
rect 19165 23545 19199 23579
rect 20913 23545 20947 23579
rect 1593 23477 1627 23511
rect 19349 23477 19383 23511
rect 23397 23477 23431 23511
rect 23857 23477 23891 23511
rect 27537 23477 27571 23511
rect 16221 23273 16255 23307
rect 16773 23273 16807 23307
rect 17877 23273 17911 23307
rect 19717 23273 19751 23307
rect 20536 23273 20570 23307
rect 20729 23273 20763 23307
rect 24777 23273 24811 23307
rect 25605 23273 25639 23307
rect 27721 23273 27755 23307
rect 18337 23205 18371 23239
rect 22201 23205 22235 23239
rect 25789 23205 25823 23239
rect 26433 23205 26467 23239
rect 21189 23137 21223 23171
rect 21373 23069 21407 23103
rect 21465 23069 21499 23103
rect 21649 23069 21683 23103
rect 21741 23069 21775 23103
rect 23581 23069 23615 23103
rect 26249 23069 26283 23103
rect 26433 23069 26467 23103
rect 27077 23069 27111 23103
rect 28365 23069 28399 23103
rect 19901 23001 19935 23035
rect 20361 23001 20395 23035
rect 23336 23001 23370 23035
rect 24593 23001 24627 23035
rect 25421 23001 25455 23035
rect 25621 23001 25655 23035
rect 17325 22933 17359 22967
rect 19533 22933 19567 22967
rect 19701 22933 19735 22967
rect 20561 22933 20595 22967
rect 24803 22933 24837 22967
rect 24961 22933 24995 22967
rect 26893 22933 26927 22967
rect 16865 22729 16899 22763
rect 18061 22729 18095 22763
rect 19073 22729 19107 22763
rect 19809 22729 19843 22763
rect 21297 22729 21331 22763
rect 21465 22729 21499 22763
rect 24041 22729 24075 22763
rect 24209 22729 24243 22763
rect 25037 22729 25071 22763
rect 25789 22729 25823 22763
rect 28181 22729 28215 22763
rect 20437 22661 20471 22695
rect 20637 22661 20671 22695
rect 21097 22661 21131 22695
rect 23489 22661 23523 22695
rect 24409 22661 24443 22695
rect 25237 22661 25271 22695
rect 22007 22599 22041 22633
rect 22109 22593 22143 22627
rect 22301 22593 22335 22627
rect 22393 22593 22427 22627
rect 23029 22593 23063 22627
rect 23213 22593 23247 22627
rect 23581 22593 23615 22627
rect 25973 22593 26007 22627
rect 27721 22593 27755 22627
rect 28365 22593 28399 22627
rect 26617 22525 26651 22559
rect 20269 22457 20303 22491
rect 24869 22457 24903 22491
rect 1593 22389 1627 22423
rect 17509 22389 17543 22423
rect 20453 22389 20487 22423
rect 21281 22389 21315 22423
rect 22569 22389 22603 22423
rect 24225 22389 24259 22423
rect 25053 22389 25087 22423
rect 18889 22185 18923 22219
rect 22017 22185 22051 22219
rect 22845 22185 22879 22219
rect 23029 22185 23063 22219
rect 23673 22185 23707 22219
rect 25789 22185 25823 22219
rect 27077 22185 27111 22219
rect 27537 22185 27571 22219
rect 19717 22117 19751 22151
rect 20177 22117 20211 22151
rect 21097 22117 21131 22151
rect 23489 22117 23523 22151
rect 26433 22117 26467 22151
rect 18337 22049 18371 22083
rect 17785 21981 17819 22015
rect 21281 21981 21315 22015
rect 24777 21981 24811 22015
rect 27721 21981 27755 22015
rect 28365 21981 28399 22015
rect 22001 21913 22035 21947
rect 22201 21913 22235 21947
rect 22661 21913 22695 21947
rect 23857 21913 23891 21947
rect 21833 21845 21867 21879
rect 22871 21845 22905 21879
rect 23647 21845 23681 21879
rect 24685 21845 24719 21879
rect 19349 21641 19383 21675
rect 22109 21641 22143 21675
rect 23857 21641 23891 21675
rect 26433 21641 26467 21675
rect 22261 21573 22295 21607
rect 22477 21573 22511 21607
rect 23305 21573 23339 21607
rect 25145 21573 25179 21607
rect 25697 21573 25731 21607
rect 23075 21539 23109 21573
rect 23765 21505 23799 21539
rect 24409 21505 24443 21539
rect 26617 21505 26651 21539
rect 27169 21505 27203 21539
rect 1593 21437 1627 21471
rect 19809 21369 19843 21403
rect 20729 21369 20763 21403
rect 18797 21301 18831 21335
rect 21373 21301 21407 21335
rect 22293 21301 22327 21335
rect 22937 21301 22971 21335
rect 23121 21301 23155 21335
rect 28365 21301 28399 21335
rect 19901 21097 19935 21131
rect 20453 21097 20487 21131
rect 20913 21097 20947 21131
rect 21465 21097 21499 21131
rect 23121 21097 23155 21131
rect 25145 21097 25179 21131
rect 25789 21097 25823 21131
rect 26249 21097 26283 21131
rect 28365 21097 28399 21131
rect 23765 21029 23799 21063
rect 24593 21029 24627 21063
rect 27721 21029 27755 21063
rect 27077 20961 27111 20995
rect 22385 20893 22419 20927
rect 23213 20893 23247 20927
rect 22569 20825 22603 20859
rect 19993 20553 20027 20587
rect 21005 20553 21039 20587
rect 22109 20553 22143 20587
rect 22661 20553 22695 20587
rect 23213 20553 23247 20587
rect 26065 20553 26099 20587
rect 27261 20553 27295 20587
rect 28181 20553 28215 20587
rect 23857 20485 23891 20519
rect 20545 20417 20579 20451
rect 24317 20417 24351 20451
rect 28365 20417 28399 20451
rect 1593 20213 1627 20247
rect 24961 20213 24995 20247
rect 25513 20213 25547 20247
rect 26617 20213 26651 20247
rect 20637 20009 20671 20043
rect 21649 20009 21683 20043
rect 22293 20009 22327 20043
rect 23121 20009 23155 20043
rect 23673 20009 23707 20043
rect 25145 20009 25179 20043
rect 27169 20009 27203 20043
rect 27721 20009 27755 20043
rect 24593 19941 24627 19975
rect 21189 19873 21223 19907
rect 1593 19805 1627 19839
rect 28365 19805 28399 19839
rect 25789 19669 25823 19703
rect 26341 19669 26375 19703
rect 22017 19465 22051 19499
rect 22845 19465 22879 19499
rect 23489 19465 23523 19499
rect 26157 19465 26191 19499
rect 27721 19465 27755 19499
rect 25145 19397 25179 19431
rect 24041 19261 24075 19295
rect 24593 19193 24627 19227
rect 28365 19125 28399 19159
rect 23581 18921 23615 18955
rect 24869 18921 24903 18955
rect 26249 18853 26283 18887
rect 28089 18785 28123 18819
rect 28365 18717 28399 18751
rect 22385 18581 22419 18615
rect 23029 18581 23063 18615
rect 25421 18581 25455 18615
rect 26893 18581 26927 18615
rect 25881 18377 25915 18411
rect 26525 18377 26559 18411
rect 27721 18377 27755 18411
rect 23765 18309 23799 18343
rect 27169 18309 27203 18343
rect 28365 18309 28399 18343
rect 1593 18037 1627 18071
rect 24869 18037 24903 18071
rect 25421 18037 25455 18071
rect 24593 17833 24627 17867
rect 25605 17833 25639 17867
rect 26249 17833 26283 17867
rect 26985 17833 27019 17867
rect 27721 17833 27755 17867
rect 1593 17629 1627 17663
rect 28365 17629 28399 17663
rect 25053 17289 25087 17323
rect 25513 17289 25547 17323
rect 27169 17289 27203 17323
rect 26065 17221 26099 17255
rect 28365 16949 28399 16983
rect 26249 16745 26283 16779
rect 27813 16745 27847 16779
rect 26985 16677 27019 16711
rect 27629 16201 27663 16235
rect 1593 15997 1627 16031
rect 28365 15861 28399 15895
rect 1593 15453 1627 15487
rect 28365 14841 28399 14875
rect 1593 14365 1627 14399
rect 28365 13685 28399 13719
rect 1593 13277 1627 13311
rect 28365 13277 28399 13311
rect 1593 12189 1627 12223
rect 1593 11509 1627 11543
rect 28365 11509 28399 11543
rect 28365 11101 28399 11135
rect 1593 10013 1627 10047
rect 28365 9401 28399 9435
rect 1593 9333 1627 9367
rect 28365 9061 28399 9095
rect 1593 7837 1627 7871
rect 28365 7837 28399 7871
rect 1593 7157 1627 7191
rect 28365 6749 28399 6783
rect 1593 6069 1627 6103
rect 28365 5661 28399 5695
rect 1593 5117 1627 5151
rect 28365 4981 28399 5015
rect 1593 3893 1627 3927
rect 28365 3621 28399 3655
rect 1593 3485 1627 3519
rect 28365 2805 28399 2839
<< metal1 >>
rect 11790 32172 11796 32224
rect 11848 32212 11854 32224
rect 14918 32212 14924 32224
rect 11848 32184 14924 32212
rect 11848 32172 11854 32184
rect 14918 32172 14924 32184
rect 14976 32172 14982 32224
rect 20254 32036 20260 32088
rect 20312 32076 20318 32088
rect 21542 32076 21548 32088
rect 20312 32048 21548 32076
rect 20312 32036 20318 32048
rect 21542 32036 21548 32048
rect 21600 32036 21606 32088
rect 8386 31900 8392 31952
rect 8444 31940 8450 31952
rect 26878 31940 26884 31952
rect 8444 31912 26884 31940
rect 8444 31900 8450 31912
rect 26878 31900 26884 31912
rect 26936 31900 26942 31952
rect 13998 31832 14004 31884
rect 14056 31872 14062 31884
rect 18690 31872 18696 31884
rect 14056 31844 18696 31872
rect 14056 31832 14062 31844
rect 18690 31832 18696 31844
rect 18748 31832 18754 31884
rect 11698 31764 11704 31816
rect 11756 31804 11762 31816
rect 11756 31776 19334 31804
rect 11756 31764 11762 31776
rect 8570 31696 8576 31748
rect 8628 31736 8634 31748
rect 13814 31736 13820 31748
rect 8628 31708 13820 31736
rect 8628 31696 8634 31708
rect 13814 31696 13820 31708
rect 13872 31696 13878 31748
rect 16574 31696 16580 31748
rect 16632 31736 16638 31748
rect 18782 31736 18788 31748
rect 16632 31708 18788 31736
rect 16632 31696 16638 31708
rect 18782 31696 18788 31708
rect 18840 31696 18846 31748
rect 13722 31628 13728 31680
rect 13780 31668 13786 31680
rect 18506 31668 18512 31680
rect 13780 31640 18512 31668
rect 13780 31628 13786 31640
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 19306 31668 19334 31776
rect 19978 31696 19984 31748
rect 20036 31736 20042 31748
rect 21634 31736 21640 31748
rect 20036 31708 21640 31736
rect 20036 31696 20042 31708
rect 21634 31696 21640 31708
rect 21692 31696 21698 31748
rect 22646 31668 22652 31680
rect 19306 31640 22652 31668
rect 22646 31628 22652 31640
rect 22704 31628 22710 31680
rect 22738 31628 22744 31680
rect 22796 31668 22802 31680
rect 28350 31668 28356 31680
rect 22796 31640 28356 31668
rect 22796 31628 22802 31640
rect 28350 31628 28356 31640
rect 28408 31628 28414 31680
rect 1104 31578 29048 31600
rect 1104 31526 7896 31578
rect 7948 31526 7960 31578
rect 8012 31526 8024 31578
rect 8076 31526 8088 31578
rect 8140 31526 8152 31578
rect 8204 31526 14842 31578
rect 14894 31526 14906 31578
rect 14958 31526 14970 31578
rect 15022 31526 15034 31578
rect 15086 31526 15098 31578
rect 15150 31526 21788 31578
rect 21840 31526 21852 31578
rect 21904 31526 21916 31578
rect 21968 31526 21980 31578
rect 22032 31526 22044 31578
rect 22096 31526 28734 31578
rect 28786 31526 28798 31578
rect 28850 31526 28862 31578
rect 28914 31526 28926 31578
rect 28978 31526 28990 31578
rect 29042 31526 29048 31578
rect 1104 31504 29048 31526
rect 1670 31424 1676 31476
rect 1728 31464 1734 31476
rect 1857 31467 1915 31473
rect 1857 31464 1869 31467
rect 1728 31436 1869 31464
rect 1728 31424 1734 31436
rect 1857 31433 1869 31436
rect 1903 31433 1915 31467
rect 1857 31427 1915 31433
rect 4982 31424 4988 31476
rect 5040 31464 5046 31476
rect 5169 31467 5227 31473
rect 5169 31464 5181 31467
rect 5040 31436 5181 31464
rect 5040 31424 5046 31436
rect 5169 31433 5181 31436
rect 5215 31433 5227 31467
rect 5169 31427 5227 31433
rect 8294 31424 8300 31476
rect 8352 31464 8358 31476
rect 9217 31467 9275 31473
rect 9217 31464 9229 31467
rect 8352 31436 9229 31464
rect 8352 31424 8358 31436
rect 9217 31433 9229 31436
rect 9263 31433 9275 31467
rect 9217 31427 9275 31433
rect 10229 31467 10287 31473
rect 10229 31433 10241 31467
rect 10275 31464 10287 31467
rect 11606 31464 11612 31476
rect 10275 31436 11612 31464
rect 10275 31433 10287 31436
rect 10229 31427 10287 31433
rect 11606 31424 11612 31436
rect 11664 31424 11670 31476
rect 11790 31464 11796 31476
rect 11751 31436 11796 31464
rect 11790 31424 11796 31436
rect 11848 31424 11854 31476
rect 13449 31467 13507 31473
rect 12452 31436 12848 31464
rect 8478 31396 8484 31408
rect 2056 31368 8484 31396
rect 2056 31337 2084 31368
rect 8478 31356 8484 31368
rect 8536 31356 8542 31408
rect 9858 31356 9864 31408
rect 9916 31396 9922 31408
rect 12452 31405 12480 31436
rect 12437 31399 12495 31405
rect 9916 31368 12388 31396
rect 9916 31356 9922 31368
rect 2041 31331 2099 31337
rect 2041 31297 2053 31331
rect 2087 31297 2099 31331
rect 2041 31291 2099 31297
rect 3878 31288 3884 31340
rect 3936 31328 3942 31340
rect 3973 31331 4031 31337
rect 3973 31328 3985 31331
rect 3936 31300 3985 31328
rect 3936 31288 3942 31300
rect 3973 31297 3985 31300
rect 4019 31297 4031 31331
rect 5350 31328 5356 31340
rect 5311 31300 5356 31328
rect 3973 31291 4031 31297
rect 5350 31288 5356 31300
rect 5408 31288 5414 31340
rect 7101 31331 7159 31337
rect 7101 31297 7113 31331
rect 7147 31328 7159 31331
rect 7190 31328 7196 31340
rect 7147 31300 7196 31328
rect 7147 31297 7159 31300
rect 7101 31291 7159 31297
rect 7190 31288 7196 31300
rect 7248 31288 7254 31340
rect 8570 31328 8576 31340
rect 8531 31300 8576 31328
rect 8570 31288 8576 31300
rect 8628 31288 8634 31340
rect 9401 31331 9459 31337
rect 9401 31297 9413 31331
rect 9447 31297 9459 31331
rect 9401 31291 9459 31297
rect 10413 31331 10471 31337
rect 10413 31297 10425 31331
rect 10459 31297 10471 31331
rect 10413 31291 10471 31297
rect 566 31220 572 31272
rect 624 31260 630 31272
rect 2501 31263 2559 31269
rect 2501 31260 2513 31263
rect 624 31232 2513 31260
rect 624 31220 630 31232
rect 2501 31229 2513 31232
rect 2547 31229 2559 31263
rect 2501 31223 2559 31229
rect 9416 31192 9444 31291
rect 10428 31260 10456 31291
rect 11146 31288 11152 31340
rect 11204 31328 11210 31340
rect 11974 31328 11980 31340
rect 11204 31300 11249 31328
rect 11935 31300 11980 31328
rect 11204 31288 11210 31300
rect 11974 31288 11980 31300
rect 12032 31288 12038 31340
rect 12360 31328 12388 31368
rect 12437 31365 12449 31399
rect 12483 31365 12495 31399
rect 12820 31396 12848 31436
rect 13449 31433 13461 31467
rect 13495 31464 13507 31467
rect 13538 31464 13544 31476
rect 13495 31436 13544 31464
rect 13495 31433 13507 31436
rect 13449 31427 13507 31433
rect 13538 31424 13544 31436
rect 13596 31424 13602 31476
rect 14921 31467 14979 31473
rect 14921 31464 14933 31467
rect 13786 31436 14933 31464
rect 13786 31396 13814 31436
rect 14921 31433 14933 31436
rect 14967 31464 14979 31467
rect 19150 31464 19156 31476
rect 14967 31436 19156 31464
rect 14967 31433 14979 31436
rect 14921 31427 14979 31433
rect 19150 31424 19156 31436
rect 19208 31424 19214 31476
rect 23198 31464 23204 31476
rect 19628 31436 23204 31464
rect 12437 31359 12495 31365
rect 12667 31365 12725 31371
rect 12820 31368 13814 31396
rect 12667 31331 12679 31365
rect 12713 31331 12725 31365
rect 15562 31356 15568 31408
rect 15620 31396 15626 31408
rect 17764 31399 17822 31405
rect 15620 31368 17540 31396
rect 15620 31356 15626 31368
rect 12667 31328 12725 31331
rect 13262 31328 13268 31340
rect 12360 31325 12725 31328
rect 12360 31300 12710 31325
rect 13223 31300 13268 31328
rect 13262 31288 13268 31300
rect 13320 31288 13326 31340
rect 13354 31288 13360 31340
rect 13412 31328 13418 31340
rect 13648 31328 13860 31332
rect 14461 31331 14519 31337
rect 13412 31300 13457 31328
rect 13648 31304 14412 31328
rect 13412 31288 13418 31300
rect 13648 31260 13676 31304
rect 13832 31300 14412 31304
rect 10428 31232 13676 31260
rect 13722 31220 13728 31272
rect 13780 31260 13786 31272
rect 13780 31232 13825 31260
rect 13780 31220 13786 31232
rect 14277 31195 14335 31201
rect 14277 31192 14289 31195
rect 9416 31164 14289 31192
rect 14277 31161 14289 31164
rect 14323 31161 14335 31195
rect 14277 31155 14335 31161
rect 3421 31127 3479 31133
rect 3421 31093 3433 31127
rect 3467 31124 3479 31127
rect 5810 31124 5816 31136
rect 3467 31096 5816 31124
rect 3467 31093 3479 31096
rect 3421 31087 3479 31093
rect 5810 31084 5816 31096
rect 5868 31084 5874 31136
rect 5997 31127 6055 31133
rect 5997 31093 6009 31127
rect 6043 31124 6055 31127
rect 6178 31124 6184 31136
rect 6043 31096 6184 31124
rect 6043 31093 6055 31096
rect 5997 31087 6055 31093
rect 6178 31084 6184 31096
rect 6236 31084 6242 31136
rect 6641 31127 6699 31133
rect 6641 31093 6653 31127
rect 6687 31124 6699 31127
rect 7650 31124 7656 31136
rect 6687 31096 7656 31124
rect 6687 31093 6699 31096
rect 6641 31087 6699 31093
rect 7650 31084 7656 31096
rect 7708 31084 7714 31136
rect 7929 31127 7987 31133
rect 7929 31093 7941 31127
rect 7975 31124 7987 31127
rect 10134 31124 10140 31136
rect 7975 31096 10140 31124
rect 7975 31093 7987 31096
rect 7929 31087 7987 31093
rect 10134 31084 10140 31096
rect 10192 31084 10198 31136
rect 10965 31127 11023 31133
rect 10965 31093 10977 31127
rect 11011 31124 11023 31127
rect 12158 31124 12164 31136
rect 11011 31096 12164 31124
rect 11011 31093 11023 31096
rect 10965 31087 11023 31093
rect 12158 31084 12164 31096
rect 12216 31084 12222 31136
rect 12621 31127 12679 31133
rect 12621 31093 12633 31127
rect 12667 31124 12679 31127
rect 12710 31124 12716 31136
rect 12667 31096 12716 31124
rect 12667 31093 12679 31096
rect 12621 31087 12679 31093
rect 12710 31084 12716 31096
rect 12768 31084 12774 31136
rect 12805 31127 12863 31133
rect 12805 31093 12817 31127
rect 12851 31124 12863 31127
rect 13906 31124 13912 31136
rect 12851 31096 13912 31124
rect 12851 31093 12863 31096
rect 12805 31087 12863 31093
rect 13906 31084 13912 31096
rect 13964 31084 13970 31136
rect 14384 31124 14412 31300
rect 14461 31297 14473 31331
rect 14507 31328 14519 31331
rect 15470 31328 15476 31340
rect 14507 31300 15476 31328
rect 14507 31297 14519 31300
rect 14461 31291 14519 31297
rect 15470 31288 15476 31300
rect 15528 31288 15534 31340
rect 16045 31331 16103 31337
rect 16045 31297 16057 31331
rect 16091 31328 16103 31331
rect 16758 31328 16764 31340
rect 16091 31300 16764 31328
rect 16091 31297 16103 31300
rect 16045 31291 16103 31297
rect 16758 31288 16764 31300
rect 16816 31288 16822 31340
rect 17034 31328 17040 31340
rect 16995 31300 17040 31328
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 17512 31337 17540 31368
rect 17764 31365 17776 31399
rect 17810 31396 17822 31399
rect 18138 31396 18144 31408
rect 17810 31368 18144 31396
rect 17810 31365 17822 31368
rect 17764 31359 17822 31365
rect 18138 31356 18144 31368
rect 18196 31356 18202 31408
rect 17497 31331 17555 31337
rect 17497 31297 17509 31331
rect 17543 31328 17555 31331
rect 18874 31328 18880 31340
rect 17543 31300 18880 31328
rect 17543 31297 17555 31300
rect 17497 31291 17555 31297
rect 18874 31288 18880 31300
rect 18932 31328 18938 31340
rect 19518 31328 19524 31340
rect 18932 31300 19524 31328
rect 18932 31288 18938 31300
rect 19518 31288 19524 31300
rect 19576 31288 19582 31340
rect 19628 31337 19656 31436
rect 23198 31424 23204 31436
rect 23256 31424 23262 31476
rect 28166 31464 28172 31476
rect 28127 31436 28172 31464
rect 28166 31424 28172 31436
rect 28224 31424 28230 31476
rect 20622 31356 20628 31408
rect 20680 31396 20686 31408
rect 21082 31396 21088 31408
rect 20680 31368 21088 31396
rect 20680 31356 20686 31368
rect 21082 31356 21088 31368
rect 21140 31356 21146 31408
rect 21174 31356 21180 31408
rect 21232 31405 21238 31408
rect 21232 31396 21244 31405
rect 21232 31368 21277 31396
rect 21232 31359 21244 31368
rect 21232 31356 21238 31359
rect 21358 31356 21364 31408
rect 21416 31396 21422 31408
rect 21416 31368 26648 31396
rect 21416 31356 21422 31368
rect 19613 31331 19671 31337
rect 19613 31297 19625 31331
rect 19659 31297 19671 31331
rect 20806 31328 20812 31340
rect 19613 31291 19671 31297
rect 20456 31300 20812 31328
rect 16301 31263 16359 31269
rect 16301 31229 16313 31263
rect 16347 31260 16359 31263
rect 16482 31260 16488 31272
rect 16347 31232 16488 31260
rect 16347 31229 16359 31232
rect 16301 31223 16359 31229
rect 16482 31220 16488 31232
rect 16540 31220 16546 31272
rect 18506 31220 18512 31272
rect 18564 31260 18570 31272
rect 20456 31260 20484 31300
rect 20806 31288 20812 31300
rect 20864 31288 20870 31340
rect 20898 31288 20904 31340
rect 20956 31328 20962 31340
rect 20956 31300 21496 31328
rect 20956 31288 20962 31300
rect 21468 31269 21496 31300
rect 21542 31288 21548 31340
rect 21600 31328 21606 31340
rect 24854 31337 24860 31340
rect 23118 31331 23176 31337
rect 23118 31328 23130 31331
rect 21600 31300 23130 31328
rect 21600 31288 21606 31300
rect 23118 31297 23130 31300
rect 23164 31297 23176 31331
rect 23118 31291 23176 31297
rect 24848 31291 24860 31337
rect 24912 31328 24918 31340
rect 26620 31337 26648 31368
rect 26605 31331 26663 31337
rect 24912 31300 24948 31328
rect 24854 31288 24860 31291
rect 24912 31288 24918 31300
rect 26605 31297 26617 31331
rect 26651 31297 26663 31331
rect 26605 31291 26663 31297
rect 26694 31288 26700 31340
rect 26752 31328 26758 31340
rect 27157 31331 27215 31337
rect 27157 31328 27169 31331
rect 26752 31300 27169 31328
rect 26752 31288 26758 31300
rect 27157 31297 27169 31300
rect 27203 31297 27215 31331
rect 27157 31291 27215 31297
rect 27246 31288 27252 31340
rect 27304 31328 27310 31340
rect 27433 31331 27491 31337
rect 27304 31300 27349 31328
rect 27304 31288 27310 31300
rect 27433 31297 27445 31331
rect 27479 31297 27491 31331
rect 27433 31291 27491 31297
rect 27525 31331 27583 31337
rect 27525 31297 27537 31331
rect 27571 31328 27583 31331
rect 27890 31328 27896 31340
rect 27571 31300 27896 31328
rect 27571 31297 27583 31300
rect 27525 31291 27583 31297
rect 18564 31232 20484 31260
rect 21453 31263 21511 31269
rect 18564 31220 18570 31232
rect 21453 31229 21465 31263
rect 21499 31260 21511 31263
rect 22094 31260 22100 31272
rect 21499 31232 22100 31260
rect 21499 31229 21511 31232
rect 21453 31223 21511 31229
rect 22094 31220 22100 31232
rect 22152 31220 22158 31272
rect 23385 31263 23443 31269
rect 23385 31229 23397 31263
rect 23431 31260 23443 31263
rect 23934 31260 23940 31272
rect 23431 31232 23940 31260
rect 23431 31229 23443 31232
rect 23385 31223 23443 31229
rect 23934 31220 23940 31232
rect 23992 31220 23998 31272
rect 24486 31220 24492 31272
rect 24544 31260 24550 31272
rect 24581 31263 24639 31269
rect 24581 31260 24593 31263
rect 24544 31232 24593 31260
rect 24544 31220 24550 31232
rect 24581 31229 24593 31232
rect 24627 31229 24639 31263
rect 24581 31223 24639 31229
rect 26142 31220 26148 31272
rect 26200 31260 26206 31272
rect 27448 31260 27476 31291
rect 27890 31288 27896 31300
rect 27948 31288 27954 31340
rect 28350 31328 28356 31340
rect 28311 31300 28356 31328
rect 28350 31288 28356 31300
rect 28408 31288 28414 31340
rect 26200 31232 27476 31260
rect 26200 31220 26206 31232
rect 20073 31195 20131 31201
rect 20073 31192 20085 31195
rect 18432 31164 20085 31192
rect 16853 31127 16911 31133
rect 16853 31124 16865 31127
rect 14384 31096 16865 31124
rect 16853 31093 16865 31096
rect 16899 31093 16911 31127
rect 16853 31087 16911 31093
rect 16942 31084 16948 31136
rect 17000 31124 17006 31136
rect 18432 31124 18460 31164
rect 20073 31161 20085 31164
rect 20119 31161 20131 31195
rect 20073 31155 20131 31161
rect 21910 31152 21916 31204
rect 21968 31192 21974 31204
rect 22005 31195 22063 31201
rect 22005 31192 22017 31195
rect 21968 31164 22017 31192
rect 21968 31152 21974 31164
rect 22005 31161 22017 31164
rect 22051 31161 22063 31195
rect 27709 31195 27767 31201
rect 27709 31192 27721 31195
rect 22005 31155 22063 31161
rect 23768 31164 24072 31192
rect 17000 31096 18460 31124
rect 18877 31127 18935 31133
rect 17000 31084 17006 31096
rect 18877 31093 18889 31127
rect 18923 31124 18935 31127
rect 19242 31124 19248 31136
rect 18923 31096 19248 31124
rect 18923 31093 18935 31096
rect 18877 31087 18935 31093
rect 19242 31084 19248 31096
rect 19300 31084 19306 31136
rect 19426 31124 19432 31136
rect 19387 31096 19432 31124
rect 19426 31084 19432 31096
rect 19484 31084 19490 31136
rect 19886 31084 19892 31136
rect 19944 31124 19950 31136
rect 20530 31124 20536 31136
rect 19944 31096 20536 31124
rect 19944 31084 19950 31096
rect 20530 31084 20536 31096
rect 20588 31084 20594 31136
rect 20714 31084 20720 31136
rect 20772 31124 20778 31136
rect 23768 31124 23796 31164
rect 20772 31096 23796 31124
rect 20772 31084 20778 31096
rect 23842 31084 23848 31136
rect 23900 31124 23906 31136
rect 24044 31124 24072 31164
rect 25792 31164 27721 31192
rect 25792 31124 25820 31164
rect 27709 31161 27721 31164
rect 27755 31161 27767 31195
rect 27709 31155 27767 31161
rect 25958 31124 25964 31136
rect 23900 31096 23945 31124
rect 24044 31096 25820 31124
rect 25919 31096 25964 31124
rect 23900 31084 23906 31096
rect 25958 31084 25964 31096
rect 26016 31084 26022 31136
rect 26418 31124 26424 31136
rect 26379 31096 26424 31124
rect 26418 31084 26424 31096
rect 26476 31084 26482 31136
rect 1104 31034 28888 31056
rect 1104 30982 4423 31034
rect 4475 30982 4487 31034
rect 4539 30982 4551 31034
rect 4603 30982 4615 31034
rect 4667 30982 4679 31034
rect 4731 30982 11369 31034
rect 11421 30982 11433 31034
rect 11485 30982 11497 31034
rect 11549 30982 11561 31034
rect 11613 30982 11625 31034
rect 11677 30982 18315 31034
rect 18367 30982 18379 31034
rect 18431 30982 18443 31034
rect 18495 30982 18507 31034
rect 18559 30982 18571 31034
rect 18623 30982 25261 31034
rect 25313 30982 25325 31034
rect 25377 30982 25389 31034
rect 25441 30982 25453 31034
rect 25505 30982 25517 31034
rect 25569 30982 28888 31034
rect 1104 30960 28888 30982
rect 6178 30920 6184 30932
rect 6139 30892 6184 30920
rect 6178 30880 6184 30892
rect 6236 30920 6242 30932
rect 7742 30920 7748 30932
rect 6236 30892 7748 30920
rect 6236 30880 6242 30892
rect 7742 30880 7748 30892
rect 7800 30880 7806 30932
rect 8478 30880 8484 30932
rect 8536 30920 8542 30932
rect 9309 30923 9367 30929
rect 9309 30920 9321 30923
rect 8536 30892 9321 30920
rect 8536 30880 8542 30892
rect 9309 30889 9321 30892
rect 9355 30889 9367 30923
rect 11238 30920 11244 30932
rect 9309 30883 9367 30889
rect 10060 30892 11244 30920
rect 7929 30855 7987 30861
rect 7929 30821 7941 30855
rect 7975 30852 7987 30855
rect 8662 30852 8668 30864
rect 7975 30824 8668 30852
rect 7975 30821 7987 30824
rect 7929 30815 7987 30821
rect 8662 30812 8668 30824
rect 8720 30812 8726 30864
rect 5169 30787 5227 30793
rect 5169 30753 5181 30787
rect 5215 30784 5227 30787
rect 7098 30784 7104 30796
rect 5215 30756 7104 30784
rect 5215 30753 5227 30756
rect 5169 30747 5227 30753
rect 7098 30744 7104 30756
rect 7156 30744 7162 30796
rect 10060 30784 10088 30892
rect 11238 30880 11244 30892
rect 11296 30920 11302 30932
rect 11609 30923 11667 30929
rect 11609 30920 11621 30923
rect 11296 30892 11621 30920
rect 11296 30880 11302 30892
rect 11609 30889 11621 30892
rect 11655 30889 11667 30923
rect 11790 30920 11796 30932
rect 11751 30892 11796 30920
rect 11609 30883 11667 30889
rect 11790 30880 11796 30892
rect 11848 30880 11854 30932
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 13262 30920 13268 30932
rect 12492 30892 13268 30920
rect 12492 30880 12498 30892
rect 13262 30880 13268 30892
rect 13320 30880 13326 30932
rect 16132 30892 18920 30920
rect 10137 30855 10195 30861
rect 10137 30821 10149 30855
rect 10183 30852 10195 30855
rect 16132 30852 16160 30892
rect 17494 30852 17500 30864
rect 10183 30824 16160 30852
rect 17455 30824 17500 30852
rect 10183 30821 10195 30824
rect 10137 30815 10195 30821
rect 17494 30812 17500 30824
rect 17552 30812 17558 30864
rect 18892 30852 18920 30892
rect 18966 30880 18972 30932
rect 19024 30920 19030 30932
rect 20346 30920 20352 30932
rect 19024 30892 20352 30920
rect 19024 30880 19030 30892
rect 20346 30880 20352 30892
rect 20404 30880 20410 30932
rect 20622 30920 20628 30932
rect 20583 30892 20628 30920
rect 20622 30880 20628 30892
rect 20680 30880 20686 30932
rect 21726 30880 21732 30932
rect 21784 30920 21790 30932
rect 25958 30920 25964 30932
rect 21784 30892 25964 30920
rect 21784 30880 21790 30892
rect 25958 30880 25964 30892
rect 26016 30880 26022 30932
rect 20254 30852 20260 30864
rect 18892 30824 20260 30852
rect 20254 30812 20260 30824
rect 20312 30812 20318 30864
rect 20364 30824 21128 30852
rect 11698 30784 11704 30796
rect 8220 30756 10088 30784
rect 1578 30716 1584 30728
rect 1539 30688 1584 30716
rect 1578 30676 1584 30688
rect 1636 30676 1642 30728
rect 4065 30719 4123 30725
rect 4065 30685 4077 30719
rect 4111 30716 4123 30719
rect 8220 30716 8248 30756
rect 11697 30744 11704 30784
rect 11756 30784 11762 30796
rect 11882 30784 11888 30796
rect 11756 30756 11888 30784
rect 11756 30744 11762 30756
rect 11882 30744 11888 30756
rect 11940 30744 11946 30796
rect 12434 30784 12440 30796
rect 12268 30756 12440 30784
rect 8386 30716 8392 30728
rect 4111 30688 8248 30716
rect 8347 30688 8392 30716
rect 4111 30685 4123 30688
rect 4065 30679 4123 30685
rect 8386 30676 8392 30688
rect 8444 30676 8450 30728
rect 9306 30676 9312 30728
rect 9364 30716 9370 30728
rect 9493 30719 9551 30725
rect 9493 30716 9505 30719
rect 9364 30688 9505 30716
rect 9364 30676 9370 30688
rect 9493 30685 9505 30688
rect 9539 30685 9551 30719
rect 9493 30679 9551 30685
rect 9953 30719 10011 30725
rect 9953 30685 9965 30719
rect 9999 30685 10011 30719
rect 11697 30691 11725 30744
rect 12268 30725 12296 30756
rect 12434 30744 12440 30756
rect 12492 30744 12498 30796
rect 12713 30787 12771 30793
rect 12713 30753 12725 30787
rect 12759 30784 12771 30787
rect 17310 30784 17316 30796
rect 12759 30756 16088 30784
rect 12759 30753 12771 30756
rect 12713 30747 12771 30753
rect 9953 30679 10011 30685
rect 11655 30685 11725 30691
rect 6825 30651 6883 30657
rect 6825 30617 6837 30651
rect 6871 30648 6883 30651
rect 8478 30648 8484 30660
rect 6871 30620 8484 30648
rect 6871 30617 6883 30620
rect 6825 30611 6883 30617
rect 8478 30608 8484 30620
rect 8536 30608 8542 30660
rect 9968 30648 9996 30679
rect 8588 30620 9996 30648
rect 3418 30580 3424 30592
rect 3379 30552 3424 30580
rect 3418 30540 3424 30552
rect 3476 30540 3482 30592
rect 4617 30583 4675 30589
rect 4617 30549 4629 30583
rect 4663 30580 4675 30583
rect 4798 30580 4804 30592
rect 4663 30552 4804 30580
rect 4663 30549 4675 30552
rect 4617 30543 4675 30549
rect 4798 30540 4804 30552
rect 4856 30540 4862 30592
rect 5718 30580 5724 30592
rect 5679 30552 5724 30580
rect 5718 30540 5724 30552
rect 5776 30540 5782 30592
rect 7374 30580 7380 30592
rect 7335 30552 7380 30580
rect 7374 30540 7380 30552
rect 7432 30540 7438 30592
rect 8588 30589 8616 30620
rect 10042 30608 10048 30660
rect 10100 30648 10106 30660
rect 10781 30651 10839 30657
rect 10781 30648 10793 30651
rect 10100 30620 10793 30648
rect 10100 30608 10106 30620
rect 10781 30617 10793 30620
rect 10827 30648 10839 30651
rect 11146 30648 11152 30660
rect 10827 30620 11152 30648
rect 10827 30617 10839 30620
rect 10781 30611 10839 30617
rect 11146 30608 11152 30620
rect 11204 30608 11210 30660
rect 11425 30651 11483 30657
rect 11425 30617 11437 30651
rect 11471 30617 11483 30651
rect 11655 30651 11667 30685
rect 11701 30654 11725 30685
rect 12253 30719 12311 30725
rect 12253 30685 12265 30719
rect 12299 30685 12311 30719
rect 12253 30679 12311 30685
rect 12342 30676 12348 30728
rect 12400 30676 12406 30728
rect 13170 30716 13176 30728
rect 13131 30688 13176 30716
rect 13170 30676 13176 30688
rect 13228 30676 13234 30728
rect 13262 30676 13268 30728
rect 13320 30716 13326 30728
rect 13446 30716 13452 30728
rect 13320 30688 13365 30716
rect 13407 30688 13452 30716
rect 13320 30676 13326 30688
rect 13446 30676 13452 30688
rect 13504 30676 13510 30728
rect 13541 30719 13599 30725
rect 13541 30685 13553 30719
rect 13587 30685 13599 30719
rect 13541 30679 13599 30685
rect 13725 30719 13783 30725
rect 13725 30685 13737 30719
rect 13771 30716 13783 30719
rect 13998 30716 14004 30728
rect 13771 30688 14004 30716
rect 13771 30685 13783 30688
rect 13725 30679 13783 30685
rect 11701 30651 11713 30654
rect 11655 30645 11713 30651
rect 12066 30648 12072 30660
rect 11425 30611 11483 30617
rect 11808 30620 12072 30648
rect 8573 30583 8631 30589
rect 8573 30549 8585 30583
rect 8619 30549 8631 30583
rect 8573 30543 8631 30549
rect 8662 30540 8668 30592
rect 8720 30580 8726 30592
rect 10873 30583 10931 30589
rect 10873 30580 10885 30583
rect 8720 30552 10885 30580
rect 8720 30540 8726 30552
rect 10873 30549 10885 30552
rect 10919 30580 10931 30583
rect 11054 30580 11060 30592
rect 10919 30552 11060 30580
rect 10919 30549 10931 30552
rect 10873 30543 10931 30549
rect 11054 30540 11060 30552
rect 11112 30540 11118 30592
rect 11440 30580 11468 30611
rect 11808 30580 11836 30620
rect 12066 30608 12072 30620
rect 12124 30608 12130 30660
rect 12360 30648 12388 30676
rect 13556 30648 13584 30679
rect 13998 30676 14004 30688
rect 14056 30676 14062 30728
rect 14550 30676 14556 30728
rect 14608 30716 14614 30728
rect 14829 30719 14887 30725
rect 14829 30716 14841 30719
rect 14608 30688 14841 30716
rect 14608 30676 14614 30688
rect 14829 30685 14841 30688
rect 14875 30685 14887 30719
rect 14829 30679 14887 30685
rect 14921 30719 14979 30725
rect 14921 30685 14933 30719
rect 14967 30685 14979 30719
rect 15102 30716 15108 30728
rect 15063 30688 15108 30716
rect 14921 30679 14979 30685
rect 12360 30620 13584 30648
rect 14936 30648 14964 30679
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 15197 30719 15255 30725
rect 15197 30685 15209 30719
rect 15243 30716 15255 30719
rect 15286 30716 15292 30728
rect 15243 30688 15292 30716
rect 15243 30685 15255 30688
rect 15197 30679 15255 30685
rect 15286 30676 15292 30688
rect 15344 30676 15350 30728
rect 16060 30716 16088 30756
rect 16960 30756 17316 30784
rect 16960 30716 16988 30756
rect 17310 30744 17316 30756
rect 17368 30744 17374 30796
rect 18874 30784 18880 30796
rect 18835 30756 18880 30784
rect 18874 30744 18880 30756
rect 18932 30744 18938 30796
rect 19886 30784 19892 30796
rect 19306 30756 19892 30784
rect 16060 30688 16988 30716
rect 17037 30719 17095 30725
rect 17037 30685 17049 30719
rect 17083 30716 17095 30719
rect 17678 30716 17684 30728
rect 17083 30688 17684 30716
rect 17083 30685 17095 30688
rect 17037 30679 17095 30685
rect 17678 30676 17684 30688
rect 17736 30676 17742 30728
rect 18230 30716 18236 30728
rect 17880 30688 18236 30716
rect 16298 30648 16304 30660
rect 14936 30620 16304 30648
rect 16298 30608 16304 30620
rect 16356 30608 16362 30660
rect 16792 30651 16850 30657
rect 16792 30617 16804 30651
rect 16838 30648 16850 30651
rect 17880 30648 17908 30688
rect 18230 30676 18236 30688
rect 18288 30676 18294 30728
rect 19058 30676 19064 30728
rect 19116 30716 19122 30728
rect 19306 30716 19334 30756
rect 19886 30744 19892 30756
rect 19944 30744 19950 30796
rect 20162 30744 20168 30796
rect 20220 30784 20226 30796
rect 20364 30784 20392 30824
rect 20530 30784 20536 30796
rect 20220 30756 20392 30784
rect 20456 30756 20536 30784
rect 20220 30744 20226 30756
rect 19116 30688 19334 30716
rect 19981 30719 20039 30725
rect 19116 30676 19122 30688
rect 19981 30685 19993 30719
rect 20027 30685 20039 30719
rect 20346 30716 20352 30728
rect 20307 30688 20352 30716
rect 19981 30679 20039 30685
rect 16838 30620 17908 30648
rect 16838 30617 16850 30620
rect 16792 30611 16850 30617
rect 17954 30608 17960 30660
rect 18012 30648 18018 30660
rect 18632 30651 18690 30657
rect 18632 30648 18644 30651
rect 18012 30620 18644 30648
rect 18012 30608 18018 30620
rect 18632 30617 18644 30620
rect 18678 30648 18690 30651
rect 19610 30648 19616 30660
rect 18678 30620 19616 30648
rect 18678 30617 18690 30620
rect 18632 30611 18690 30617
rect 19610 30608 19616 30620
rect 19668 30608 19674 30660
rect 11440 30552 11836 30580
rect 11974 30540 11980 30592
rect 12032 30580 12038 30592
rect 12345 30583 12403 30589
rect 12345 30580 12357 30583
rect 12032 30552 12357 30580
rect 12032 30540 12038 30552
rect 12345 30549 12357 30552
rect 12391 30549 12403 30583
rect 12345 30543 12403 30549
rect 12437 30583 12495 30589
rect 12437 30549 12449 30583
rect 12483 30580 12495 30583
rect 13630 30580 13636 30592
rect 12483 30552 13636 30580
rect 12483 30549 12495 30552
rect 12437 30543 12495 30549
rect 13630 30540 13636 30552
rect 13688 30540 13694 30592
rect 14642 30580 14648 30592
rect 14603 30552 14648 30580
rect 14642 30540 14648 30552
rect 14700 30540 14706 30592
rect 15654 30580 15660 30592
rect 15615 30552 15660 30580
rect 15654 30540 15660 30552
rect 15712 30540 15718 30592
rect 17862 30540 17868 30592
rect 17920 30580 17926 30592
rect 19429 30583 19487 30589
rect 19429 30580 19441 30583
rect 17920 30552 19441 30580
rect 17920 30540 17926 30552
rect 19429 30549 19441 30552
rect 19475 30549 19487 30583
rect 19996 30580 20024 30679
rect 20346 30676 20352 30688
rect 20404 30676 20410 30728
rect 20456 30725 20484 30756
rect 20530 30744 20536 30756
rect 20588 30744 20594 30796
rect 21100 30793 21128 30824
rect 21085 30787 21143 30793
rect 21085 30753 21097 30787
rect 21131 30753 21143 30787
rect 21085 30747 21143 30753
rect 20441 30719 20499 30725
rect 20441 30685 20453 30719
rect 20487 30685 20499 30719
rect 21100 30716 21128 30747
rect 22094 30744 22100 30796
rect 22152 30784 22158 30796
rect 22152 30756 23980 30784
rect 22152 30744 22158 30756
rect 23952 30728 23980 30756
rect 25884 30756 26188 30784
rect 21174 30716 21180 30728
rect 21100 30688 21180 30716
rect 20441 30679 20499 30685
rect 21174 30676 21180 30688
rect 21232 30676 21238 30728
rect 21910 30716 21916 30728
rect 21284 30688 21916 30716
rect 20070 30608 20076 30660
rect 20128 30657 20134 30660
rect 20128 30651 20177 30657
rect 20128 30617 20131 30651
rect 20165 30617 20177 30651
rect 20128 30611 20177 30617
rect 20128 30608 20134 30611
rect 20254 30608 20260 30660
rect 20312 30648 20318 30660
rect 20312 30620 20357 30648
rect 20312 30608 20318 30620
rect 20530 30608 20536 30660
rect 20588 30648 20594 30660
rect 21284 30648 21312 30688
rect 21910 30676 21916 30688
rect 21968 30676 21974 30728
rect 22646 30676 22652 30728
rect 22704 30716 22710 30728
rect 23474 30716 23480 30728
rect 22704 30688 23480 30716
rect 22704 30676 22710 30688
rect 23474 30676 23480 30688
rect 23532 30676 23538 30728
rect 23750 30716 23756 30728
rect 23711 30688 23756 30716
rect 23750 30676 23756 30688
rect 23808 30676 23814 30728
rect 23934 30676 23940 30728
rect 23992 30716 23998 30728
rect 25884 30716 25912 30756
rect 23992 30688 25912 30716
rect 23992 30676 23998 30688
rect 25958 30676 25964 30728
rect 26016 30716 26022 30728
rect 26160 30716 26188 30756
rect 27801 30719 27859 30725
rect 27801 30716 27813 30719
rect 26016 30688 26061 30716
rect 26160 30688 27813 30716
rect 26016 30676 26022 30688
rect 27801 30685 27813 30688
rect 27847 30716 27859 30719
rect 28074 30716 28080 30728
rect 27847 30688 28080 30716
rect 27847 30685 27859 30688
rect 27801 30679 27859 30685
rect 28074 30676 28080 30688
rect 28132 30676 28138 30728
rect 20588 30620 21312 30648
rect 21352 30651 21410 30657
rect 20588 30608 20594 30620
rect 21352 30617 21364 30651
rect 21398 30648 21410 30651
rect 21634 30648 21640 30660
rect 21398 30620 21640 30648
rect 21398 30617 21410 30620
rect 21352 30611 21410 30617
rect 21634 30608 21640 30620
rect 21692 30608 21698 30660
rect 21726 30608 21732 30660
rect 21784 30648 21790 30660
rect 25694 30651 25752 30657
rect 25694 30648 25706 30651
rect 21784 30620 25706 30648
rect 21784 30608 21790 30620
rect 25694 30617 25706 30620
rect 25740 30617 25752 30651
rect 27534 30651 27592 30657
rect 27534 30648 27546 30651
rect 25694 30611 25752 30617
rect 25792 30620 27546 30648
rect 21542 30580 21548 30592
rect 19996 30552 21548 30580
rect 19429 30543 19487 30549
rect 21542 30540 21548 30552
rect 21600 30540 21606 30592
rect 22465 30583 22523 30589
rect 22465 30549 22477 30583
rect 22511 30580 22523 30583
rect 22646 30580 22652 30592
rect 22511 30552 22652 30580
rect 22511 30549 22523 30552
rect 22465 30543 22523 30549
rect 22646 30540 22652 30552
rect 22704 30540 22710 30592
rect 23474 30540 23480 30592
rect 23532 30580 23538 30592
rect 24302 30580 24308 30592
rect 23532 30552 24308 30580
rect 23532 30540 23538 30552
rect 24302 30540 24308 30552
rect 24360 30540 24366 30592
rect 24578 30580 24584 30592
rect 24539 30552 24584 30580
rect 24578 30540 24584 30552
rect 24636 30540 24642 30592
rect 25038 30540 25044 30592
rect 25096 30580 25102 30592
rect 25792 30580 25820 30620
rect 27534 30617 27546 30620
rect 27580 30617 27592 30651
rect 27534 30611 27592 30617
rect 26418 30580 26424 30592
rect 25096 30552 25820 30580
rect 26379 30552 26424 30580
rect 25096 30540 25102 30552
rect 26418 30540 26424 30552
rect 26476 30540 26482 30592
rect 28258 30580 28264 30592
rect 28219 30552 28264 30580
rect 28258 30540 28264 30552
rect 28316 30540 28322 30592
rect 1104 30490 29048 30512
rect 1104 30438 7896 30490
rect 7948 30438 7960 30490
rect 8012 30438 8024 30490
rect 8076 30438 8088 30490
rect 8140 30438 8152 30490
rect 8204 30438 14842 30490
rect 14894 30438 14906 30490
rect 14958 30438 14970 30490
rect 15022 30438 15034 30490
rect 15086 30438 15098 30490
rect 15150 30438 21788 30490
rect 21840 30438 21852 30490
rect 21904 30438 21916 30490
rect 21968 30438 21980 30490
rect 22032 30438 22044 30490
rect 22096 30438 28734 30490
rect 28786 30438 28798 30490
rect 28850 30438 28862 30490
rect 28914 30438 28926 30490
rect 28978 30438 28990 30490
rect 29042 30438 29048 30490
rect 1104 30416 29048 30438
rect 3418 30336 3424 30388
rect 3476 30376 3482 30388
rect 6546 30376 6552 30388
rect 3476 30348 6552 30376
rect 3476 30336 3482 30348
rect 6546 30336 6552 30348
rect 6604 30336 6610 30388
rect 9950 30376 9956 30388
rect 7116 30348 9956 30376
rect 7116 30320 7144 30348
rect 9950 30336 9956 30348
rect 10008 30336 10014 30388
rect 10134 30336 10140 30388
rect 10192 30376 10198 30388
rect 16390 30376 16396 30388
rect 10192 30348 16396 30376
rect 10192 30336 10198 30348
rect 16390 30336 16396 30348
rect 16448 30336 16454 30388
rect 17034 30336 17040 30388
rect 17092 30376 17098 30388
rect 17129 30379 17187 30385
rect 17129 30376 17141 30379
rect 17092 30348 17141 30376
rect 17092 30336 17098 30348
rect 17129 30345 17141 30348
rect 17175 30345 17187 30379
rect 17129 30339 17187 30345
rect 17310 30336 17316 30388
rect 17368 30376 17374 30388
rect 24578 30376 24584 30388
rect 17368 30348 24584 30376
rect 17368 30336 17374 30348
rect 24578 30336 24584 30348
rect 24636 30336 24642 30388
rect 25038 30376 25044 30388
rect 24688 30348 25044 30376
rect 5445 30311 5503 30317
rect 5445 30277 5457 30311
rect 5491 30308 5503 30311
rect 5718 30308 5724 30320
rect 5491 30280 5724 30308
rect 5491 30277 5503 30280
rect 5445 30271 5503 30277
rect 5718 30268 5724 30280
rect 5776 30268 5782 30320
rect 7098 30308 7104 30320
rect 7059 30280 7104 30308
rect 7098 30268 7104 30280
rect 7156 30268 7162 30320
rect 7650 30268 7656 30320
rect 7708 30308 7714 30320
rect 8205 30311 8263 30317
rect 8205 30308 8217 30311
rect 7708 30280 8217 30308
rect 7708 30268 7714 30280
rect 8205 30277 8217 30280
rect 8251 30308 8263 30311
rect 8938 30308 8944 30320
rect 8251 30280 8944 30308
rect 8251 30277 8263 30280
rect 8205 30271 8263 30277
rect 8938 30268 8944 30280
rect 8996 30268 9002 30320
rect 10594 30308 10600 30320
rect 9232 30280 10600 30308
rect 4341 30243 4399 30249
rect 4341 30209 4353 30243
rect 4387 30240 4399 30243
rect 9232 30240 9260 30280
rect 10594 30268 10600 30280
rect 10652 30268 10658 30320
rect 10781 30311 10839 30317
rect 10781 30277 10793 30311
rect 10827 30277 10839 30311
rect 10781 30271 10839 30277
rect 9398 30240 9404 30252
rect 4387 30212 9260 30240
rect 9359 30212 9404 30240
rect 4387 30209 4399 30212
rect 4341 30203 4399 30209
rect 9398 30200 9404 30212
rect 9456 30200 9462 30252
rect 10229 30243 10287 30249
rect 10229 30209 10241 30243
rect 10275 30240 10287 30243
rect 10796 30240 10824 30271
rect 10870 30268 10876 30320
rect 10928 30308 10934 30320
rect 10981 30311 11039 30317
rect 10981 30308 10993 30311
rect 10928 30280 10993 30308
rect 10928 30268 10934 30280
rect 10981 30277 10993 30280
rect 11027 30277 11039 30311
rect 10981 30271 11039 30277
rect 11146 30268 11152 30320
rect 11204 30308 11210 30320
rect 12894 30308 12900 30320
rect 11204 30280 12900 30308
rect 11204 30268 11210 30280
rect 11698 30240 11704 30252
rect 10275 30212 10732 30240
rect 10796 30212 11704 30240
rect 10275 30209 10287 30212
rect 10229 30203 10287 30209
rect 5534 30132 5540 30184
rect 5592 30172 5598 30184
rect 5997 30175 6055 30181
rect 5997 30172 6009 30175
rect 5592 30144 6009 30172
rect 5592 30132 5598 30144
rect 5997 30141 6009 30144
rect 6043 30172 6055 30175
rect 8570 30172 8576 30184
rect 6043 30144 8576 30172
rect 6043 30141 6055 30144
rect 5997 30135 6055 30141
rect 8570 30132 8576 30144
rect 8628 30132 8634 30184
rect 8941 30175 8999 30181
rect 8941 30141 8953 30175
rect 8987 30172 8999 30175
rect 10502 30172 10508 30184
rect 8987 30144 10508 30172
rect 8987 30141 8999 30144
rect 8941 30135 8999 30141
rect 10502 30132 10508 30144
rect 10560 30132 10566 30184
rect 10704 30172 10732 30212
rect 11698 30200 11704 30212
rect 11756 30200 11762 30252
rect 12250 30240 12256 30252
rect 12211 30212 12256 30240
rect 12250 30200 12256 30212
rect 12308 30200 12314 30252
rect 12544 30249 12572 30280
rect 12894 30268 12900 30280
rect 12952 30268 12958 30320
rect 14366 30308 14372 30320
rect 13004 30280 14372 30308
rect 12345 30243 12403 30249
rect 12345 30209 12357 30243
rect 12391 30209 12403 30243
rect 12345 30203 12403 30209
rect 12529 30243 12587 30249
rect 12529 30209 12541 30243
rect 12575 30209 12587 30243
rect 12529 30203 12587 30209
rect 10778 30172 10784 30184
rect 10704 30144 10784 30172
rect 10778 30132 10784 30144
rect 10836 30132 10842 30184
rect 12268 30172 12296 30200
rect 10888 30144 12296 30172
rect 12360 30172 12388 30203
rect 12618 30200 12624 30252
rect 12676 30240 12682 30252
rect 12676 30212 12721 30240
rect 12676 30200 12682 30212
rect 13004 30172 13032 30280
rect 14366 30268 14372 30280
rect 14424 30268 14430 30320
rect 14642 30268 14648 30320
rect 14700 30308 14706 30320
rect 17615 30311 17673 30317
rect 17615 30308 17627 30311
rect 14700 30280 17627 30308
rect 14700 30268 14706 30280
rect 17615 30277 17627 30280
rect 17661 30277 17673 30311
rect 17615 30271 17673 30277
rect 19368 30311 19426 30317
rect 19368 30277 19380 30311
rect 19414 30308 19426 30311
rect 20622 30308 20628 30320
rect 19414 30280 20628 30308
rect 19414 30277 19426 30280
rect 19368 30271 19426 30277
rect 20622 30268 20628 30280
rect 20680 30268 20686 30320
rect 23842 30308 23848 30320
rect 22066 30280 23848 30308
rect 13354 30249 13360 30252
rect 13348 30240 13360 30249
rect 13315 30212 13360 30240
rect 13348 30203 13360 30212
rect 13354 30200 13360 30203
rect 13412 30200 13418 30252
rect 15746 30240 15752 30252
rect 14384 30212 15752 30240
rect 12360 30144 13032 30172
rect 13081 30175 13139 30181
rect 7745 30107 7803 30113
rect 7745 30073 7757 30107
rect 7791 30104 7803 30107
rect 9766 30104 9772 30116
rect 7791 30076 9772 30104
rect 7791 30073 7803 30076
rect 7745 30067 7803 30073
rect 9766 30064 9772 30076
rect 9824 30064 9830 30116
rect 9950 30064 9956 30116
rect 10008 30104 10014 30116
rect 10318 30104 10324 30116
rect 10008 30076 10324 30104
rect 10008 30064 10014 30076
rect 10318 30064 10324 30076
rect 10376 30064 10382 30116
rect 10888 30104 10916 30144
rect 13081 30141 13093 30175
rect 13127 30141 13139 30175
rect 13081 30135 13139 30141
rect 11146 30104 11152 30116
rect 10520 30076 10916 30104
rect 11107 30076 11152 30104
rect 4893 30039 4951 30045
rect 4893 30005 4905 30039
rect 4939 30036 4951 30039
rect 6822 30036 6828 30048
rect 4939 30008 6828 30036
rect 4939 30005 4951 30008
rect 4893 29999 4951 30005
rect 6822 29996 6828 30008
rect 6880 29996 6886 30048
rect 8294 29996 8300 30048
rect 8352 30036 8358 30048
rect 9582 30036 9588 30048
rect 8352 30008 9588 30036
rect 8352 29996 8358 30008
rect 9582 29996 9588 30008
rect 9640 29996 9646 30048
rect 10134 30036 10140 30048
rect 10047 30008 10140 30036
rect 10134 29996 10140 30008
rect 10192 30036 10198 30048
rect 10520 30036 10548 30076
rect 11146 30064 11152 30076
rect 11204 30064 11210 30116
rect 12802 30064 12808 30116
rect 12860 30104 12866 30116
rect 13096 30104 13124 30135
rect 12860 30076 13124 30104
rect 12860 30064 12866 30076
rect 10192 30008 10548 30036
rect 10192 29996 10198 30008
rect 10594 29996 10600 30048
rect 10652 30036 10658 30048
rect 10962 30036 10968 30048
rect 10652 30008 10968 30036
rect 10652 29996 10658 30008
rect 10962 29996 10968 30008
rect 11020 29996 11026 30048
rect 12066 30036 12072 30048
rect 12027 30008 12072 30036
rect 12066 29996 12072 30008
rect 12124 29996 12130 30048
rect 12158 29996 12164 30048
rect 12216 30036 12222 30048
rect 14384 30036 14412 30212
rect 15746 30200 15752 30212
rect 15804 30200 15810 30252
rect 16022 30240 16028 30252
rect 16080 30249 16086 30252
rect 16080 30243 16103 30249
rect 15955 30212 16028 30240
rect 16022 30200 16028 30212
rect 16091 30240 16103 30243
rect 16942 30240 16948 30252
rect 16091 30212 16948 30240
rect 16091 30209 16103 30212
rect 16080 30203 16103 30209
rect 16080 30200 16086 30203
rect 16942 30200 16948 30212
rect 17000 30200 17006 30252
rect 17313 30243 17371 30249
rect 17313 30240 17325 30243
rect 17052 30212 17325 30240
rect 16301 30175 16359 30181
rect 16301 30141 16313 30175
rect 16347 30141 16359 30175
rect 16301 30135 16359 30141
rect 14458 30064 14464 30116
rect 14516 30104 14522 30116
rect 16316 30104 16344 30135
rect 16850 30132 16856 30184
rect 16908 30172 16914 30184
rect 17052 30172 17080 30212
rect 17313 30209 17325 30212
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 17405 30243 17463 30249
rect 17405 30209 17417 30243
rect 17451 30209 17463 30243
rect 17405 30203 17463 30209
rect 16908 30144 17080 30172
rect 16908 30132 16914 30144
rect 17218 30132 17224 30184
rect 17276 30172 17282 30184
rect 17420 30172 17448 30203
rect 17494 30200 17500 30252
rect 17552 30240 17558 30252
rect 17552 30212 17597 30240
rect 17630 30212 19656 30240
rect 17552 30200 17558 30212
rect 17276 30144 17448 30172
rect 17276 30132 17282 30144
rect 16482 30104 16488 30116
rect 14516 30076 15056 30104
rect 16316 30076 16488 30104
rect 14516 30064 14522 30076
rect 12216 30008 14412 30036
rect 12216 29996 12222 30008
rect 14826 29996 14832 30048
rect 14884 30036 14890 30048
rect 14921 30039 14979 30045
rect 14921 30036 14933 30039
rect 14884 30008 14933 30036
rect 14884 29996 14890 30008
rect 14921 30005 14933 30008
rect 14967 30005 14979 30039
rect 15028 30036 15056 30076
rect 16482 30064 16488 30076
rect 16540 30104 16546 30116
rect 17630 30104 17658 30212
rect 17773 30175 17831 30181
rect 17773 30141 17785 30175
rect 17819 30172 17831 30175
rect 18598 30172 18604 30184
rect 17819 30144 18604 30172
rect 17819 30141 17831 30144
rect 17773 30135 17831 30141
rect 18598 30132 18604 30144
rect 18656 30132 18662 30184
rect 19628 30181 19656 30212
rect 19702 30200 19708 30252
rect 19760 30240 19766 30252
rect 20346 30249 20352 30252
rect 20073 30243 20131 30249
rect 20073 30240 20085 30243
rect 19760 30212 20085 30240
rect 19760 30200 19766 30212
rect 20073 30209 20085 30212
rect 20119 30209 20131 30243
rect 20340 30240 20352 30249
rect 20307 30212 20352 30240
rect 20073 30203 20131 30209
rect 20340 30203 20352 30212
rect 20346 30200 20352 30203
rect 20404 30200 20410 30252
rect 22066 30240 22094 30280
rect 23842 30268 23848 30280
rect 23900 30268 23906 30320
rect 24210 30268 24216 30320
rect 24268 30308 24274 30320
rect 24688 30308 24716 30348
rect 25038 30336 25044 30348
rect 25096 30336 25102 30388
rect 25222 30376 25228 30388
rect 25183 30348 25228 30376
rect 25222 30336 25228 30348
rect 25280 30336 25286 30388
rect 27154 30376 27160 30388
rect 27115 30348 27160 30376
rect 27154 30336 27160 30348
rect 27212 30336 27218 30388
rect 27338 30336 27344 30388
rect 27396 30376 27402 30388
rect 27396 30348 27476 30376
rect 27396 30336 27402 30348
rect 27448 30317 27476 30348
rect 27522 30336 27528 30388
rect 27580 30336 27586 30388
rect 24268 30280 24716 30308
rect 27433 30311 27491 30317
rect 24268 30268 24274 30280
rect 27433 30277 27445 30311
rect 27479 30308 27491 30311
rect 27549 30308 27577 30336
rect 27643 30311 27701 30317
rect 27643 30308 27655 30311
rect 27479 30280 27513 30308
rect 27549 30280 27655 30308
rect 27479 30277 27491 30280
rect 27433 30271 27491 30277
rect 27643 30277 27655 30280
rect 27689 30277 27701 30311
rect 27643 30271 27701 30277
rect 22278 30249 22284 30252
rect 21100 30212 22094 30240
rect 19613 30175 19671 30181
rect 19613 30141 19625 30175
rect 19659 30172 19671 30175
rect 19794 30172 19800 30184
rect 19659 30144 19800 30172
rect 19659 30141 19671 30144
rect 19613 30135 19671 30141
rect 19794 30132 19800 30144
rect 19852 30132 19858 30184
rect 16540 30076 17658 30104
rect 16540 30064 16546 30076
rect 15654 30036 15660 30048
rect 15028 30008 15660 30036
rect 14921 29999 14979 30005
rect 15654 29996 15660 30008
rect 15712 29996 15718 30048
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 18046 30036 18052 30048
rect 15988 30008 18052 30036
rect 15988 29996 15994 30008
rect 18046 29996 18052 30008
rect 18104 29996 18110 30048
rect 18138 29996 18144 30048
rect 18196 30036 18202 30048
rect 18233 30039 18291 30045
rect 18233 30036 18245 30039
rect 18196 30008 18245 30036
rect 18196 29996 18202 30008
rect 18233 30005 18245 30008
rect 18279 30005 18291 30039
rect 18233 29999 18291 30005
rect 18322 29996 18328 30048
rect 18380 30036 18386 30048
rect 21100 30036 21128 30212
rect 22272 30203 22284 30249
rect 22336 30240 22342 30252
rect 24101 30243 24159 30249
rect 24101 30240 24113 30243
rect 22336 30212 22372 30240
rect 23032 30212 24113 30240
rect 22278 30200 22284 30203
rect 22336 30200 22342 30212
rect 21174 30132 21180 30184
rect 21232 30172 21238 30184
rect 22005 30175 22063 30181
rect 22005 30172 22017 30175
rect 21232 30144 22017 30172
rect 21232 30132 21238 30144
rect 22005 30141 22017 30144
rect 22051 30141 22063 30175
rect 22005 30135 22063 30141
rect 21266 30064 21272 30116
rect 21324 30104 21330 30116
rect 21324 30076 22048 30104
rect 21324 30064 21330 30076
rect 18380 30008 21128 30036
rect 18380 29996 18386 30008
rect 21174 29996 21180 30048
rect 21232 30036 21238 30048
rect 21453 30039 21511 30045
rect 21453 30036 21465 30039
rect 21232 30008 21465 30036
rect 21232 29996 21238 30008
rect 21453 30005 21465 30008
rect 21499 30005 21511 30039
rect 22020 30036 22048 30076
rect 23032 30036 23060 30212
rect 24101 30209 24113 30212
rect 24147 30209 24159 30243
rect 24101 30203 24159 30209
rect 26237 30243 26295 30249
rect 26237 30209 26249 30243
rect 26283 30240 26295 30243
rect 26602 30240 26608 30252
rect 26283 30212 26608 30240
rect 26283 30209 26295 30212
rect 26237 30203 26295 30209
rect 26602 30200 26608 30212
rect 26660 30200 26666 30252
rect 26970 30200 26976 30252
rect 27028 30240 27034 30252
rect 27341 30243 27399 30249
rect 27341 30240 27353 30243
rect 27028 30212 27353 30240
rect 27028 30200 27034 30212
rect 27341 30209 27353 30212
rect 27387 30209 27399 30243
rect 27522 30240 27528 30252
rect 27483 30212 27528 30240
rect 27341 30203 27399 30209
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 23842 30172 23848 30184
rect 23803 30144 23848 30172
rect 23842 30132 23848 30144
rect 23900 30132 23906 30184
rect 26513 30175 26571 30181
rect 26513 30141 26525 30175
rect 26559 30172 26571 30175
rect 26694 30172 26700 30184
rect 26559 30144 26700 30172
rect 26559 30141 26571 30144
rect 26513 30135 26571 30141
rect 26694 30132 26700 30144
rect 26752 30132 26758 30184
rect 27801 30175 27859 30181
rect 27801 30141 27813 30175
rect 27847 30141 27859 30175
rect 27801 30135 27859 30141
rect 25682 30064 25688 30116
rect 25740 30104 25746 30116
rect 27816 30104 27844 30135
rect 25740 30076 27844 30104
rect 25740 30064 25746 30076
rect 23382 30036 23388 30048
rect 22020 30008 23060 30036
rect 23343 30008 23388 30036
rect 21453 29999 21511 30005
rect 23382 29996 23388 30008
rect 23440 29996 23446 30048
rect 25038 29996 25044 30048
rect 25096 30036 25102 30048
rect 28261 30039 28319 30045
rect 28261 30036 28273 30039
rect 25096 30008 28273 30036
rect 25096 29996 25102 30008
rect 28261 30005 28273 30008
rect 28307 30005 28319 30039
rect 28261 29999 28319 30005
rect 1104 29946 28888 29968
rect 1104 29894 4423 29946
rect 4475 29894 4487 29946
rect 4539 29894 4551 29946
rect 4603 29894 4615 29946
rect 4667 29894 4679 29946
rect 4731 29894 11369 29946
rect 11421 29894 11433 29946
rect 11485 29894 11497 29946
rect 11549 29894 11561 29946
rect 11613 29894 11625 29946
rect 11677 29894 18315 29946
rect 18367 29894 18379 29946
rect 18431 29894 18443 29946
rect 18495 29894 18507 29946
rect 18559 29894 18571 29946
rect 18623 29894 25261 29946
rect 25313 29894 25325 29946
rect 25377 29894 25389 29946
rect 25441 29894 25453 29946
rect 25505 29894 25517 29946
rect 25569 29894 28888 29946
rect 1104 29872 28888 29894
rect 5534 29792 5540 29844
rect 5592 29832 5598 29844
rect 5721 29835 5779 29841
rect 5721 29832 5733 29835
rect 5592 29804 5733 29832
rect 5592 29792 5598 29804
rect 5721 29801 5733 29804
rect 5767 29801 5779 29835
rect 5721 29795 5779 29801
rect 5810 29792 5816 29844
rect 5868 29832 5874 29844
rect 7929 29835 7987 29841
rect 7929 29832 7941 29835
rect 5868 29804 7941 29832
rect 5868 29792 5874 29804
rect 7929 29801 7941 29804
rect 7975 29832 7987 29835
rect 8294 29832 8300 29844
rect 7975 29804 8300 29832
rect 7975 29801 7987 29804
rect 7929 29795 7987 29801
rect 8294 29792 8300 29804
rect 8352 29792 8358 29844
rect 8478 29832 8484 29844
rect 8439 29804 8484 29832
rect 8478 29792 8484 29804
rect 8536 29832 8542 29844
rect 9628 29832 9634 29844
rect 8536 29804 9634 29832
rect 8536 29792 8542 29804
rect 9628 29792 9634 29804
rect 9686 29792 9692 29844
rect 9769 29835 9827 29841
rect 9769 29801 9781 29835
rect 9815 29832 9827 29835
rect 12526 29832 12532 29844
rect 9815 29804 12532 29832
rect 9815 29801 9827 29804
rect 9769 29795 9827 29801
rect 9876 29764 9904 29804
rect 12526 29792 12532 29804
rect 12584 29792 12590 29844
rect 12618 29792 12624 29844
rect 12676 29832 12682 29844
rect 14274 29832 14280 29844
rect 12676 29804 14280 29832
rect 12676 29792 12682 29804
rect 14274 29792 14280 29804
rect 14332 29792 14338 29844
rect 14384 29804 14872 29832
rect 9692 29736 9904 29764
rect 9953 29767 10011 29773
rect 4709 29699 4767 29705
rect 4709 29665 4721 29699
rect 4755 29696 4767 29699
rect 4798 29696 4804 29708
rect 4755 29668 4804 29696
rect 4755 29665 4767 29668
rect 4709 29659 4767 29665
rect 4798 29656 4804 29668
rect 4856 29696 4862 29708
rect 9692 29696 9720 29736
rect 9953 29733 9965 29767
rect 9999 29733 10011 29767
rect 9953 29727 10011 29733
rect 4856 29668 9720 29696
rect 9968 29696 9996 29727
rect 11054 29724 11060 29776
rect 11112 29764 11118 29776
rect 11606 29764 11612 29776
rect 11112 29736 11612 29764
rect 11112 29724 11118 29736
rect 11606 29724 11612 29736
rect 11664 29764 11670 29776
rect 11664 29736 11744 29764
rect 11664 29724 11670 29736
rect 9968 29668 10272 29696
rect 4856 29656 4862 29668
rect 1578 29628 1584 29640
rect 1539 29600 1584 29628
rect 1578 29588 1584 29600
rect 1636 29588 1642 29640
rect 5718 29588 5724 29640
rect 5776 29628 5782 29640
rect 7469 29631 7527 29637
rect 7469 29628 7481 29631
rect 5776 29600 7481 29628
rect 5776 29588 5782 29600
rect 7469 29597 7481 29600
rect 7515 29628 7527 29631
rect 10134 29628 10140 29640
rect 7515 29600 10140 29628
rect 7515 29597 7527 29600
rect 7469 29591 7527 29597
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 6273 29563 6331 29569
rect 6273 29529 6285 29563
rect 6319 29560 6331 29563
rect 9582 29560 9588 29572
rect 6319 29532 9444 29560
rect 9543 29532 9588 29560
rect 6319 29529 6331 29532
rect 6273 29523 6331 29529
rect 5258 29492 5264 29504
rect 5219 29464 5264 29492
rect 5258 29452 5264 29464
rect 5316 29452 5322 29504
rect 6914 29492 6920 29504
rect 6875 29464 6920 29492
rect 6914 29452 6920 29464
rect 6972 29452 6978 29504
rect 9416 29492 9444 29532
rect 9582 29520 9588 29532
rect 9640 29520 9646 29572
rect 10244 29560 10272 29668
rect 10502 29656 10508 29708
rect 10560 29696 10566 29708
rect 10778 29696 10784 29708
rect 10560 29668 10784 29696
rect 10560 29656 10566 29668
rect 10778 29656 10784 29668
rect 10836 29656 10842 29708
rect 11330 29696 11336 29708
rect 11291 29668 11336 29696
rect 11330 29656 11336 29668
rect 11388 29656 11394 29708
rect 11716 29696 11744 29736
rect 13446 29724 13452 29776
rect 13504 29764 13510 29776
rect 13722 29764 13728 29776
rect 13504 29736 13728 29764
rect 13504 29724 13510 29736
rect 13722 29724 13728 29736
rect 13780 29724 13786 29776
rect 14384 29764 14412 29804
rect 14844 29773 14872 29804
rect 15562 29792 15568 29844
rect 15620 29832 15626 29844
rect 15838 29832 15844 29844
rect 15620 29804 15844 29832
rect 15620 29792 15626 29804
rect 13832 29736 14412 29764
rect 14829 29767 14887 29773
rect 13832 29696 13860 29736
rect 14829 29733 14841 29767
rect 14875 29733 14887 29767
rect 14829 29727 14887 29733
rect 14921 29767 14979 29773
rect 14921 29733 14933 29767
rect 14967 29764 14979 29767
rect 15286 29764 15292 29776
rect 14967 29736 15292 29764
rect 14967 29733 14979 29736
rect 14921 29727 14979 29733
rect 15286 29724 15292 29736
rect 15344 29724 15350 29776
rect 15562 29696 15568 29708
rect 11716 29668 11836 29696
rect 10410 29628 10416 29640
rect 10371 29600 10416 29628
rect 10410 29588 10416 29600
rect 10468 29588 10474 29640
rect 10870 29628 10876 29640
rect 10831 29600 10876 29628
rect 10870 29588 10876 29600
rect 10928 29588 10934 29640
rect 11054 29588 11060 29640
rect 11112 29628 11118 29640
rect 11808 29637 11836 29668
rect 13363 29668 13860 29696
rect 14752 29668 15568 29696
rect 11517 29631 11575 29637
rect 11517 29628 11529 29631
rect 11112 29600 11529 29628
rect 11112 29588 11118 29600
rect 11517 29597 11529 29600
rect 11563 29597 11575 29631
rect 11517 29591 11575 29597
rect 11609 29631 11667 29637
rect 11609 29597 11621 29631
rect 11655 29597 11667 29631
rect 11609 29591 11667 29597
rect 11793 29631 11851 29637
rect 11793 29597 11805 29631
rect 11839 29597 11851 29631
rect 11793 29591 11851 29597
rect 10778 29560 10784 29572
rect 10244 29532 10784 29560
rect 10778 29520 10784 29532
rect 10836 29520 10842 29572
rect 9795 29495 9853 29501
rect 9795 29492 9807 29495
rect 9416 29464 9807 29492
rect 9795 29461 9807 29464
rect 9841 29492 9853 29495
rect 9950 29492 9956 29504
rect 9841 29464 9956 29492
rect 9841 29461 9853 29464
rect 9795 29455 9853 29461
rect 9950 29452 9956 29464
rect 10008 29452 10014 29504
rect 10318 29452 10324 29504
rect 10376 29492 10382 29504
rect 10505 29495 10563 29501
rect 10505 29492 10517 29495
rect 10376 29464 10517 29492
rect 10376 29452 10382 29464
rect 10505 29461 10517 29464
rect 10551 29461 10563 29495
rect 10505 29455 10563 29461
rect 10594 29452 10600 29504
rect 10652 29492 10658 29504
rect 11624 29492 11652 29591
rect 11882 29588 11888 29640
rect 11940 29628 11946 29640
rect 11940 29600 11985 29628
rect 11940 29588 11946 29600
rect 12158 29588 12164 29640
rect 12216 29628 12222 29640
rect 12345 29631 12403 29637
rect 12345 29628 12357 29631
rect 12216 29600 12357 29628
rect 12216 29588 12222 29600
rect 12345 29597 12357 29600
rect 12391 29597 12403 29631
rect 12345 29591 12403 29597
rect 12434 29520 12440 29572
rect 12492 29560 12498 29572
rect 12590 29563 12648 29569
rect 12590 29560 12602 29563
rect 12492 29532 12602 29560
rect 12492 29520 12498 29532
rect 12590 29529 12602 29532
rect 12636 29529 12648 29563
rect 12590 29523 12648 29529
rect 12986 29520 12992 29572
rect 13044 29560 13050 29572
rect 13363 29560 13391 29668
rect 14752 29637 14780 29668
rect 15562 29656 15568 29668
rect 15620 29656 15626 29708
rect 15672 29705 15700 29804
rect 15838 29792 15844 29804
rect 15896 29792 15902 29844
rect 16390 29792 16396 29844
rect 16448 29832 16454 29844
rect 20438 29832 20444 29844
rect 16448 29804 20444 29832
rect 16448 29792 16454 29804
rect 20438 29792 20444 29804
rect 20496 29792 20502 29844
rect 26421 29835 26479 29841
rect 26421 29832 26433 29835
rect 20539 29804 26433 29832
rect 17034 29764 17040 29776
rect 16995 29736 17040 29764
rect 17034 29724 17040 29736
rect 17092 29724 17098 29776
rect 18782 29724 18788 29776
rect 18840 29764 18846 29776
rect 20539 29764 20567 29804
rect 26421 29801 26433 29804
rect 26467 29801 26479 29835
rect 26421 29795 26479 29801
rect 21266 29764 21272 29776
rect 18840 29736 20567 29764
rect 20732 29736 21272 29764
rect 18840 29724 18846 29736
rect 15657 29699 15715 29705
rect 15657 29665 15669 29699
rect 15703 29665 15715 29699
rect 15657 29659 15715 29665
rect 17310 29656 17316 29708
rect 17368 29696 17374 29708
rect 17497 29699 17555 29705
rect 17497 29696 17509 29699
rect 17368 29668 17509 29696
rect 17368 29656 17374 29668
rect 17497 29665 17509 29668
rect 17543 29665 17555 29699
rect 17497 29659 17555 29665
rect 18690 29656 18696 29708
rect 18748 29696 18754 29708
rect 19426 29696 19432 29708
rect 18748 29668 19432 29696
rect 18748 29656 18754 29668
rect 19426 29656 19432 29668
rect 19484 29656 19490 29708
rect 19610 29656 19616 29708
rect 19668 29696 19674 29708
rect 20732 29696 20760 29736
rect 21266 29724 21272 29736
rect 21324 29724 21330 29776
rect 23382 29764 23388 29776
rect 22756 29736 23388 29764
rect 19668 29668 20760 29696
rect 19668 29656 19674 29668
rect 20806 29656 20812 29708
rect 20864 29696 20870 29708
rect 20864 29668 21220 29696
rect 20864 29656 20870 29668
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29597 14795 29631
rect 15010 29628 15016 29640
rect 14923 29600 15016 29628
rect 14737 29591 14795 29597
rect 15010 29588 15016 29600
rect 15068 29588 15074 29640
rect 15378 29588 15384 29640
rect 15436 29628 15442 29640
rect 16482 29628 16488 29640
rect 15436 29600 16488 29628
rect 15436 29588 15442 29600
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 17402 29588 17408 29640
rect 17460 29628 17466 29640
rect 17764 29631 17822 29637
rect 17460 29622 17724 29628
rect 17764 29622 17776 29631
rect 17460 29600 17776 29622
rect 17460 29588 17466 29600
rect 17696 29597 17776 29600
rect 17810 29597 17822 29631
rect 17696 29594 17822 29597
rect 17764 29591 17822 29594
rect 18046 29588 18052 29640
rect 18104 29628 18110 29640
rect 19702 29628 19708 29640
rect 18104 29600 19708 29628
rect 18104 29588 18110 29600
rect 19702 29588 19708 29600
rect 19760 29588 19766 29640
rect 19886 29588 19892 29640
rect 19944 29628 19950 29640
rect 20257 29631 20315 29637
rect 20257 29628 20269 29631
rect 19944 29600 20269 29628
rect 19944 29588 19950 29600
rect 20257 29597 20269 29600
rect 20303 29597 20315 29631
rect 20257 29591 20315 29597
rect 20533 29631 20591 29637
rect 20533 29597 20545 29631
rect 20579 29628 20591 29631
rect 21082 29628 21088 29640
rect 20579 29600 21088 29628
rect 20579 29597 20591 29600
rect 20533 29591 20591 29597
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 21192 29628 21220 29668
rect 22106 29631 22164 29637
rect 22106 29628 22118 29631
rect 21192 29600 22118 29628
rect 22106 29597 22118 29600
rect 22152 29597 22164 29631
rect 22370 29628 22376 29640
rect 22331 29600 22376 29628
rect 22106 29591 22164 29597
rect 22370 29588 22376 29600
rect 22428 29588 22434 29640
rect 13044 29532 13391 29560
rect 13044 29520 13050 29532
rect 13998 29520 14004 29572
rect 14056 29560 14062 29572
rect 14826 29560 14832 29572
rect 14056 29532 14832 29560
rect 14056 29520 14062 29532
rect 14826 29520 14832 29532
rect 14884 29520 14890 29572
rect 15028 29560 15056 29588
rect 15746 29560 15752 29572
rect 15028 29532 15752 29560
rect 15746 29520 15752 29532
rect 15804 29520 15810 29572
rect 15924 29563 15982 29569
rect 15924 29529 15936 29563
rect 15970 29560 15982 29563
rect 18138 29560 18144 29572
rect 15970 29532 18144 29560
rect 15970 29529 15982 29532
rect 15924 29523 15982 29529
rect 18138 29520 18144 29532
rect 18196 29520 18202 29572
rect 18322 29520 18328 29572
rect 18380 29560 18386 29572
rect 20162 29560 20168 29572
rect 18380 29532 20168 29560
rect 18380 29520 18386 29532
rect 20162 29520 20168 29532
rect 20220 29520 20226 29572
rect 20438 29520 20444 29572
rect 20496 29560 20502 29572
rect 20496 29532 22160 29560
rect 20496 29520 20502 29532
rect 14642 29492 14648 29504
rect 10652 29464 10697 29492
rect 11624 29464 14648 29492
rect 10652 29452 10658 29464
rect 14642 29452 14648 29464
rect 14700 29452 14706 29504
rect 15197 29495 15255 29501
rect 15197 29461 15209 29495
rect 15243 29492 15255 29495
rect 16942 29492 16948 29504
rect 15243 29464 16948 29492
rect 15243 29461 15255 29464
rect 15197 29455 15255 29461
rect 16942 29452 16948 29464
rect 17000 29452 17006 29504
rect 17954 29452 17960 29504
rect 18012 29492 18018 29504
rect 18506 29492 18512 29504
rect 18012 29464 18512 29492
rect 18012 29452 18018 29464
rect 18506 29452 18512 29464
rect 18564 29452 18570 29504
rect 18690 29452 18696 29504
rect 18748 29492 18754 29504
rect 18877 29495 18935 29501
rect 18877 29492 18889 29495
rect 18748 29464 18889 29492
rect 18748 29452 18754 29464
rect 18877 29461 18889 29464
rect 18923 29461 18935 29495
rect 18877 29455 18935 29461
rect 20993 29495 21051 29501
rect 20993 29461 21005 29495
rect 21039 29492 21051 29495
rect 21082 29492 21088 29504
rect 21039 29464 21088 29492
rect 21039 29461 21051 29464
rect 20993 29455 21051 29461
rect 21082 29452 21088 29464
rect 21140 29452 21146 29504
rect 22132 29492 22160 29532
rect 22756 29492 22784 29736
rect 23382 29724 23388 29736
rect 23440 29724 23446 29776
rect 23400 29696 23428 29724
rect 22848 29668 23336 29696
rect 23400 29668 24716 29696
rect 22848 29637 22876 29668
rect 22833 29631 22891 29637
rect 22833 29597 22845 29631
rect 22879 29597 22891 29631
rect 22833 29591 22891 29597
rect 22922 29588 22928 29640
rect 22980 29628 22986 29640
rect 23109 29631 23167 29637
rect 23109 29628 23121 29631
rect 22980 29600 23121 29628
rect 22980 29588 22986 29600
rect 23109 29597 23121 29600
rect 23155 29597 23167 29631
rect 23308 29628 23336 29668
rect 24118 29628 24124 29640
rect 23308 29600 24124 29628
rect 23109 29591 23167 29597
rect 22132 29464 22784 29492
rect 23124 29492 23152 29591
rect 24118 29588 24124 29600
rect 24176 29588 24182 29640
rect 24581 29631 24639 29637
rect 24581 29597 24593 29631
rect 24627 29597 24639 29631
rect 24688 29628 24716 29668
rect 24837 29631 24895 29637
rect 24837 29628 24849 29631
rect 24688 29600 24849 29628
rect 24581 29591 24639 29597
rect 24837 29597 24849 29600
rect 24883 29597 24895 29631
rect 24837 29591 24895 29597
rect 23842 29520 23848 29572
rect 23900 29560 23906 29572
rect 24596 29560 24624 29591
rect 25958 29588 25964 29640
rect 26016 29628 26022 29640
rect 27801 29631 27859 29637
rect 27801 29628 27813 29631
rect 26016 29600 27813 29628
rect 26016 29588 26022 29600
rect 27801 29597 27813 29600
rect 27847 29628 27859 29631
rect 28258 29628 28264 29640
rect 27847 29600 28264 29628
rect 27847 29597 27859 29600
rect 27801 29591 27859 29597
rect 28258 29588 28264 29600
rect 28316 29628 28322 29640
rect 28626 29628 28632 29640
rect 28316 29600 28632 29628
rect 28316 29588 28322 29600
rect 28626 29588 28632 29600
rect 28684 29588 28690 29640
rect 23900 29532 24624 29560
rect 23900 29520 23906 29532
rect 25130 29520 25136 29572
rect 25188 29560 25194 29572
rect 27534 29563 27592 29569
rect 27534 29560 27546 29563
rect 25188 29532 27546 29560
rect 25188 29520 25194 29532
rect 27534 29529 27546 29532
rect 27580 29529 27592 29563
rect 27534 29523 27592 29529
rect 24670 29492 24676 29504
rect 23124 29464 24676 29492
rect 24670 29452 24676 29464
rect 24728 29452 24734 29504
rect 25038 29452 25044 29504
rect 25096 29492 25102 29504
rect 25961 29495 26019 29501
rect 25961 29492 25973 29495
rect 25096 29464 25973 29492
rect 25096 29452 25102 29464
rect 25961 29461 25973 29464
rect 26007 29461 26019 29495
rect 25961 29455 26019 29461
rect 27982 29452 27988 29504
rect 28040 29492 28046 29504
rect 28261 29495 28319 29501
rect 28261 29492 28273 29495
rect 28040 29464 28273 29492
rect 28040 29452 28046 29464
rect 28261 29461 28273 29464
rect 28307 29461 28319 29495
rect 28261 29455 28319 29461
rect 1104 29402 29048 29424
rect 1104 29350 7896 29402
rect 7948 29350 7960 29402
rect 8012 29350 8024 29402
rect 8076 29350 8088 29402
rect 8140 29350 8152 29402
rect 8204 29350 14842 29402
rect 14894 29350 14906 29402
rect 14958 29350 14970 29402
rect 15022 29350 15034 29402
rect 15086 29350 15098 29402
rect 15150 29350 21788 29402
rect 21840 29350 21852 29402
rect 21904 29350 21916 29402
rect 21968 29350 21980 29402
rect 22032 29350 22044 29402
rect 22096 29350 28734 29402
rect 28786 29350 28798 29402
rect 28850 29350 28862 29402
rect 28914 29350 28926 29402
rect 28978 29350 28990 29402
rect 29042 29350 29048 29402
rect 1104 29328 29048 29350
rect 5258 29248 5264 29300
rect 5316 29288 5322 29300
rect 6733 29291 6791 29297
rect 6733 29288 6745 29291
rect 5316 29260 6745 29288
rect 5316 29248 5322 29260
rect 6733 29257 6745 29260
rect 6779 29257 6791 29291
rect 6733 29251 6791 29257
rect 6748 29152 6776 29251
rect 6914 29248 6920 29300
rect 6972 29288 6978 29300
rect 7837 29291 7895 29297
rect 7837 29288 7849 29291
rect 6972 29260 7849 29288
rect 6972 29248 6978 29260
rect 7837 29257 7849 29260
rect 7883 29257 7895 29291
rect 8478 29288 8484 29300
rect 8439 29260 8484 29288
rect 7837 29251 7895 29257
rect 7852 29220 7880 29251
rect 8478 29248 8484 29260
rect 8536 29248 8542 29300
rect 8754 29248 8760 29300
rect 8812 29288 8818 29300
rect 9858 29288 9864 29300
rect 8812 29260 9864 29288
rect 8812 29248 8818 29260
rect 9858 29248 9864 29260
rect 9916 29248 9922 29300
rect 16574 29288 16580 29300
rect 10796 29260 16580 29288
rect 9490 29220 9496 29232
rect 7852 29192 9496 29220
rect 9490 29180 9496 29192
rect 9548 29180 9554 29232
rect 10686 29220 10692 29232
rect 9600 29192 10692 29220
rect 9600 29152 9628 29192
rect 10686 29180 10692 29192
rect 10744 29180 10750 29232
rect 10796 29229 10824 29260
rect 16574 29248 16580 29260
rect 16632 29248 16638 29300
rect 17144 29260 17448 29288
rect 10781 29223 10839 29229
rect 10781 29189 10793 29223
rect 10827 29189 10839 29223
rect 10981 29223 11039 29229
rect 10981 29220 10993 29223
rect 10781 29183 10839 29189
rect 10888 29192 10993 29220
rect 6748 29124 9628 29152
rect 9858 29112 9864 29164
rect 9916 29152 9922 29164
rect 10137 29155 10195 29161
rect 10137 29152 10149 29155
rect 9916 29124 10149 29152
rect 9916 29112 9922 29124
rect 10137 29121 10149 29124
rect 10183 29152 10195 29155
rect 10502 29152 10508 29164
rect 10183 29124 10508 29152
rect 10183 29121 10195 29124
rect 10137 29115 10195 29121
rect 10502 29112 10508 29124
rect 10560 29112 10566 29164
rect 10704 29152 10732 29180
rect 10888 29152 10916 29192
rect 10981 29189 10993 29192
rect 11027 29189 11039 29223
rect 10981 29183 11039 29189
rect 12158 29180 12164 29232
rect 12216 29220 12222 29232
rect 12216 29192 13124 29220
rect 12216 29180 12222 29192
rect 12250 29152 12256 29164
rect 10704 29124 10916 29152
rect 12211 29124 12256 29152
rect 12250 29112 12256 29124
rect 12308 29112 12314 29164
rect 12434 29161 12440 29164
rect 12418 29155 12440 29161
rect 12418 29121 12430 29155
rect 12418 29115 12440 29121
rect 12434 29112 12440 29115
rect 12492 29112 12498 29164
rect 12529 29155 12587 29161
rect 12529 29121 12541 29155
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 7377 29087 7435 29093
rect 7377 29053 7389 29087
rect 7423 29084 7435 29087
rect 12544 29084 12572 29115
rect 12618 29112 12624 29164
rect 12676 29152 12682 29164
rect 13096 29161 13124 29192
rect 13538 29180 13544 29232
rect 13596 29220 13602 29232
rect 15010 29220 15016 29232
rect 13596 29192 15016 29220
rect 13596 29180 13602 29192
rect 15010 29180 15016 29192
rect 15068 29180 15074 29232
rect 15378 29220 15384 29232
rect 15120 29192 15384 29220
rect 13081 29155 13139 29161
rect 12676 29124 12721 29152
rect 12676 29112 12682 29124
rect 13081 29121 13093 29155
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13348 29155 13406 29161
rect 13348 29121 13360 29155
rect 13394 29152 13406 29155
rect 14458 29152 14464 29164
rect 13394 29124 14464 29152
rect 13394 29121 13406 29124
rect 13348 29115 13406 29121
rect 14458 29112 14464 29124
rect 14516 29112 14522 29164
rect 15120 29152 15148 29192
rect 15378 29180 15384 29192
rect 15436 29180 15442 29232
rect 15470 29180 15476 29232
rect 15528 29220 15534 29232
rect 15528 29192 16068 29220
rect 15528 29180 15534 29192
rect 14936 29124 15148 29152
rect 15188 29155 15246 29161
rect 7423 29056 13124 29084
rect 7423 29053 7435 29056
rect 7377 29047 7435 29053
rect 13096 29028 13124 29056
rect 14734 29044 14740 29096
rect 14792 29084 14798 29096
rect 14936 29093 14964 29124
rect 15188 29121 15200 29155
rect 15234 29152 15246 29155
rect 15746 29152 15752 29164
rect 15234 29124 15752 29152
rect 15234 29121 15246 29124
rect 15188 29115 15246 29121
rect 15746 29112 15752 29124
rect 15804 29112 15810 29164
rect 16040 29152 16068 29192
rect 16758 29180 16764 29232
rect 16816 29220 16822 29232
rect 17144 29220 17172 29260
rect 17420 29229 17448 29260
rect 18340 29260 18532 29288
rect 16816 29192 17172 29220
rect 17405 29223 17463 29229
rect 16816 29180 16822 29192
rect 17405 29189 17417 29223
rect 17451 29189 17463 29223
rect 17405 29183 17463 29189
rect 17635 29223 17693 29229
rect 17635 29189 17647 29223
rect 17681 29220 17693 29223
rect 18340 29220 18368 29260
rect 17681 29192 18368 29220
rect 18504 29220 18532 29260
rect 18874 29248 18880 29300
rect 18932 29288 18938 29300
rect 20438 29288 20444 29300
rect 18932 29260 20444 29288
rect 18932 29248 18938 29260
rect 20438 29248 20444 29260
rect 20496 29248 20502 29300
rect 21082 29288 21088 29300
rect 20916 29260 21088 29288
rect 20714 29220 20720 29232
rect 18504 29192 20720 29220
rect 17681 29189 17693 29192
rect 17635 29183 17693 29189
rect 20714 29180 20720 29192
rect 20772 29180 20778 29232
rect 17129 29155 17187 29161
rect 17129 29152 17141 29155
rect 16040 29124 17141 29152
rect 17129 29121 17141 29124
rect 17175 29121 17187 29155
rect 17310 29152 17316 29164
rect 17271 29124 17316 29152
rect 17129 29115 17187 29121
rect 17310 29112 17316 29124
rect 17368 29112 17374 29164
rect 17494 29152 17500 29164
rect 17455 29124 17500 29152
rect 17494 29112 17500 29124
rect 17552 29112 17558 29164
rect 17954 29112 17960 29164
rect 18012 29152 18018 29164
rect 18233 29155 18291 29161
rect 18233 29152 18245 29155
rect 18012 29124 18245 29152
rect 18012 29112 18018 29124
rect 18233 29121 18245 29124
rect 18279 29121 18291 29155
rect 18500 29155 18558 29161
rect 18500 29152 18512 29155
rect 18233 29115 18291 29121
rect 18340 29124 18512 29152
rect 14921 29087 14979 29093
rect 14921 29084 14933 29087
rect 14792 29056 14933 29084
rect 14792 29044 14798 29056
rect 14921 29053 14933 29056
rect 14967 29053 14979 29087
rect 14921 29047 14979 29053
rect 16942 29044 16948 29096
rect 17000 29084 17006 29096
rect 17773 29087 17831 29093
rect 17773 29084 17785 29087
rect 17000 29056 17785 29084
rect 17000 29044 17006 29056
rect 17773 29053 17785 29056
rect 17819 29053 17831 29087
rect 17773 29047 17831 29053
rect 18046 29044 18052 29096
rect 18104 29084 18110 29096
rect 18340 29084 18368 29124
rect 18500 29121 18512 29124
rect 18546 29152 18558 29155
rect 18782 29152 18788 29164
rect 18546 29124 18788 29152
rect 18546 29121 18558 29124
rect 18500 29115 18558 29121
rect 18782 29112 18788 29124
rect 18840 29112 18846 29164
rect 18874 29112 18880 29164
rect 18932 29152 18938 29164
rect 20916 29152 20944 29260
rect 21082 29248 21088 29260
rect 21140 29248 21146 29300
rect 21266 29248 21272 29300
rect 21324 29288 21330 29300
rect 25130 29288 25136 29300
rect 21324 29260 25136 29288
rect 21324 29248 21330 29260
rect 25130 29248 25136 29260
rect 25188 29248 25194 29300
rect 26878 29248 26884 29300
rect 26936 29288 26942 29300
rect 27157 29291 27215 29297
rect 27157 29288 27169 29291
rect 26936 29260 27169 29288
rect 26936 29248 26942 29260
rect 27157 29257 27169 29260
rect 27203 29257 27215 29291
rect 27157 29251 27215 29257
rect 20990 29180 20996 29232
rect 21048 29220 21054 29232
rect 24090 29223 24148 29229
rect 24090 29220 24102 29223
rect 21048 29192 24102 29220
rect 21048 29180 21054 29192
rect 24090 29189 24102 29192
rect 24136 29189 24148 29223
rect 24090 29183 24148 29189
rect 24762 29180 24768 29232
rect 24820 29220 24826 29232
rect 27433 29223 27491 29229
rect 27433 29220 27445 29223
rect 24820 29192 27445 29220
rect 24820 29180 24826 29192
rect 27433 29189 27445 29192
rect 27479 29189 27491 29223
rect 27433 29183 27491 29189
rect 21186 29155 21244 29161
rect 21186 29152 21198 29155
rect 18932 29124 21198 29152
rect 18932 29112 18938 29124
rect 21186 29121 21198 29124
rect 21232 29121 21244 29155
rect 21186 29115 21244 29121
rect 23106 29112 23112 29164
rect 23164 29161 23170 29164
rect 23164 29152 23176 29161
rect 23164 29124 24900 29152
rect 23164 29115 23176 29124
rect 23164 29112 23170 29115
rect 18104 29056 18368 29084
rect 21453 29087 21511 29093
rect 18104 29044 18110 29056
rect 21453 29053 21465 29087
rect 21499 29084 21511 29087
rect 22370 29084 22376 29096
rect 21499 29056 22376 29084
rect 21499 29053 21511 29056
rect 21453 29047 21511 29053
rect 22370 29044 22376 29056
rect 22428 29044 22434 29096
rect 23382 29084 23388 29096
rect 23343 29056 23388 29084
rect 23382 29044 23388 29056
rect 23440 29084 23446 29096
rect 23842 29084 23848 29096
rect 23440 29056 23848 29084
rect 23440 29044 23446 29056
rect 23842 29044 23848 29056
rect 23900 29044 23906 29096
rect 5997 29019 6055 29025
rect 5997 28985 6009 29019
rect 6043 29016 6055 29019
rect 8938 29016 8944 29028
rect 6043 28988 8616 29016
rect 8899 28988 8944 29016
rect 6043 28985 6055 28988
rect 5997 28979 6055 28985
rect 8588 28948 8616 28988
rect 8938 28976 8944 28988
rect 8996 28976 9002 29028
rect 11054 29016 11060 29028
rect 10244 28988 11060 29016
rect 8754 28948 8760 28960
rect 8588 28920 8760 28948
rect 8754 28908 8760 28920
rect 8812 28908 8818 28960
rect 9214 28908 9220 28960
rect 9272 28948 9278 28960
rect 10244 28957 10272 28988
rect 11054 28976 11060 28988
rect 11112 28976 11118 29028
rect 11149 29019 11207 29025
rect 11149 28985 11161 29019
rect 11195 29016 11207 29019
rect 12986 29016 12992 29028
rect 11195 28988 12992 29016
rect 11195 28985 11207 28988
rect 11149 28979 11207 28985
rect 12986 28976 12992 28988
rect 13044 28976 13050 29028
rect 13078 28976 13084 29028
rect 13136 28976 13142 29028
rect 16758 29016 16764 29028
rect 14384 28988 14688 29016
rect 9493 28951 9551 28957
rect 9493 28948 9505 28951
rect 9272 28920 9505 28948
rect 9272 28908 9278 28920
rect 9493 28917 9505 28920
rect 9539 28948 9551 28951
rect 10229 28951 10287 28957
rect 10229 28948 10241 28951
rect 9539 28920 10241 28948
rect 9539 28917 9551 28920
rect 9493 28911 9551 28917
rect 10229 28917 10241 28920
rect 10275 28917 10287 28951
rect 10229 28911 10287 28917
rect 10594 28908 10600 28960
rect 10652 28948 10658 28960
rect 10962 28948 10968 28960
rect 10652 28920 10968 28948
rect 10652 28908 10658 28920
rect 10962 28908 10968 28920
rect 11020 28908 11026 28960
rect 11072 28948 11100 28976
rect 11238 28948 11244 28960
rect 11072 28920 11244 28948
rect 11238 28908 11244 28920
rect 11296 28908 11302 28960
rect 12069 28951 12127 28957
rect 12069 28917 12081 28951
rect 12115 28948 12127 28951
rect 14384 28948 14412 28988
rect 12115 28920 14412 28948
rect 12115 28917 12127 28920
rect 12069 28911 12127 28917
rect 14458 28908 14464 28960
rect 14516 28948 14522 28960
rect 14660 28948 14688 28988
rect 16224 28988 16764 29016
rect 16224 28948 16252 28988
rect 16758 28976 16764 28988
rect 16816 28976 16822 29028
rect 20073 29019 20131 29025
rect 20073 29016 20085 29019
rect 17512 28988 18276 29016
rect 14516 28920 14561 28948
rect 14660 28920 16252 28948
rect 16301 28951 16359 28957
rect 14516 28908 14522 28920
rect 16301 28917 16313 28951
rect 16347 28948 16359 28951
rect 16390 28948 16396 28960
rect 16347 28920 16396 28948
rect 16347 28917 16359 28920
rect 16301 28911 16359 28917
rect 16390 28908 16396 28920
rect 16448 28908 16454 28960
rect 16482 28908 16488 28960
rect 16540 28948 16546 28960
rect 17512 28948 17540 28988
rect 16540 28920 17540 28948
rect 18248 28948 18276 28988
rect 19168 28988 20085 29016
rect 19168 28948 19196 28988
rect 20073 28985 20085 28988
rect 20119 29016 20131 29019
rect 20346 29016 20352 29028
rect 20119 28988 20352 29016
rect 20119 28985 20131 28988
rect 20073 28979 20131 28985
rect 20346 28976 20352 28988
rect 20404 28976 20410 29028
rect 21634 28976 21640 29028
rect 21692 29016 21698 29028
rect 22005 29019 22063 29025
rect 22005 29016 22017 29019
rect 21692 28988 22017 29016
rect 21692 28976 21698 28988
rect 22005 28985 22017 28988
rect 22051 28985 22063 29019
rect 22005 28979 22063 28985
rect 18248 28920 19196 28948
rect 16540 28908 16546 28920
rect 19426 28908 19432 28960
rect 19484 28948 19490 28960
rect 19610 28948 19616 28960
rect 19484 28920 19616 28948
rect 19484 28908 19490 28920
rect 19610 28908 19616 28920
rect 19668 28908 19674 28960
rect 19886 28908 19892 28960
rect 19944 28948 19950 28960
rect 20254 28948 20260 28960
rect 19944 28920 20260 28948
rect 19944 28908 19950 28920
rect 20254 28908 20260 28920
rect 20312 28908 20318 28960
rect 20438 28908 20444 28960
rect 20496 28948 20502 28960
rect 23842 28948 23848 28960
rect 20496 28920 23848 28948
rect 20496 28908 20502 28920
rect 23842 28908 23848 28920
rect 23900 28908 23906 28960
rect 24872 28948 24900 29124
rect 27154 29112 27160 29164
rect 27212 29152 27218 29164
rect 27341 29155 27399 29161
rect 27341 29152 27353 29155
rect 27212 29124 27353 29152
rect 27212 29112 27218 29124
rect 27341 29121 27353 29124
rect 27387 29121 27399 29155
rect 27522 29152 27528 29164
rect 27483 29124 27528 29152
rect 27341 29115 27399 29121
rect 27522 29112 27528 29124
rect 27580 29112 27586 29164
rect 27614 29112 27620 29164
rect 27672 29161 27678 29164
rect 27672 29155 27701 29161
rect 27689 29121 27701 29155
rect 27672 29115 27701 29121
rect 27672 29112 27678 29115
rect 27798 29112 27804 29164
rect 27856 29152 27862 29164
rect 27856 29124 27901 29152
rect 27856 29112 27862 29124
rect 25685 29087 25743 29093
rect 25685 29053 25697 29087
rect 25731 29053 25743 29087
rect 25958 29084 25964 29096
rect 25919 29056 25964 29084
rect 25685 29047 25743 29053
rect 24946 28976 24952 29028
rect 25004 29016 25010 29028
rect 25700 29016 25728 29047
rect 25958 29044 25964 29056
rect 26016 29044 26022 29096
rect 26694 29016 26700 29028
rect 25004 28988 26700 29016
rect 25004 28976 25010 28988
rect 26694 28976 26700 28988
rect 26752 29016 26758 29028
rect 26878 29016 26884 29028
rect 26752 28988 26884 29016
rect 26752 28976 26758 28988
rect 26878 28976 26884 28988
rect 26936 28976 26942 29028
rect 25225 28951 25283 28957
rect 25225 28948 25237 28951
rect 24872 28920 25237 28948
rect 25225 28917 25237 28920
rect 25271 28917 25283 28951
rect 28350 28948 28356 28960
rect 28311 28920 28356 28948
rect 25225 28911 25283 28917
rect 28350 28908 28356 28920
rect 28408 28948 28414 28960
rect 28626 28948 28632 28960
rect 28408 28920 28632 28948
rect 28408 28908 28414 28920
rect 28626 28908 28632 28920
rect 28684 28908 28690 28960
rect 1104 28858 28888 28880
rect 1104 28806 4423 28858
rect 4475 28806 4487 28858
rect 4539 28806 4551 28858
rect 4603 28806 4615 28858
rect 4667 28806 4679 28858
rect 4731 28806 11369 28858
rect 11421 28806 11433 28858
rect 11485 28806 11497 28858
rect 11549 28806 11561 28858
rect 11613 28806 11625 28858
rect 11677 28806 18315 28858
rect 18367 28806 18379 28858
rect 18431 28806 18443 28858
rect 18495 28806 18507 28858
rect 18559 28806 18571 28858
rect 18623 28806 25261 28858
rect 25313 28806 25325 28858
rect 25377 28806 25389 28858
rect 25441 28806 25453 28858
rect 25505 28806 25517 28858
rect 25569 28806 28888 28858
rect 1104 28784 28888 28806
rect 6365 28747 6423 28753
rect 6365 28713 6377 28747
rect 6411 28744 6423 28747
rect 8386 28744 8392 28756
rect 6411 28716 8392 28744
rect 6411 28713 6423 28716
rect 6365 28707 6423 28713
rect 8386 28704 8392 28716
rect 8444 28704 8450 28756
rect 8573 28747 8631 28753
rect 8573 28713 8585 28747
rect 8619 28744 8631 28747
rect 8662 28744 8668 28756
rect 8619 28716 8668 28744
rect 8619 28713 8631 28716
rect 8573 28707 8631 28713
rect 8662 28704 8668 28716
rect 8720 28704 8726 28756
rect 9490 28704 9496 28756
rect 9548 28744 9554 28756
rect 10873 28747 10931 28753
rect 10873 28744 10885 28747
rect 9548 28716 10885 28744
rect 9548 28704 9554 28716
rect 10873 28713 10885 28716
rect 10919 28744 10931 28747
rect 11054 28744 11060 28756
rect 10919 28716 11060 28744
rect 10919 28713 10931 28716
rect 10873 28707 10931 28713
rect 11054 28704 11060 28716
rect 11112 28704 11118 28756
rect 11146 28704 11152 28756
rect 11204 28744 11210 28756
rect 11606 28744 11612 28756
rect 11204 28716 11612 28744
rect 11204 28704 11210 28716
rect 11606 28704 11612 28716
rect 11664 28704 11670 28756
rect 11793 28747 11851 28753
rect 11793 28713 11805 28747
rect 11839 28744 11851 28747
rect 13170 28744 13176 28756
rect 11839 28716 13176 28744
rect 11839 28713 11851 28716
rect 11793 28707 11851 28713
rect 13170 28704 13176 28716
rect 13228 28704 13234 28756
rect 14645 28747 14703 28753
rect 14645 28713 14657 28747
rect 14691 28744 14703 28747
rect 20070 28744 20076 28756
rect 14691 28716 20076 28744
rect 14691 28713 14703 28716
rect 14645 28707 14703 28713
rect 20070 28704 20076 28716
rect 20128 28704 20134 28756
rect 20254 28704 20260 28756
rect 20312 28744 20318 28756
rect 23658 28744 23664 28756
rect 20312 28716 23664 28744
rect 20312 28704 20318 28716
rect 23658 28704 23664 28716
rect 23716 28704 23722 28756
rect 23842 28704 23848 28756
rect 23900 28744 23906 28756
rect 25498 28744 25504 28756
rect 23900 28716 25504 28744
rect 23900 28704 23906 28716
rect 25498 28704 25504 28716
rect 25556 28704 25562 28756
rect 6917 28679 6975 28685
rect 6917 28645 6929 28679
rect 6963 28676 6975 28679
rect 7098 28676 7104 28688
rect 6963 28648 7104 28676
rect 6963 28645 6975 28648
rect 6917 28639 6975 28645
rect 7098 28636 7104 28648
rect 7156 28676 7162 28688
rect 7377 28679 7435 28685
rect 7377 28676 7389 28679
rect 7156 28648 7389 28676
rect 7156 28636 7162 28648
rect 7377 28645 7389 28648
rect 7423 28645 7435 28679
rect 7377 28639 7435 28645
rect 7742 28636 7748 28688
rect 7800 28676 7806 28688
rect 7929 28679 7987 28685
rect 7929 28676 7941 28679
rect 7800 28648 7941 28676
rect 7800 28636 7806 28648
rect 7929 28645 7941 28648
rect 7975 28645 7987 28679
rect 8680 28676 8708 28704
rect 9677 28679 9735 28685
rect 9677 28676 9689 28679
rect 8680 28648 9689 28676
rect 7929 28639 7987 28645
rect 9508 28620 9536 28648
rect 9677 28645 9689 28648
rect 9723 28645 9735 28679
rect 11072 28676 11100 28704
rect 12158 28676 12164 28688
rect 11072 28648 12164 28676
rect 9677 28639 9735 28645
rect 12158 28636 12164 28648
rect 12216 28636 12222 28688
rect 14550 28676 14556 28688
rect 13372 28648 14556 28676
rect 9490 28568 9496 28620
rect 9548 28568 9554 28620
rect 11238 28568 11244 28620
rect 11296 28608 11302 28620
rect 13372 28608 13400 28648
rect 14550 28636 14556 28648
rect 14608 28636 14614 28688
rect 15010 28636 15016 28688
rect 15068 28676 15074 28688
rect 15470 28676 15476 28688
rect 15068 28648 15476 28676
rect 15068 28636 15074 28648
rect 15470 28636 15476 28648
rect 15528 28636 15534 28688
rect 16758 28636 16764 28688
rect 16816 28676 16822 28688
rect 17037 28679 17095 28685
rect 17037 28676 17049 28679
rect 16816 28648 17049 28676
rect 16816 28636 16822 28648
rect 17037 28645 17049 28648
rect 17083 28645 17095 28679
rect 19426 28676 19432 28688
rect 17037 28639 17095 28645
rect 18892 28648 19432 28676
rect 13814 28608 13820 28620
rect 11296 28580 13400 28608
rect 11296 28568 11302 28580
rect 1578 28540 1584 28552
rect 1539 28512 1584 28540
rect 1578 28500 1584 28512
rect 1636 28500 1642 28552
rect 8938 28500 8944 28552
rect 8996 28540 9002 28552
rect 10134 28540 10140 28552
rect 8996 28512 10140 28540
rect 8996 28500 9002 28512
rect 10134 28500 10140 28512
rect 10192 28500 10198 28552
rect 10410 28500 10416 28552
rect 10468 28540 10474 28552
rect 12253 28543 12311 28549
rect 12253 28540 12265 28543
rect 10468 28512 12265 28540
rect 10468 28500 10474 28512
rect 12253 28509 12265 28512
rect 12299 28540 12311 28543
rect 12342 28540 12348 28552
rect 12299 28512 12348 28540
rect 12299 28509 12311 28512
rect 12253 28503 12311 28509
rect 12342 28500 12348 28512
rect 12400 28500 12406 28552
rect 12526 28540 12532 28552
rect 12487 28512 12532 28540
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 13372 28549 13400 28580
rect 13648 28580 13820 28608
rect 13648 28549 13676 28580
rect 13814 28568 13820 28580
rect 13872 28608 13878 28620
rect 13872 28580 15056 28608
rect 13872 28568 13878 28580
rect 12713 28543 12771 28549
rect 12713 28509 12725 28543
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28509 13415 28543
rect 13357 28503 13415 28509
rect 13449 28543 13507 28549
rect 13449 28509 13461 28543
rect 13495 28509 13507 28543
rect 13449 28503 13507 28509
rect 13633 28543 13691 28549
rect 13633 28509 13645 28543
rect 13679 28509 13691 28543
rect 13633 28503 13691 28509
rect 9674 28432 9680 28484
rect 9732 28472 9738 28484
rect 10781 28475 10839 28481
rect 10781 28472 10793 28475
rect 9732 28444 10793 28472
rect 9732 28432 9738 28444
rect 10781 28441 10793 28444
rect 10827 28441 10839 28475
rect 11422 28472 11428 28484
rect 11383 28444 11428 28472
rect 10781 28435 10839 28441
rect 11422 28432 11428 28444
rect 11480 28432 11486 28484
rect 11641 28475 11699 28481
rect 11641 28441 11653 28475
rect 11687 28472 11699 28475
rect 11790 28472 11796 28484
rect 11687 28444 11796 28472
rect 11687 28441 11699 28444
rect 11641 28435 11699 28441
rect 11790 28432 11796 28444
rect 11848 28432 11854 28484
rect 12728 28472 12756 28503
rect 13464 28472 13492 28503
rect 13722 28500 13728 28552
rect 13780 28540 13786 28552
rect 13780 28512 13825 28540
rect 13780 28500 13786 28512
rect 14550 28500 14556 28552
rect 14608 28540 14614 28552
rect 14829 28543 14887 28549
rect 14829 28540 14841 28543
rect 14608 28512 14841 28540
rect 14608 28500 14614 28512
rect 14829 28509 14841 28512
rect 14875 28509 14887 28543
rect 14829 28503 14887 28509
rect 14921 28543 14979 28549
rect 14921 28509 14933 28543
rect 14967 28509 14979 28543
rect 15028 28540 15056 28580
rect 15286 28568 15292 28620
rect 15344 28608 15350 28620
rect 15657 28611 15715 28617
rect 15657 28608 15669 28611
rect 15344 28580 15669 28608
rect 15344 28568 15350 28580
rect 15657 28577 15669 28580
rect 15703 28577 15715 28611
rect 15657 28571 15715 28577
rect 16666 28568 16672 28620
rect 16724 28608 16730 28620
rect 17770 28608 17776 28620
rect 16724 28580 17776 28608
rect 16724 28568 16730 28580
rect 17770 28568 17776 28580
rect 17828 28568 17834 28620
rect 18892 28608 18920 28648
rect 19426 28636 19432 28648
rect 19484 28636 19490 28688
rect 20806 28636 20812 28688
rect 20864 28676 20870 28688
rect 20993 28679 21051 28685
rect 20993 28676 21005 28679
rect 20864 28648 21005 28676
rect 20864 28636 20870 28648
rect 20993 28645 21005 28648
rect 21039 28645 21051 28679
rect 20993 28639 21051 28645
rect 22370 28636 22376 28688
rect 22428 28676 22434 28688
rect 22428 28648 23474 28676
rect 22428 28636 22434 28648
rect 19334 28608 19340 28620
rect 18800 28580 18920 28608
rect 18984 28580 19340 28608
rect 15102 28540 15108 28552
rect 15015 28512 15108 28540
rect 14921 28503 14979 28509
rect 15028 28508 15108 28512
rect 13998 28472 14004 28484
rect 12728 28444 13400 28472
rect 13464 28444 14004 28472
rect 11882 28364 11888 28416
rect 11940 28404 11946 28416
rect 12345 28407 12403 28413
rect 12345 28404 12357 28407
rect 11940 28376 12357 28404
rect 11940 28364 11946 28376
rect 12345 28373 12357 28376
rect 12391 28404 12403 28407
rect 13078 28404 13084 28416
rect 12391 28376 13084 28404
rect 12391 28373 12403 28376
rect 12345 28367 12403 28373
rect 13078 28364 13084 28376
rect 13136 28364 13142 28416
rect 13173 28407 13231 28413
rect 13173 28373 13185 28407
rect 13219 28404 13231 28407
rect 13262 28404 13268 28416
rect 13219 28376 13268 28404
rect 13219 28373 13231 28376
rect 13173 28367 13231 28373
rect 13262 28364 13268 28376
rect 13320 28364 13326 28416
rect 13372 28404 13400 28444
rect 13998 28432 14004 28444
rect 14056 28432 14062 28484
rect 14936 28472 14964 28503
rect 15102 28500 15108 28508
rect 15160 28500 15166 28552
rect 15197 28543 15255 28549
rect 15197 28509 15209 28543
rect 15243 28540 15255 28543
rect 15378 28540 15384 28552
rect 15243 28512 15384 28540
rect 15243 28509 15255 28512
rect 15197 28503 15255 28509
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 18621 28543 18679 28549
rect 18621 28540 18633 28543
rect 15478 28534 17882 28540
rect 17972 28534 18633 28540
rect 15478 28512 18633 28534
rect 15478 28472 15506 28512
rect 17854 28506 18000 28512
rect 18621 28509 18633 28512
rect 18667 28540 18679 28543
rect 18800 28540 18828 28580
rect 18667 28512 18828 28540
rect 18877 28543 18935 28549
rect 18667 28509 18679 28512
rect 18621 28503 18679 28509
rect 18877 28509 18889 28543
rect 18923 28540 18935 28543
rect 18984 28540 19012 28580
rect 19334 28568 19340 28580
rect 19392 28568 19398 28620
rect 20438 28608 20444 28620
rect 20399 28580 20444 28608
rect 20438 28568 20444 28580
rect 20496 28568 20502 28620
rect 22287 28580 22539 28608
rect 22287 28540 22315 28580
rect 18923 28512 19012 28540
rect 19076 28512 22315 28540
rect 18923 28509 18935 28512
rect 18877 28503 18935 28509
rect 14936 28444 15506 28472
rect 15924 28475 15982 28481
rect 15924 28441 15936 28475
rect 15970 28472 15982 28475
rect 17586 28472 17592 28484
rect 15970 28444 17592 28472
rect 15970 28441 15982 28444
rect 15924 28435 15982 28441
rect 17586 28432 17592 28444
rect 17644 28432 17650 28484
rect 17770 28432 17776 28484
rect 17828 28472 17834 28484
rect 18506 28472 18512 28484
rect 17828 28444 18512 28472
rect 17828 28432 17834 28444
rect 18506 28432 18512 28444
rect 18564 28432 18570 28484
rect 19076 28472 19104 28512
rect 22370 28500 22376 28552
rect 22428 28540 22434 28552
rect 22428 28512 22473 28540
rect 22428 28500 22434 28512
rect 18636 28444 19104 28472
rect 16114 28404 16120 28416
rect 13372 28376 16120 28404
rect 16114 28364 16120 28376
rect 16172 28364 16178 28416
rect 16298 28364 16304 28416
rect 16356 28404 16362 28416
rect 17497 28407 17555 28413
rect 17497 28404 17509 28407
rect 16356 28376 17509 28404
rect 16356 28364 16362 28376
rect 17497 28373 17509 28376
rect 17543 28404 17555 28407
rect 18636 28404 18664 28444
rect 19242 28432 19248 28484
rect 19300 28472 19306 28484
rect 22002 28472 22008 28484
rect 19300 28444 22008 28472
rect 19300 28432 19306 28444
rect 22002 28432 22008 28444
rect 22060 28432 22066 28484
rect 22128 28475 22186 28481
rect 22128 28441 22140 28475
rect 22174 28472 22186 28475
rect 22278 28472 22284 28484
rect 22174 28444 22284 28472
rect 22174 28441 22186 28444
rect 22128 28435 22186 28441
rect 22278 28432 22284 28444
rect 22336 28432 22342 28484
rect 22511 28472 22539 28580
rect 23106 28568 23112 28620
rect 23164 28608 23170 28620
rect 23164 28580 23209 28608
rect 23164 28568 23170 28580
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28540 22891 28543
rect 22922 28540 22928 28552
rect 22879 28512 22928 28540
rect 22879 28509 22891 28512
rect 22833 28503 22891 28509
rect 22922 28500 22928 28512
rect 22980 28500 22986 28552
rect 23446 28540 23474 28648
rect 24394 28608 24400 28620
rect 23768 28580 24400 28608
rect 23768 28540 23796 28580
rect 24394 28568 24400 28580
rect 24452 28608 24458 28620
rect 24581 28611 24639 28617
rect 24581 28608 24593 28611
rect 24452 28580 24593 28608
rect 24452 28568 24458 28580
rect 24581 28577 24593 28580
rect 24627 28577 24639 28611
rect 24581 28571 24639 28577
rect 23446 28512 23796 28540
rect 24670 28500 24676 28552
rect 24728 28540 24734 28552
rect 25406 28540 25412 28552
rect 24728 28512 25412 28540
rect 24728 28500 24734 28512
rect 25406 28500 25412 28512
rect 25464 28540 25470 28552
rect 26421 28543 26479 28549
rect 26421 28540 26433 28543
rect 25464 28512 26433 28540
rect 25464 28500 25470 28512
rect 26421 28509 26433 28512
rect 26467 28509 26479 28543
rect 26421 28503 26479 28509
rect 24826 28475 24884 28481
rect 24826 28472 24838 28475
rect 22511 28444 24838 28472
rect 24826 28441 24838 28444
rect 24872 28441 24884 28475
rect 24826 28435 24884 28441
rect 26510 28432 26516 28484
rect 26568 28472 26574 28484
rect 26666 28475 26724 28481
rect 26666 28472 26678 28475
rect 26568 28444 26678 28472
rect 26568 28432 26574 28444
rect 26666 28441 26678 28444
rect 26712 28441 26724 28475
rect 26666 28435 26724 28441
rect 17543 28376 18664 28404
rect 17543 28373 17555 28376
rect 17497 28367 17555 28373
rect 18782 28364 18788 28416
rect 18840 28404 18846 28416
rect 19797 28407 19855 28413
rect 19797 28404 19809 28407
rect 18840 28376 19809 28404
rect 18840 28364 18846 28376
rect 19797 28373 19809 28376
rect 19843 28373 19855 28407
rect 20162 28404 20168 28416
rect 20123 28376 20168 28404
rect 19797 28367 19855 28373
rect 20162 28364 20168 28376
rect 20220 28364 20226 28416
rect 20257 28407 20315 28413
rect 20257 28373 20269 28407
rect 20303 28404 20315 28407
rect 20438 28404 20444 28416
rect 20303 28376 20444 28404
rect 20303 28373 20315 28376
rect 20257 28367 20315 28373
rect 20438 28364 20444 28376
rect 20496 28364 20502 28416
rect 21082 28364 21088 28416
rect 21140 28404 21146 28416
rect 24946 28404 24952 28416
rect 21140 28376 24952 28404
rect 21140 28364 21146 28376
rect 24946 28364 24952 28376
rect 25004 28404 25010 28416
rect 25222 28404 25228 28416
rect 25004 28376 25228 28404
rect 25004 28364 25010 28376
rect 25222 28364 25228 28376
rect 25280 28364 25286 28416
rect 25590 28364 25596 28416
rect 25648 28404 25654 28416
rect 25961 28407 26019 28413
rect 25961 28404 25973 28407
rect 25648 28376 25973 28404
rect 25648 28364 25654 28376
rect 25961 28373 25973 28376
rect 26007 28404 26019 28407
rect 26142 28404 26148 28416
rect 26007 28376 26148 28404
rect 26007 28373 26019 28376
rect 25961 28367 26019 28373
rect 26142 28364 26148 28376
rect 26200 28364 26206 28416
rect 27798 28404 27804 28416
rect 27759 28376 27804 28404
rect 27798 28364 27804 28376
rect 27856 28364 27862 28416
rect 28350 28404 28356 28416
rect 28311 28376 28356 28404
rect 28350 28364 28356 28376
rect 28408 28364 28414 28416
rect 1104 28314 29048 28336
rect 1104 28262 7896 28314
rect 7948 28262 7960 28314
rect 8012 28262 8024 28314
rect 8076 28262 8088 28314
rect 8140 28262 8152 28314
rect 8204 28262 14842 28314
rect 14894 28262 14906 28314
rect 14958 28262 14970 28314
rect 15022 28262 15034 28314
rect 15086 28262 15098 28314
rect 15150 28262 21788 28314
rect 21840 28262 21852 28314
rect 21904 28262 21916 28314
rect 21968 28262 21980 28314
rect 22032 28262 22044 28314
rect 22096 28262 28734 28314
rect 28786 28262 28798 28314
rect 28850 28262 28862 28314
rect 28914 28262 28926 28314
rect 28978 28262 28990 28314
rect 29042 28262 29048 28314
rect 1104 28240 29048 28262
rect 7285 28203 7343 28209
rect 7285 28169 7297 28203
rect 7331 28200 7343 28203
rect 9306 28200 9312 28212
rect 7331 28172 9312 28200
rect 7331 28169 7343 28172
rect 7285 28163 7343 28169
rect 9306 28160 9312 28172
rect 9364 28160 9370 28212
rect 10042 28200 10048 28212
rect 10003 28172 10048 28200
rect 10042 28160 10048 28172
rect 10100 28160 10106 28212
rect 10134 28160 10140 28212
rect 10192 28200 10198 28212
rect 10502 28200 10508 28212
rect 10192 28172 10508 28200
rect 10192 28160 10198 28172
rect 10502 28160 10508 28172
rect 10560 28160 10566 28212
rect 11054 28200 11060 28212
rect 11015 28172 11060 28200
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11790 28160 11796 28212
rect 11848 28200 11854 28212
rect 13078 28200 13084 28212
rect 11848 28172 12296 28200
rect 13039 28172 13084 28200
rect 11848 28160 11854 28172
rect 7374 28092 7380 28144
rect 7432 28132 7438 28144
rect 7745 28135 7803 28141
rect 7745 28132 7757 28135
rect 7432 28104 7757 28132
rect 7432 28092 7438 28104
rect 7745 28101 7757 28104
rect 7791 28132 7803 28135
rect 8297 28135 8355 28141
rect 8297 28132 8309 28135
rect 7791 28104 8309 28132
rect 7791 28101 7803 28104
rect 7745 28095 7803 28101
rect 8297 28101 8309 28104
rect 8343 28132 8355 28135
rect 9214 28132 9220 28144
rect 8343 28104 9220 28132
rect 8343 28101 8355 28104
rect 8297 28095 8355 28101
rect 9214 28092 9220 28104
rect 9272 28092 9278 28144
rect 10318 28092 10324 28144
rect 10376 28132 10382 28144
rect 11882 28132 11888 28144
rect 10376 28104 11888 28132
rect 10376 28092 10382 28104
rect 11882 28092 11888 28104
rect 11940 28092 11946 28144
rect 12161 28135 12219 28141
rect 12161 28101 12173 28135
rect 12207 28101 12219 28135
rect 12268 28132 12296 28172
rect 13078 28160 13084 28172
rect 13136 28160 13142 28212
rect 14461 28203 14519 28209
rect 14461 28169 14473 28203
rect 14507 28200 14519 28203
rect 17678 28200 17684 28212
rect 14507 28172 17684 28200
rect 14507 28169 14519 28172
rect 14461 28163 14519 28169
rect 17678 28160 17684 28172
rect 17736 28160 17742 28212
rect 18230 28200 18236 28212
rect 18143 28172 18236 28200
rect 18230 28160 18236 28172
rect 18288 28200 18294 28212
rect 19058 28200 19064 28212
rect 18288 28172 19064 28200
rect 18288 28160 18294 28172
rect 19058 28160 19064 28172
rect 19116 28160 19122 28212
rect 27798 28200 27804 28212
rect 19444 28172 27804 28200
rect 12342 28132 12348 28144
rect 12400 28141 12406 28144
rect 12400 28135 12419 28141
rect 12268 28104 12348 28132
rect 12161 28095 12219 28101
rect 12176 28064 12204 28095
rect 12342 28092 12348 28104
rect 12407 28132 12419 28135
rect 12407 28104 12493 28132
rect 12407 28101 12419 28104
rect 12400 28095 12419 28101
rect 12400 28092 12406 28095
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 15188 28135 15246 28141
rect 15188 28132 15200 28135
rect 14700 28104 15200 28132
rect 14700 28092 14706 28104
rect 15188 28101 15200 28104
rect 15234 28132 15246 28135
rect 16298 28132 16304 28144
rect 15234 28104 16304 28132
rect 15234 28101 15246 28104
rect 15188 28095 15246 28101
rect 16298 28092 16304 28104
rect 16356 28092 16362 28144
rect 17405 28135 17463 28141
rect 17405 28101 17417 28135
rect 17451 28101 17463 28135
rect 17405 28095 17463 28101
rect 17496 28135 17554 28141
rect 17496 28101 17508 28135
rect 17542 28132 17554 28135
rect 17542 28104 19196 28132
rect 17542 28101 17554 28104
rect 17496 28095 17554 28101
rect 12526 28064 12532 28076
rect 12176 28036 12532 28064
rect 12526 28024 12532 28036
rect 12584 28024 12590 28076
rect 12986 28064 12992 28076
rect 12947 28036 12992 28064
rect 12986 28024 12992 28036
rect 13044 28024 13050 28076
rect 13909 28067 13967 28073
rect 13909 28064 13921 28067
rect 13740 28036 13921 28064
rect 6822 27956 6828 28008
rect 6880 27996 6886 28008
rect 8941 27999 8999 28005
rect 8941 27996 8953 27999
rect 6880 27968 8953 27996
rect 6880 27956 6886 27968
rect 8941 27965 8953 27968
rect 8987 27996 8999 27999
rect 11790 27996 11796 28008
rect 8987 27968 11796 27996
rect 8987 27965 8999 27968
rect 8941 27959 8999 27965
rect 11790 27956 11796 27968
rect 11848 27956 11854 28008
rect 11974 27956 11980 28008
rect 12032 27996 12038 28008
rect 12250 27996 12256 28008
rect 12032 27968 12256 27996
rect 12032 27956 12038 27968
rect 12250 27956 12256 27968
rect 12308 27956 12314 28008
rect 13262 27996 13268 28008
rect 13223 27968 13268 27996
rect 13262 27956 13268 27968
rect 13320 27956 13326 28008
rect 13449 27999 13507 28005
rect 13449 27965 13461 27999
rect 13495 27996 13507 27999
rect 13538 27996 13544 28008
rect 13495 27968 13544 27996
rect 13495 27965 13507 27968
rect 13449 27959 13507 27965
rect 13538 27956 13544 27968
rect 13596 27956 13602 28008
rect 11606 27888 11612 27940
rect 11664 27928 11670 27940
rect 13740 27928 13768 28036
rect 13909 28033 13921 28036
rect 13955 28033 13967 28067
rect 13909 28027 13967 28033
rect 14001 28067 14059 28073
rect 14001 28033 14013 28067
rect 14047 28033 14059 28067
rect 14001 28027 14059 28033
rect 14152 28067 14210 28073
rect 14152 28033 14164 28067
rect 14198 28033 14210 28067
rect 14152 28027 14210 28033
rect 14277 28067 14335 28073
rect 14277 28033 14289 28067
rect 14323 28064 14335 28067
rect 14323 28036 14688 28064
rect 14323 28033 14335 28036
rect 14277 28027 14335 28033
rect 14016 27996 14044 28027
rect 14168 27996 14196 28027
rect 14660 28008 14688 28036
rect 14734 28024 14740 28076
rect 14792 28064 14798 28076
rect 14921 28067 14979 28073
rect 14921 28064 14933 28067
rect 14792 28036 14933 28064
rect 14792 28024 14798 28036
rect 14921 28033 14933 28036
rect 14967 28033 14979 28067
rect 14921 28027 14979 28033
rect 16022 28024 16028 28076
rect 16080 28064 16086 28076
rect 17267 28067 17325 28073
rect 17267 28064 17279 28067
rect 16080 28036 17279 28064
rect 16080 28024 16086 28036
rect 17267 28033 17279 28036
rect 17313 28033 17325 28067
rect 17420 28064 17448 28095
rect 17589 28067 17647 28073
rect 17420 28036 17547 28064
rect 17267 28027 17325 28033
rect 17519 28008 17547 28036
rect 17589 28033 17601 28067
rect 17635 28064 17647 28067
rect 17678 28064 17684 28076
rect 17635 28036 17684 28064
rect 17635 28033 17647 28036
rect 17589 28027 17647 28033
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 17770 28024 17776 28076
rect 17828 28064 17834 28076
rect 19058 28064 19064 28076
rect 17828 28036 17873 28064
rect 17972 28036 19064 28064
rect 17828 28024 17834 28036
rect 17972 28008 18000 28036
rect 19058 28024 19064 28036
rect 19116 28024 19122 28076
rect 19168 28064 19196 28104
rect 19242 28092 19248 28144
rect 19300 28132 19306 28144
rect 19346 28135 19404 28141
rect 19346 28132 19358 28135
rect 19300 28104 19358 28132
rect 19300 28092 19306 28104
rect 19346 28101 19358 28104
rect 19392 28132 19404 28135
rect 19444 28132 19472 28172
rect 27798 28160 27804 28172
rect 27856 28160 27862 28212
rect 19392 28104 19472 28132
rect 19392 28101 19404 28104
rect 19346 28095 19404 28101
rect 19518 28092 19524 28144
rect 19576 28132 19582 28144
rect 19978 28132 19984 28144
rect 19576 28104 19984 28132
rect 19576 28092 19582 28104
rect 19978 28092 19984 28104
rect 20036 28092 20042 28144
rect 20806 28092 20812 28144
rect 20864 28132 20870 28144
rect 21174 28132 21180 28144
rect 21232 28141 21238 28144
rect 20864 28104 21180 28132
rect 20864 28092 20870 28104
rect 21174 28092 21180 28104
rect 21232 28095 21244 28141
rect 21232 28092 21238 28095
rect 21726 28092 21732 28144
rect 21784 28132 21790 28144
rect 22738 28132 22744 28144
rect 21784 28104 22744 28132
rect 21784 28092 21790 28104
rect 22738 28092 22744 28104
rect 22796 28092 22802 28144
rect 23032 28104 24256 28132
rect 20254 28064 20260 28076
rect 19168 28036 20260 28064
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 21453 28067 21511 28073
rect 21453 28064 21465 28067
rect 20456 28036 21465 28064
rect 14458 27996 14464 28008
rect 14016 27968 14136 27996
rect 14168 27968 14464 27996
rect 14108 27940 14136 27968
rect 14458 27956 14464 27968
rect 14516 27956 14522 28008
rect 14642 27956 14648 28008
rect 14700 27956 14706 28008
rect 16114 27956 16120 28008
rect 16172 27996 16178 28008
rect 17034 27996 17040 28008
rect 16172 27968 17040 27996
rect 16172 27956 16178 27968
rect 17034 27956 17040 27968
rect 17092 27956 17098 28008
rect 17129 27999 17187 28005
rect 17129 27965 17141 27999
rect 17175 27965 17187 27999
rect 17494 27996 17500 28008
rect 17414 27968 17500 27996
rect 17129 27959 17187 27965
rect 13906 27928 13912 27940
rect 11664 27900 12388 27928
rect 13740 27900 13912 27928
rect 11664 27888 11670 27900
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 8478 27820 8484 27872
rect 8536 27860 8542 27872
rect 9401 27863 9459 27869
rect 9401 27860 9413 27863
rect 8536 27832 9413 27860
rect 8536 27820 8542 27832
rect 9401 27829 9413 27832
rect 9447 27860 9459 27863
rect 10410 27860 10416 27872
rect 9447 27832 10416 27860
rect 9447 27829 9459 27832
rect 9401 27823 9459 27829
rect 10410 27820 10416 27832
rect 10468 27820 10474 27872
rect 10594 27820 10600 27872
rect 10652 27860 10658 27872
rect 12250 27860 12256 27872
rect 10652 27832 12256 27860
rect 10652 27820 10658 27832
rect 12250 27820 12256 27832
rect 12308 27820 12314 27872
rect 12360 27869 12388 27900
rect 13906 27888 13912 27900
rect 13964 27888 13970 27940
rect 14090 27888 14096 27940
rect 14148 27888 14154 27940
rect 14550 27888 14556 27940
rect 14608 27928 14614 27940
rect 14826 27928 14832 27940
rect 14608 27900 14832 27928
rect 14608 27888 14614 27900
rect 14826 27888 14832 27900
rect 14884 27888 14890 27940
rect 12345 27863 12403 27869
rect 12345 27829 12357 27863
rect 12391 27829 12403 27863
rect 12345 27823 12403 27829
rect 12529 27863 12587 27869
rect 12529 27829 12541 27863
rect 12575 27860 12587 27863
rect 13078 27860 13084 27872
rect 12575 27832 13084 27860
rect 12575 27829 12587 27832
rect 12529 27823 12587 27829
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 14918 27820 14924 27872
rect 14976 27860 14982 27872
rect 15930 27860 15936 27872
rect 14976 27832 15936 27860
rect 14976 27820 14982 27832
rect 15930 27820 15936 27832
rect 15988 27820 15994 27872
rect 16301 27863 16359 27869
rect 16301 27829 16313 27863
rect 16347 27860 16359 27863
rect 17034 27860 17040 27872
rect 16347 27832 17040 27860
rect 16347 27829 16359 27832
rect 16301 27823 16359 27829
rect 17034 27820 17040 27832
rect 17092 27820 17098 27872
rect 17144 27860 17172 27959
rect 17494 27956 17500 27968
rect 17552 27996 17558 28008
rect 17954 27996 17960 28008
rect 17552 27968 17960 27996
rect 17552 27956 17558 27968
rect 17954 27956 17960 27968
rect 18012 27956 18018 28008
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27996 19671 27999
rect 19702 27996 19708 28008
rect 19659 27968 19708 27996
rect 19659 27965 19671 27968
rect 19613 27959 19671 27965
rect 19702 27956 19708 27968
rect 19760 27956 19766 28008
rect 19978 27956 19984 28008
rect 20036 27996 20042 28008
rect 20456 27996 20484 28036
rect 21453 28033 21465 28036
rect 21499 28033 21511 28067
rect 21453 28027 21511 28033
rect 20036 27968 20484 27996
rect 21468 27996 21496 28027
rect 21542 28024 21548 28076
rect 21600 28064 21606 28076
rect 23032 28064 23060 28104
rect 21600 28036 23060 28064
rect 23129 28067 23187 28073
rect 21600 28024 21606 28036
rect 23129 28033 23141 28067
rect 23175 28064 23187 28067
rect 23290 28064 23296 28076
rect 23175 28036 23296 28064
rect 23175 28033 23187 28036
rect 23129 28027 23187 28033
rect 23290 28024 23296 28036
rect 23348 28024 23354 28076
rect 23750 28024 23756 28076
rect 23808 28068 23814 28076
rect 23808 28064 23888 28068
rect 24101 28067 24159 28073
rect 24101 28064 24113 28067
rect 23808 28040 24113 28064
rect 23808 28024 23814 28040
rect 23860 28036 24113 28040
rect 24101 28033 24113 28036
rect 24147 28033 24159 28067
rect 24228 28064 24256 28104
rect 24486 28092 24492 28144
rect 24544 28132 24550 28144
rect 25869 28135 25927 28141
rect 25869 28132 25881 28135
rect 24544 28104 25881 28132
rect 24544 28092 24550 28104
rect 25869 28101 25881 28104
rect 25915 28101 25927 28135
rect 25869 28095 25927 28101
rect 26053 28135 26111 28141
rect 26053 28101 26065 28135
rect 26099 28132 26111 28135
rect 26326 28132 26332 28144
rect 26099 28104 26332 28132
rect 26099 28101 26111 28104
rect 26053 28095 26111 28101
rect 26326 28092 26332 28104
rect 26384 28092 26390 28144
rect 26878 28092 26884 28144
rect 26936 28132 26942 28144
rect 27982 28132 27988 28144
rect 26936 28104 27988 28132
rect 26936 28092 26942 28104
rect 27982 28092 27988 28104
rect 28040 28132 28046 28144
rect 28040 28104 28396 28132
rect 28040 28092 28046 28104
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 24228 28036 27169 28064
rect 24101 28027 24159 28033
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 27338 28064 27344 28076
rect 27299 28036 27344 28064
rect 27157 28027 27215 28033
rect 27338 28024 27344 28036
rect 27396 28024 27402 28076
rect 27614 28064 27620 28076
rect 27575 28036 27620 28064
rect 27614 28024 27620 28036
rect 27672 28024 27678 28076
rect 27798 28024 27804 28076
rect 27856 28064 27862 28076
rect 28368 28073 28396 28104
rect 28169 28067 28227 28073
rect 28169 28064 28181 28067
rect 27856 28036 28181 28064
rect 27856 28024 27862 28036
rect 28169 28033 28181 28036
rect 28215 28033 28227 28067
rect 28169 28027 28227 28033
rect 28353 28067 28411 28073
rect 28353 28033 28365 28067
rect 28399 28033 28411 28067
rect 28353 28027 28411 28033
rect 22370 27996 22376 28008
rect 21468 27968 22376 27996
rect 20036 27956 20042 27968
rect 22370 27956 22376 27968
rect 22428 27956 22434 28008
rect 23382 27996 23388 28008
rect 23295 27968 23388 27996
rect 23382 27956 23388 27968
rect 23440 27956 23446 28008
rect 23842 27956 23848 28008
rect 23900 27996 23906 28008
rect 23900 27968 23945 27996
rect 23900 27956 23906 27968
rect 24946 27956 24952 28008
rect 25004 27996 25010 28008
rect 25004 27968 25360 27996
rect 25004 27956 25010 27968
rect 17586 27888 17592 27940
rect 17644 27928 17650 27940
rect 17644 27900 18752 27928
rect 17644 27888 17650 27900
rect 18598 27860 18604 27872
rect 17144 27832 18604 27860
rect 18598 27820 18604 27832
rect 18656 27820 18662 27872
rect 18724 27860 18752 27900
rect 19996 27900 20592 27928
rect 19996 27860 20024 27900
rect 18724 27832 20024 27860
rect 20070 27820 20076 27872
rect 20128 27860 20134 27872
rect 20564 27860 20592 27900
rect 20806 27860 20812 27872
rect 20128 27832 20173 27860
rect 20564 27832 20812 27860
rect 20128 27820 20134 27832
rect 20806 27820 20812 27832
rect 20864 27820 20870 27872
rect 21542 27820 21548 27872
rect 21600 27860 21606 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 21600 27832 22017 27860
rect 21600 27820 21606 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22005 27823 22063 27829
rect 22370 27820 22376 27872
rect 22428 27860 22434 27872
rect 23400 27860 23428 27956
rect 25222 27928 25228 27940
rect 25183 27900 25228 27928
rect 25222 27888 25228 27900
rect 25280 27888 25286 27940
rect 25332 27928 25360 27968
rect 25498 27956 25504 28008
rect 25556 27996 25562 28008
rect 25777 27999 25835 28005
rect 25777 27996 25789 27999
rect 25556 27968 25789 27996
rect 25556 27956 25562 27968
rect 25777 27965 25789 27968
rect 25823 27965 25835 27999
rect 25777 27959 25835 27965
rect 26142 27956 26148 28008
rect 26200 27996 26206 28008
rect 27525 27999 27583 28005
rect 27525 27996 27537 27999
rect 26200 27968 27537 27996
rect 26200 27956 26206 27968
rect 27525 27965 27537 27968
rect 27571 27965 27583 27999
rect 27525 27959 27583 27965
rect 26786 27928 26792 27940
rect 25332 27900 26792 27928
rect 26786 27888 26792 27900
rect 26844 27888 26850 27940
rect 27430 27928 27436 27940
rect 27391 27900 27436 27928
rect 27430 27888 27436 27900
rect 27488 27888 27494 27940
rect 22428 27832 23428 27860
rect 22428 27820 22434 27832
rect 23842 27820 23848 27872
rect 23900 27860 23906 27872
rect 25038 27860 25044 27872
rect 23900 27832 25044 27860
rect 23900 27820 23906 27832
rect 25038 27820 25044 27832
rect 25096 27820 25102 27872
rect 25314 27820 25320 27872
rect 25372 27860 25378 27872
rect 26050 27860 26056 27872
rect 25372 27832 26056 27860
rect 25372 27820 25378 27832
rect 26050 27820 26056 27832
rect 26108 27820 26114 27872
rect 26329 27863 26387 27869
rect 26329 27829 26341 27863
rect 26375 27860 26387 27863
rect 26418 27860 26424 27872
rect 26375 27832 26424 27860
rect 26375 27829 26387 27832
rect 26329 27823 26387 27829
rect 26418 27820 26424 27832
rect 26476 27820 26482 27872
rect 28258 27860 28264 27872
rect 28219 27832 28264 27860
rect 28258 27820 28264 27832
rect 28316 27820 28322 27872
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 7742 27616 7748 27668
rect 7800 27656 7806 27668
rect 8478 27656 8484 27668
rect 7800 27628 8484 27656
rect 7800 27616 7806 27628
rect 8478 27616 8484 27628
rect 8536 27616 8542 27668
rect 9214 27616 9220 27668
rect 9272 27656 9278 27668
rect 10965 27659 11023 27665
rect 10965 27656 10977 27659
rect 9272 27628 10977 27656
rect 9272 27616 9278 27628
rect 10965 27625 10977 27628
rect 11011 27625 11023 27659
rect 12158 27656 12164 27668
rect 10965 27619 11023 27625
rect 11532 27628 11836 27656
rect 12119 27628 12164 27656
rect 9401 27591 9459 27597
rect 9401 27557 9413 27591
rect 9447 27588 9459 27591
rect 9674 27588 9680 27600
rect 9447 27560 9680 27588
rect 9447 27557 9459 27560
rect 9401 27551 9459 27557
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 9953 27591 10011 27597
rect 9953 27557 9965 27591
rect 9999 27588 10011 27591
rect 10318 27588 10324 27600
rect 9999 27560 10324 27588
rect 9999 27557 10011 27560
rect 9953 27551 10011 27557
rect 10318 27548 10324 27560
rect 10376 27548 10382 27600
rect 10502 27548 10508 27600
rect 10560 27588 10566 27600
rect 11532 27588 11560 27628
rect 10560 27560 11560 27588
rect 11609 27591 11667 27597
rect 10560 27548 10566 27560
rect 11609 27557 11621 27591
rect 11655 27588 11667 27591
rect 11698 27588 11704 27600
rect 11655 27560 11704 27588
rect 11655 27557 11667 27560
rect 11609 27551 11667 27557
rect 11698 27548 11704 27560
rect 11756 27548 11762 27600
rect 11808 27588 11836 27628
rect 12158 27616 12164 27628
rect 12216 27616 12222 27668
rect 12250 27616 12256 27668
rect 12308 27656 12314 27668
rect 13541 27659 13599 27665
rect 13541 27656 13553 27659
rect 12308 27628 13553 27656
rect 12308 27616 12314 27628
rect 13541 27625 13553 27628
rect 13587 27625 13599 27659
rect 14734 27656 14740 27668
rect 13541 27619 13599 27625
rect 13786 27628 14740 27656
rect 12802 27588 12808 27600
rect 11808 27560 12808 27588
rect 12802 27548 12808 27560
rect 12860 27588 12866 27600
rect 12897 27591 12955 27597
rect 12897 27588 12909 27591
rect 12860 27560 12909 27588
rect 12860 27548 12866 27560
rect 12897 27557 12909 27560
rect 12943 27588 12955 27591
rect 13786 27588 13814 27628
rect 14734 27616 14740 27628
rect 14792 27616 14798 27668
rect 15657 27659 15715 27665
rect 15657 27656 15669 27659
rect 15120 27628 15669 27656
rect 12943 27560 13814 27588
rect 12943 27557 12955 27560
rect 12897 27551 12955 27557
rect 14366 27548 14372 27600
rect 14424 27588 14430 27600
rect 15120 27588 15148 27628
rect 15657 27625 15669 27628
rect 15703 27656 15715 27659
rect 15930 27656 15936 27668
rect 15703 27628 15936 27656
rect 15703 27625 15715 27628
rect 15657 27619 15715 27625
rect 15930 27616 15936 27628
rect 15988 27616 15994 27668
rect 16022 27616 16028 27668
rect 16080 27616 16086 27668
rect 16298 27616 16304 27668
rect 16356 27656 16362 27668
rect 23842 27656 23848 27668
rect 16356 27628 23848 27656
rect 16356 27616 16362 27628
rect 23842 27616 23848 27628
rect 23900 27616 23906 27668
rect 24854 27616 24860 27668
rect 24912 27656 24918 27668
rect 25682 27656 25688 27668
rect 24912 27628 25688 27656
rect 24912 27616 24918 27628
rect 25682 27616 25688 27628
rect 25740 27616 25746 27668
rect 25866 27616 25872 27668
rect 25924 27656 25930 27668
rect 25961 27659 26019 27665
rect 25961 27656 25973 27659
rect 25924 27628 25973 27656
rect 25924 27616 25930 27628
rect 25961 27625 25973 27628
rect 26007 27625 26019 27659
rect 25961 27619 26019 27625
rect 26050 27616 26056 27668
rect 26108 27656 26114 27668
rect 27801 27659 27859 27665
rect 27801 27656 27813 27659
rect 26108 27628 27813 27656
rect 26108 27616 26114 27628
rect 27801 27625 27813 27628
rect 27847 27656 27859 27659
rect 27890 27656 27896 27668
rect 27847 27628 27896 27656
rect 27847 27625 27859 27628
rect 27801 27619 27859 27625
rect 27890 27616 27896 27628
rect 27948 27616 27954 27668
rect 14424 27560 15148 27588
rect 15197 27591 15255 27597
rect 14424 27548 14430 27560
rect 15197 27557 15209 27591
rect 15243 27588 15255 27591
rect 16040 27588 16068 27616
rect 15243 27560 16068 27588
rect 15243 27557 15255 27560
rect 15197 27551 15255 27557
rect 17126 27548 17132 27600
rect 17184 27588 17190 27600
rect 17678 27588 17684 27600
rect 17184 27560 17684 27588
rect 17184 27548 17190 27560
rect 17678 27548 17684 27560
rect 17736 27548 17742 27600
rect 19058 27548 19064 27600
rect 19116 27588 19122 27600
rect 19886 27588 19892 27600
rect 19116 27560 19892 27588
rect 19116 27548 19122 27560
rect 19886 27548 19892 27560
rect 19944 27588 19950 27600
rect 19944 27560 20300 27588
rect 19944 27548 19950 27560
rect 11330 27480 11336 27532
rect 11388 27520 11394 27532
rect 13538 27520 13544 27532
rect 11388 27492 13544 27520
rect 11388 27480 11394 27492
rect 13538 27480 13544 27492
rect 13596 27480 13602 27532
rect 13814 27480 13820 27532
rect 13872 27520 13878 27532
rect 14550 27520 14556 27532
rect 13872 27492 14556 27520
rect 13872 27480 13878 27492
rect 14550 27480 14556 27492
rect 14608 27520 14614 27532
rect 14608 27492 14780 27520
rect 14608 27480 14614 27492
rect 14752 27461 14780 27492
rect 14826 27480 14832 27532
rect 14884 27520 14890 27532
rect 16022 27520 16028 27532
rect 14884 27492 16028 27520
rect 14884 27480 14890 27492
rect 10505 27455 10563 27461
rect 10505 27421 10517 27455
rect 10551 27452 10563 27455
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 10551 27424 13400 27452
rect 10551 27421 10563 27424
rect 10505 27415 10563 27421
rect 13372 27396 13400 27424
rect 13740 27424 14657 27452
rect 9674 27344 9680 27396
rect 9732 27384 9738 27396
rect 12713 27387 12771 27393
rect 12713 27384 12725 27387
rect 9732 27356 12725 27384
rect 9732 27344 9738 27356
rect 12713 27353 12725 27356
rect 12759 27384 12771 27387
rect 12894 27384 12900 27396
rect 12759 27356 12900 27384
rect 12759 27353 12771 27356
rect 12713 27347 12771 27353
rect 12894 27344 12900 27356
rect 12952 27344 12958 27396
rect 13354 27384 13360 27396
rect 13315 27356 13360 27384
rect 13354 27344 13360 27356
rect 13412 27344 13418 27396
rect 8021 27319 8079 27325
rect 8021 27285 8033 27319
rect 8067 27316 8079 27319
rect 8294 27316 8300 27328
rect 8067 27288 8300 27316
rect 8067 27285 8079 27288
rect 8021 27279 8079 27285
rect 8294 27276 8300 27288
rect 8352 27276 8358 27328
rect 10686 27276 10692 27328
rect 10744 27316 10750 27328
rect 11330 27316 11336 27328
rect 10744 27288 11336 27316
rect 10744 27276 10750 27288
rect 11330 27276 11336 27288
rect 11388 27276 11394 27328
rect 13538 27276 13544 27328
rect 13596 27325 13602 27328
rect 13740 27325 13768 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 14737 27455 14795 27461
rect 14737 27421 14749 27455
rect 14783 27421 14795 27455
rect 14918 27452 14924 27464
rect 14879 27424 14924 27452
rect 14737 27415 14795 27421
rect 14918 27412 14924 27424
rect 14976 27412 14982 27464
rect 15028 27461 15056 27492
rect 16022 27480 16028 27492
rect 16080 27480 16086 27532
rect 19334 27520 19340 27532
rect 16960 27492 17908 27520
rect 15013 27455 15071 27461
rect 15013 27421 15025 27455
rect 15059 27421 15071 27455
rect 15013 27415 15071 27421
rect 15286 27412 15292 27464
rect 15344 27452 15350 27464
rect 16960 27452 16988 27492
rect 15344 27424 16988 27452
rect 17037 27455 17095 27461
rect 15344 27412 15350 27424
rect 17037 27421 17049 27455
rect 17083 27452 17095 27455
rect 17494 27452 17500 27464
rect 17083 27424 17500 27452
rect 17083 27421 17095 27424
rect 17037 27415 17095 27421
rect 17494 27412 17500 27424
rect 17552 27412 17558 27464
rect 17880 27452 17908 27492
rect 18800 27492 19340 27520
rect 18800 27452 18828 27492
rect 19334 27480 19340 27492
rect 19392 27480 19398 27532
rect 17880 27424 18828 27452
rect 18877 27455 18935 27461
rect 18877 27421 18889 27455
rect 18923 27452 18935 27455
rect 19518 27452 19524 27464
rect 18923 27424 19524 27452
rect 18923 27421 18935 27424
rect 18877 27415 18935 27421
rect 19518 27412 19524 27424
rect 19576 27452 19582 27464
rect 19702 27452 19708 27464
rect 19576 27424 19708 27452
rect 19576 27412 19582 27424
rect 19702 27412 19708 27424
rect 19760 27412 19766 27464
rect 20162 27452 20168 27464
rect 20123 27424 20168 27452
rect 20162 27412 20168 27424
rect 20220 27412 20226 27464
rect 20272 27452 20300 27560
rect 20990 27548 20996 27600
rect 21048 27588 21054 27600
rect 21085 27591 21143 27597
rect 21085 27588 21097 27591
rect 21048 27560 21097 27588
rect 21048 27548 21054 27560
rect 21085 27557 21097 27560
rect 21131 27557 21143 27591
rect 21085 27551 21143 27557
rect 22554 27548 22560 27600
rect 22612 27588 22618 27600
rect 23566 27588 23572 27600
rect 22612 27560 23572 27588
rect 22612 27548 22618 27560
rect 20349 27455 20407 27461
rect 20349 27452 20361 27455
rect 20272 27424 20361 27452
rect 20349 27421 20361 27424
rect 20395 27421 20407 27455
rect 20622 27452 20628 27464
rect 20583 27424 20628 27452
rect 20349 27415 20407 27421
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 20714 27412 20720 27464
rect 20772 27452 20778 27464
rect 22370 27452 22376 27464
rect 20772 27424 22376 27452
rect 20772 27412 20778 27424
rect 22370 27412 22376 27424
rect 22428 27452 22434 27464
rect 22940 27461 22968 27560
rect 23566 27548 23572 27560
rect 23624 27548 23630 27600
rect 23492 27492 24716 27520
rect 22465 27455 22523 27461
rect 22465 27452 22477 27455
rect 22428 27424 22477 27452
rect 22428 27412 22434 27424
rect 22465 27421 22477 27424
rect 22511 27421 22523 27455
rect 22465 27415 22523 27421
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27421 22983 27455
rect 22925 27415 22983 27421
rect 23014 27412 23020 27464
rect 23072 27452 23078 27464
rect 23201 27455 23259 27461
rect 23201 27452 23213 27455
rect 23072 27424 23213 27452
rect 23072 27412 23078 27424
rect 23201 27421 23213 27424
rect 23247 27421 23259 27455
rect 23201 27415 23259 27421
rect 23290 27412 23296 27464
rect 23348 27452 23354 27464
rect 23492 27452 23520 27492
rect 23348 27424 23520 27452
rect 23348 27412 23354 27424
rect 23934 27412 23940 27464
rect 23992 27452 23998 27464
rect 24578 27452 24584 27464
rect 23992 27424 24584 27452
rect 23992 27412 23998 27424
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 24688 27452 24716 27492
rect 24688 27424 25084 27452
rect 25056 27396 25084 27424
rect 26050 27412 26056 27464
rect 26108 27452 26114 27464
rect 26421 27455 26479 27461
rect 26421 27452 26433 27455
rect 26108 27424 26433 27452
rect 26108 27412 26114 27424
rect 26421 27421 26433 27424
rect 26467 27421 26479 27455
rect 26421 27415 26479 27421
rect 13814 27344 13820 27396
rect 13872 27384 13878 27396
rect 16114 27384 16120 27396
rect 13872 27356 16120 27384
rect 13872 27344 13878 27356
rect 16114 27344 16120 27356
rect 16172 27344 16178 27396
rect 16792 27387 16850 27393
rect 16792 27353 16804 27387
rect 16838 27384 16850 27387
rect 16942 27384 16948 27396
rect 16838 27356 16948 27384
rect 16838 27353 16850 27356
rect 16792 27347 16850 27353
rect 16942 27344 16948 27356
rect 17000 27344 17006 27396
rect 17126 27344 17132 27396
rect 17184 27384 17190 27396
rect 18632 27387 18690 27393
rect 17184 27356 17882 27384
rect 17184 27344 17190 27356
rect 13596 27319 13615 27325
rect 13603 27285 13615 27319
rect 13596 27279 13615 27285
rect 13725 27319 13783 27325
rect 13725 27285 13737 27319
rect 13771 27285 13783 27319
rect 13725 27279 13783 27285
rect 13596 27276 13602 27279
rect 14182 27276 14188 27328
rect 14240 27316 14246 27328
rect 16666 27316 16672 27328
rect 14240 27288 16672 27316
rect 14240 27276 14246 27288
rect 16666 27276 16672 27288
rect 16724 27316 16730 27328
rect 17497 27319 17555 27325
rect 17497 27316 17509 27319
rect 16724 27288 17509 27316
rect 16724 27276 16730 27288
rect 17497 27285 17509 27288
rect 17543 27285 17555 27319
rect 17854 27316 17882 27356
rect 18632 27353 18644 27387
rect 18678 27384 18690 27387
rect 19058 27384 19064 27396
rect 18678 27356 19064 27384
rect 18678 27353 18690 27356
rect 18632 27347 18690 27353
rect 19058 27344 19064 27356
rect 19116 27344 19122 27396
rect 20257 27387 20315 27393
rect 20257 27384 20269 27387
rect 19168 27356 20269 27384
rect 19168 27316 19196 27356
rect 20257 27353 20269 27356
rect 20303 27353 20315 27387
rect 20257 27347 20315 27353
rect 20487 27387 20545 27393
rect 20487 27353 20499 27387
rect 20533 27384 20545 27387
rect 22220 27387 22278 27393
rect 20533 27356 22094 27384
rect 20533 27353 20545 27356
rect 20487 27347 20545 27353
rect 17854 27288 19196 27316
rect 19521 27319 19579 27325
rect 17497 27279 17555 27285
rect 19521 27285 19533 27319
rect 19567 27316 19579 27319
rect 19702 27316 19708 27328
rect 19567 27288 19708 27316
rect 19567 27285 19579 27288
rect 19521 27279 19579 27285
rect 19702 27276 19708 27288
rect 19760 27276 19766 27328
rect 19981 27319 20039 27325
rect 19981 27285 19993 27319
rect 20027 27316 20039 27319
rect 21726 27316 21732 27328
rect 20027 27288 21732 27316
rect 20027 27285 20039 27288
rect 19981 27279 20039 27285
rect 21726 27276 21732 27288
rect 21784 27276 21790 27328
rect 22066 27316 22094 27356
rect 22220 27353 22232 27387
rect 22266 27384 22278 27387
rect 22646 27384 22652 27396
rect 22266 27356 22652 27384
rect 22266 27353 22278 27356
rect 22220 27347 22278 27353
rect 22646 27344 22652 27356
rect 22704 27344 22710 27396
rect 23382 27344 23388 27396
rect 23440 27384 23446 27396
rect 24837 27387 24895 27393
rect 24837 27384 24849 27387
rect 23440 27356 24849 27384
rect 23440 27344 23446 27356
rect 24837 27353 24849 27356
rect 24883 27353 24895 27387
rect 24837 27347 24895 27353
rect 25038 27344 25044 27396
rect 25096 27344 25102 27396
rect 26666 27387 26724 27393
rect 26666 27353 26678 27387
rect 26712 27384 26724 27387
rect 26786 27384 26792 27396
rect 26712 27356 26792 27384
rect 26712 27353 26724 27356
rect 26666 27347 26724 27353
rect 26786 27344 26792 27356
rect 26844 27344 26850 27396
rect 27062 27344 27068 27396
rect 27120 27384 27126 27396
rect 27890 27384 27896 27396
rect 27120 27356 27896 27384
rect 27120 27344 27126 27356
rect 27890 27344 27896 27356
rect 27948 27344 27954 27396
rect 23566 27316 23572 27328
rect 22066 27288 23572 27316
rect 23566 27276 23572 27288
rect 23624 27276 23630 27328
rect 27338 27276 27344 27328
rect 27396 27316 27402 27328
rect 27522 27316 27528 27328
rect 27396 27288 27528 27316
rect 27396 27276 27402 27288
rect 27522 27276 27528 27288
rect 27580 27276 27586 27328
rect 28350 27316 28356 27328
rect 28311 27288 28356 27316
rect 28350 27276 28356 27288
rect 28408 27276 28414 27328
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 9490 27112 9496 27124
rect 9451 27084 9496 27112
rect 9490 27072 9496 27084
rect 9548 27072 9554 27124
rect 9674 27072 9680 27124
rect 9732 27112 9738 27124
rect 9953 27115 10011 27121
rect 9953 27112 9965 27115
rect 9732 27084 9965 27112
rect 9732 27072 9738 27084
rect 9953 27081 9965 27084
rect 9999 27081 10011 27115
rect 10594 27112 10600 27124
rect 10555 27084 10600 27112
rect 9953 27075 10011 27081
rect 10594 27072 10600 27084
rect 10652 27072 10658 27124
rect 11146 27112 11152 27124
rect 11107 27084 11152 27112
rect 11146 27072 11152 27084
rect 11204 27072 11210 27124
rect 11882 27072 11888 27124
rect 11940 27112 11946 27124
rect 12161 27115 12219 27121
rect 12161 27112 12173 27115
rect 11940 27084 12173 27112
rect 11940 27072 11946 27084
rect 12161 27081 12173 27084
rect 12207 27081 12219 27115
rect 12161 27075 12219 27081
rect 12618 27072 12624 27124
rect 12676 27112 12682 27124
rect 14001 27115 14059 27121
rect 14001 27112 14013 27115
rect 12676 27084 14013 27112
rect 12676 27072 12682 27084
rect 14001 27081 14013 27084
rect 14047 27081 14059 27115
rect 14001 27075 14059 27081
rect 14734 27072 14740 27124
rect 14792 27112 14798 27124
rect 15470 27112 15476 27124
rect 14792 27084 15476 27112
rect 14792 27072 14798 27084
rect 15470 27072 15476 27084
rect 15528 27072 15534 27124
rect 16301 27115 16359 27121
rect 16301 27081 16313 27115
rect 16347 27112 16359 27115
rect 16482 27112 16488 27124
rect 16347 27084 16488 27112
rect 16347 27081 16359 27084
rect 16301 27075 16359 27081
rect 16482 27072 16488 27084
rect 16540 27072 16546 27124
rect 17773 27115 17831 27121
rect 17773 27081 17785 27115
rect 17819 27112 17831 27115
rect 17862 27112 17868 27124
rect 17819 27084 17868 27112
rect 17819 27081 17831 27084
rect 17773 27075 17831 27081
rect 17862 27072 17868 27084
rect 17920 27072 17926 27124
rect 21358 27112 21364 27124
rect 17972 27084 21364 27112
rect 12342 27004 12348 27056
rect 12400 27044 12406 27056
rect 14153 27047 14211 27053
rect 14153 27044 14165 27047
rect 12400 27016 14165 27044
rect 12400 27004 12406 27016
rect 14153 27013 14165 27016
rect 14199 27013 14211 27047
rect 14366 27044 14372 27056
rect 14327 27016 14372 27044
rect 14153 27007 14211 27013
rect 14366 27004 14372 27016
rect 14424 27004 14430 27056
rect 15562 27004 15568 27056
rect 15620 27044 15626 27056
rect 17972 27044 18000 27084
rect 21358 27072 21364 27084
rect 21416 27072 21422 27124
rect 22278 27112 22284 27124
rect 22066 27084 22284 27112
rect 15620 27016 17356 27044
rect 15620 27004 15626 27016
rect 12805 26979 12863 26985
rect 12805 26945 12817 26979
rect 12851 26976 12863 26979
rect 12986 26976 12992 26988
rect 12851 26948 12992 26976
rect 12851 26945 12863 26948
rect 12805 26939 12863 26945
rect 12986 26936 12992 26948
rect 13044 26936 13050 26988
rect 13449 26979 13507 26985
rect 13449 26945 13461 26979
rect 13495 26945 13507 26979
rect 13449 26939 13507 26945
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 8628 26880 13400 26908
rect 8628 26868 8634 26880
rect 13372 26784 13400 26880
rect 13464 26840 13492 26939
rect 13630 26936 13636 26988
rect 13688 26976 13694 26988
rect 13814 26976 13820 26988
rect 13688 26948 13820 26976
rect 13688 26936 13694 26948
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 14826 26976 14832 26988
rect 14787 26948 14832 26976
rect 14826 26936 14832 26948
rect 14884 26936 14890 26988
rect 14921 26979 14979 26985
rect 14921 26945 14933 26979
rect 14967 26945 14979 26979
rect 15286 26976 15292 26988
rect 15247 26948 15292 26976
rect 14921 26939 14979 26945
rect 13906 26868 13912 26920
rect 13964 26908 13970 26920
rect 14936 26908 14964 26939
rect 15286 26936 15292 26948
rect 15344 26936 15350 26988
rect 15856 26985 15884 27016
rect 17328 27010 17356 27016
rect 17504 27016 18000 27044
rect 17504 27010 17532 27016
rect 15841 26979 15899 26985
rect 15841 26945 15853 26979
rect 15887 26945 15899 26979
rect 15841 26939 15899 26945
rect 16114 26936 16120 26988
rect 16172 26976 16178 26988
rect 17328 26985 17532 27010
rect 18322 27004 18328 27056
rect 18380 27004 18386 27056
rect 18690 27004 18696 27056
rect 18748 27044 18754 27056
rect 19242 27044 19248 27056
rect 18748 27016 19248 27044
rect 18748 27004 18754 27016
rect 19242 27004 19248 27016
rect 19300 27004 19306 27056
rect 19610 27004 19616 27056
rect 19668 27044 19674 27056
rect 19668 27016 20484 27044
rect 19668 27004 19674 27016
rect 17300 26982 17532 26985
rect 17300 26979 17358 26982
rect 16172 26948 16217 26976
rect 16172 26936 16178 26948
rect 17300 26945 17312 26979
rect 17346 26945 17358 26979
rect 17300 26939 17358 26945
rect 17589 26979 17647 26985
rect 17589 26945 17601 26979
rect 17635 26976 17647 26979
rect 17678 26976 17684 26988
rect 17635 26948 17684 26976
rect 17635 26945 17647 26948
rect 17589 26939 17647 26945
rect 17678 26936 17684 26948
rect 17736 26936 17742 26988
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18340 26976 18368 27004
rect 20346 26985 20352 26988
rect 18279 26948 18368 26976
rect 18500 26980 18558 26985
rect 18500 26979 18644 26980
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18500 26945 18512 26979
rect 18546 26976 18644 26979
rect 20340 26976 20352 26985
rect 18546 26952 19288 26976
rect 18546 26945 18558 26952
rect 18616 26948 19288 26952
rect 20307 26948 20352 26976
rect 18500 26939 18558 26945
rect 19260 26920 19288 26948
rect 20340 26939 20352 26948
rect 20346 26936 20352 26939
rect 20404 26936 20410 26988
rect 20456 26976 20484 27016
rect 20530 27004 20536 27056
rect 20588 27044 20594 27056
rect 22066 27044 22094 27084
rect 22278 27072 22284 27084
rect 22336 27072 22342 27124
rect 23842 27112 23848 27124
rect 23803 27084 23848 27112
rect 23842 27072 23848 27084
rect 23900 27072 23906 27124
rect 24118 27072 24124 27124
rect 24176 27112 24182 27124
rect 25038 27112 25044 27124
rect 24176 27084 25044 27112
rect 24176 27072 24182 27084
rect 25038 27072 25044 27084
rect 25096 27072 25102 27124
rect 25130 27072 25136 27124
rect 25188 27112 25194 27124
rect 25685 27115 25743 27121
rect 25685 27112 25697 27115
rect 25188 27084 25697 27112
rect 25188 27072 25194 27084
rect 25685 27081 25697 27084
rect 25731 27081 25743 27115
rect 25685 27075 25743 27081
rect 25866 27072 25872 27124
rect 25924 27112 25930 27124
rect 25924 27084 27384 27112
rect 25924 27072 25930 27084
rect 27157 27047 27215 27053
rect 27157 27044 27169 27047
rect 20588 27016 22094 27044
rect 22132 27016 27169 27044
rect 20588 27004 20594 27016
rect 22132 26976 22160 27016
rect 27157 27013 27169 27016
rect 27203 27013 27215 27047
rect 27157 27007 27215 27013
rect 22278 26985 22284 26988
rect 22272 26976 22284 26985
rect 20456 26948 22160 26976
rect 22239 26948 22284 26976
rect 22272 26939 22284 26948
rect 22336 26976 22342 26988
rect 24578 26976 24584 26988
rect 22336 26948 24584 26976
rect 22278 26936 22284 26939
rect 22336 26936 22342 26948
rect 24578 26936 24584 26948
rect 24636 26936 24642 26988
rect 24969 26979 25027 26985
rect 24969 26945 24981 26979
rect 25015 26976 25027 26979
rect 25590 26976 25596 26988
rect 25015 26948 25596 26976
rect 25015 26945 25027 26948
rect 24969 26939 25027 26945
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 25866 26976 25872 26988
rect 25827 26948 25872 26976
rect 25866 26936 25872 26948
rect 25924 26936 25930 26988
rect 26145 26979 26203 26985
rect 26145 26945 26157 26979
rect 26191 26945 26203 26979
rect 26145 26939 26203 26945
rect 13964 26880 14964 26908
rect 15105 26911 15163 26917
rect 13964 26868 13970 26880
rect 15105 26877 15117 26911
rect 15151 26908 15163 26911
rect 16758 26908 16764 26920
rect 15151 26880 16764 26908
rect 15151 26877 15163 26880
rect 15105 26871 15163 26877
rect 16758 26868 16764 26880
rect 16816 26868 16822 26920
rect 17402 26868 17408 26920
rect 17460 26908 17466 26920
rect 17460 26880 17505 26908
rect 17460 26868 17466 26880
rect 19242 26868 19248 26920
rect 19300 26868 19306 26920
rect 19334 26868 19340 26920
rect 19392 26908 19398 26920
rect 19978 26908 19984 26920
rect 19392 26880 19984 26908
rect 19392 26868 19398 26880
rect 19978 26868 19984 26880
rect 20036 26908 20042 26920
rect 20073 26911 20131 26917
rect 20073 26908 20085 26911
rect 20036 26880 20085 26908
rect 20036 26868 20042 26880
rect 20073 26877 20085 26880
rect 20119 26877 20131 26911
rect 22002 26908 22008 26920
rect 21963 26880 22008 26908
rect 20073 26871 20131 26877
rect 22002 26868 22008 26880
rect 22060 26868 22066 26920
rect 25222 26908 25228 26920
rect 25183 26880 25228 26908
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 25682 26868 25688 26920
rect 25740 26908 25746 26920
rect 25961 26911 26019 26917
rect 25961 26908 25973 26911
rect 25740 26880 25973 26908
rect 25740 26868 25746 26880
rect 25961 26877 25973 26880
rect 26007 26877 26019 26911
rect 26160 26908 26188 26939
rect 26602 26936 26608 26988
rect 26660 26976 26666 26988
rect 27246 26976 27252 26988
rect 26660 26948 27252 26976
rect 26660 26936 26666 26948
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 27356 26985 27384 27084
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26976 27399 26979
rect 27522 26976 27528 26988
rect 27387 26948 27528 26976
rect 27387 26945 27399 26948
rect 27341 26939 27399 26945
rect 27522 26936 27528 26948
rect 27580 26936 27586 26988
rect 27614 26936 27620 26988
rect 27672 26976 27678 26988
rect 27672 26948 27717 26976
rect 27672 26936 27678 26948
rect 28074 26936 28080 26988
rect 28132 26976 28138 26988
rect 28353 26979 28411 26985
rect 28353 26976 28365 26979
rect 28132 26948 28365 26976
rect 28132 26936 28138 26948
rect 28353 26945 28365 26948
rect 28399 26945 28411 26979
rect 28353 26939 28411 26945
rect 26418 26908 26424 26920
rect 26160 26880 26424 26908
rect 25961 26871 26019 26877
rect 26418 26868 26424 26880
rect 26476 26908 26482 26920
rect 26476 26880 26648 26908
rect 26476 26868 26482 26880
rect 26620 26852 26648 26880
rect 27154 26868 27160 26920
rect 27212 26908 27218 26920
rect 27433 26911 27491 26917
rect 27433 26908 27445 26911
rect 27212 26880 27445 26908
rect 27212 26868 27218 26880
rect 27433 26877 27445 26880
rect 27479 26877 27491 26911
rect 27433 26871 27491 26877
rect 15746 26840 15752 26852
rect 13464 26812 15752 26840
rect 15746 26800 15752 26812
rect 15804 26800 15810 26852
rect 15933 26843 15991 26849
rect 15933 26809 15945 26843
rect 15979 26809 15991 26843
rect 15933 26803 15991 26809
rect 16025 26843 16083 26849
rect 16025 26809 16037 26843
rect 16071 26840 16083 26843
rect 16298 26840 16304 26852
rect 16071 26812 16304 26840
rect 16071 26809 16083 26812
rect 16025 26803 16083 26809
rect 8941 26775 8999 26781
rect 8941 26741 8953 26775
rect 8987 26772 8999 26775
rect 9766 26772 9772 26784
rect 8987 26744 9772 26772
rect 8987 26741 8999 26744
rect 8941 26735 8999 26741
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 13354 26772 13360 26784
rect 13315 26744 13360 26772
rect 13354 26732 13360 26744
rect 13412 26732 13418 26784
rect 14182 26772 14188 26784
rect 14143 26744 14188 26772
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 14550 26732 14556 26784
rect 14608 26772 14614 26784
rect 15562 26772 15568 26784
rect 14608 26744 15568 26772
rect 14608 26732 14614 26744
rect 15562 26732 15568 26744
rect 15620 26732 15626 26784
rect 15948 26772 15976 26803
rect 16298 26800 16304 26812
rect 16356 26800 16362 26852
rect 17497 26843 17555 26849
rect 17497 26809 17509 26843
rect 17543 26809 17555 26843
rect 21726 26840 21732 26852
rect 17497 26803 17555 26809
rect 21201 26812 21732 26840
rect 16114 26772 16120 26784
rect 15948 26744 16120 26772
rect 16114 26732 16120 26744
rect 16172 26732 16178 26784
rect 16758 26732 16764 26784
rect 16816 26772 16822 26784
rect 17512 26772 17540 26803
rect 16816 26744 17540 26772
rect 19613 26775 19671 26781
rect 16816 26732 16822 26744
rect 19613 26741 19625 26775
rect 19659 26772 19671 26775
rect 19794 26772 19800 26784
rect 19659 26744 19800 26772
rect 19659 26741 19671 26744
rect 19613 26735 19671 26741
rect 19794 26732 19800 26744
rect 19852 26732 19858 26784
rect 19978 26732 19984 26784
rect 20036 26772 20042 26784
rect 21201 26772 21229 26812
rect 21726 26800 21732 26812
rect 21784 26800 21790 26852
rect 23014 26800 23020 26852
rect 23072 26840 23078 26852
rect 23934 26840 23940 26852
rect 23072 26812 23940 26840
rect 23072 26800 23078 26812
rect 23934 26800 23940 26812
rect 23992 26800 23998 26852
rect 25498 26800 25504 26852
rect 25556 26840 25562 26852
rect 26053 26843 26111 26849
rect 26053 26840 26065 26843
rect 25556 26812 26065 26840
rect 25556 26800 25562 26812
rect 26053 26809 26065 26812
rect 26099 26809 26111 26843
rect 26053 26803 26111 26809
rect 26602 26800 26608 26852
rect 26660 26800 26666 26852
rect 27522 26840 27528 26852
rect 27483 26812 27528 26840
rect 27522 26800 27528 26812
rect 27580 26800 27586 26852
rect 20036 26744 21229 26772
rect 20036 26732 20042 26744
rect 21266 26732 21272 26784
rect 21324 26772 21330 26784
rect 21453 26775 21511 26781
rect 21453 26772 21465 26775
rect 21324 26744 21465 26772
rect 21324 26732 21330 26744
rect 21453 26741 21465 26744
rect 21499 26741 21511 26775
rect 21453 26735 21511 26741
rect 22278 26732 22284 26784
rect 22336 26772 22342 26784
rect 23385 26775 23443 26781
rect 23385 26772 23397 26775
rect 22336 26744 23397 26772
rect 22336 26732 22342 26744
rect 23385 26741 23397 26744
rect 23431 26772 23443 26775
rect 23658 26772 23664 26784
rect 23431 26744 23664 26772
rect 23431 26741 23443 26744
rect 23385 26735 23443 26741
rect 23658 26732 23664 26744
rect 23716 26732 23722 26784
rect 25038 26732 25044 26784
rect 25096 26772 25102 26784
rect 28169 26775 28227 26781
rect 28169 26772 28181 26775
rect 25096 26744 28181 26772
rect 25096 26732 25102 26744
rect 28169 26741 28181 26744
rect 28215 26741 28227 26775
rect 28169 26735 28227 26741
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 10413 26571 10471 26577
rect 10413 26537 10425 26571
rect 10459 26568 10471 26571
rect 10594 26568 10600 26580
rect 10459 26540 10600 26568
rect 10459 26537 10471 26540
rect 10413 26531 10471 26537
rect 10594 26528 10600 26540
rect 10652 26528 10658 26580
rect 10686 26528 10692 26580
rect 10744 26568 10750 26580
rect 11425 26571 11483 26577
rect 11425 26568 11437 26571
rect 10744 26540 11437 26568
rect 10744 26528 10750 26540
rect 11425 26537 11437 26540
rect 11471 26537 11483 26571
rect 12066 26568 12072 26580
rect 11979 26540 12072 26568
rect 11425 26531 11483 26537
rect 12066 26528 12072 26540
rect 12124 26568 12130 26580
rect 12342 26568 12348 26580
rect 12124 26540 12348 26568
rect 12124 26528 12130 26540
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 14182 26568 14188 26580
rect 12728 26540 14188 26568
rect 10965 26503 11023 26509
rect 10965 26469 10977 26503
rect 11011 26500 11023 26503
rect 11146 26500 11152 26512
rect 11011 26472 11152 26500
rect 11011 26469 11023 26472
rect 10965 26463 11023 26469
rect 11146 26460 11152 26472
rect 11204 26460 11210 26512
rect 12360 26500 12388 26528
rect 12360 26472 12480 26500
rect 11164 26432 11192 26460
rect 12342 26432 12348 26444
rect 11164 26404 12348 26432
rect 12342 26392 12348 26404
rect 12400 26392 12406 26444
rect 1578 26364 1584 26376
rect 1539 26336 1584 26364
rect 1578 26324 1584 26336
rect 1636 26324 1642 26376
rect 9858 26364 9864 26376
rect 9819 26336 9864 26364
rect 9858 26324 9864 26336
rect 9916 26324 9922 26376
rect 12452 26364 12480 26472
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 12728 26432 12756 26540
rect 14182 26528 14188 26540
rect 14240 26568 14246 26580
rect 14829 26571 14887 26577
rect 14829 26568 14841 26571
rect 14240 26540 14841 26568
rect 14240 26528 14246 26540
rect 14829 26537 14841 26540
rect 14875 26537 14887 26571
rect 16025 26571 16083 26577
rect 14829 26531 14887 26537
rect 15498 26540 15976 26568
rect 14366 26460 14372 26512
rect 14424 26500 14430 26512
rect 14642 26500 14648 26512
rect 14424 26472 14648 26500
rect 14424 26460 14430 26472
rect 14642 26460 14648 26472
rect 14700 26460 14706 26512
rect 15013 26503 15071 26509
rect 15013 26469 15025 26503
rect 15059 26500 15071 26503
rect 15498 26500 15526 26540
rect 15059 26472 15526 26500
rect 15059 26469 15071 26472
rect 15013 26463 15071 26469
rect 15654 26460 15660 26512
rect 15712 26500 15718 26512
rect 15712 26472 15792 26500
rect 15712 26460 15718 26472
rect 12676 26404 12756 26432
rect 12676 26392 12682 26404
rect 13354 26392 13360 26444
rect 13412 26432 13418 26444
rect 13412 26404 15056 26432
rect 13412 26392 13418 26404
rect 13081 26367 13139 26373
rect 13081 26364 13093 26367
rect 12452 26336 13093 26364
rect 13081 26333 13093 26336
rect 13127 26364 13139 26367
rect 13127 26336 14888 26364
rect 13127 26333 13139 26336
rect 13081 26327 13139 26333
rect 11882 26256 11888 26308
rect 11940 26296 11946 26308
rect 13906 26296 13912 26308
rect 11940 26268 13912 26296
rect 11940 26256 11946 26268
rect 13906 26256 13912 26268
rect 13964 26256 13970 26308
rect 14642 26296 14648 26308
rect 14603 26268 14648 26296
rect 14642 26256 14648 26268
rect 14700 26256 14706 26308
rect 14860 26305 14888 26336
rect 14845 26299 14903 26305
rect 14845 26265 14857 26299
rect 14891 26265 14903 26299
rect 15028 26296 15056 26404
rect 15102 26324 15108 26376
rect 15160 26364 15166 26376
rect 15463 26367 15521 26373
rect 15463 26364 15475 26367
rect 15160 26336 15475 26364
rect 15160 26324 15166 26336
rect 15463 26333 15475 26336
rect 15509 26333 15521 26367
rect 15463 26327 15521 26333
rect 15562 26324 15568 26376
rect 15620 26364 15626 26376
rect 15764 26373 15792 26472
rect 15948 26432 15976 26540
rect 16025 26537 16037 26571
rect 16071 26568 16083 26571
rect 23382 26568 23388 26580
rect 16071 26540 23388 26568
rect 16071 26537 16083 26540
rect 16025 26531 16083 26537
rect 23382 26528 23388 26540
rect 23440 26528 23446 26580
rect 27801 26571 27859 26577
rect 27801 26568 27813 26571
rect 23492 26540 27813 26568
rect 16114 26460 16120 26512
rect 16172 26500 16178 26512
rect 16482 26500 16488 26512
rect 16172 26472 16488 26500
rect 16172 26460 16178 26472
rect 16482 26460 16488 26472
rect 16540 26460 16546 26512
rect 16574 26460 16580 26512
rect 16632 26460 16638 26512
rect 17037 26503 17095 26509
rect 17037 26469 17049 26503
rect 17083 26500 17095 26503
rect 17126 26500 17132 26512
rect 17083 26472 17132 26500
rect 17083 26469 17095 26472
rect 17037 26463 17095 26469
rect 17126 26460 17132 26472
rect 17184 26460 17190 26512
rect 18690 26460 18696 26512
rect 18748 26500 18754 26512
rect 18877 26503 18935 26509
rect 18877 26500 18889 26503
rect 18748 26472 18889 26500
rect 18748 26460 18754 26472
rect 18877 26469 18889 26472
rect 18923 26469 18935 26503
rect 18877 26463 18935 26469
rect 20806 26460 20812 26512
rect 20864 26500 20870 26512
rect 20901 26503 20959 26509
rect 20901 26500 20913 26503
rect 20864 26472 20913 26500
rect 20864 26460 20870 26472
rect 20901 26469 20913 26472
rect 20947 26500 20959 26503
rect 20990 26500 20996 26512
rect 20947 26472 20996 26500
rect 20947 26469 20959 26472
rect 20901 26463 20959 26469
rect 20990 26460 20996 26472
rect 21048 26460 21054 26512
rect 23198 26500 23204 26512
rect 23159 26472 23204 26500
rect 23198 26460 23204 26472
rect 23256 26460 23262 26512
rect 16592 26432 16620 26460
rect 17494 26432 17500 26444
rect 15948 26404 16528 26432
rect 16592 26404 16896 26432
rect 17455 26404 17500 26432
rect 15749 26367 15807 26373
rect 15620 26336 15665 26364
rect 15620 26324 15626 26336
rect 15749 26333 15761 26367
rect 15795 26333 15807 26367
rect 15749 26327 15807 26333
rect 15841 26367 15899 26373
rect 15841 26333 15853 26367
rect 15887 26364 15899 26367
rect 16114 26364 16120 26376
rect 15887 26336 16120 26364
rect 15887 26333 15899 26336
rect 15841 26327 15899 26333
rect 16114 26324 16120 26336
rect 16172 26324 16178 26376
rect 16500 26373 16528 26404
rect 16485 26367 16543 26373
rect 16485 26333 16497 26367
rect 16531 26333 16543 26367
rect 16485 26327 16543 26333
rect 16577 26367 16635 26373
rect 16577 26333 16589 26367
rect 16623 26364 16635 26367
rect 16666 26364 16672 26376
rect 16623 26336 16672 26364
rect 16623 26333 16635 26336
rect 16577 26327 16635 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 16868 26373 16896 26404
rect 17494 26392 17500 26404
rect 17552 26392 17558 26444
rect 18506 26392 18512 26444
rect 18564 26432 18570 26444
rect 19518 26432 19524 26444
rect 18564 26404 19524 26432
rect 18564 26392 18570 26404
rect 19518 26392 19524 26404
rect 19576 26392 19582 26444
rect 23492 26432 23520 26540
rect 27801 26537 27813 26540
rect 27847 26537 27859 26571
rect 28350 26568 28356 26580
rect 28311 26540 28356 26568
rect 27801 26531 27859 26537
rect 28350 26528 28356 26540
rect 28408 26528 28414 26580
rect 23750 26500 23756 26512
rect 22664 26404 23520 26432
rect 23584 26472 23756 26500
rect 19794 26373 19800 26376
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26333 16819 26367
rect 16761 26327 16819 26333
rect 16853 26367 16911 26373
rect 16853 26333 16865 26367
rect 16899 26333 16911 26367
rect 19788 26364 19800 26373
rect 17650 26358 19682 26364
rect 16853 26327 16911 26333
rect 17604 26336 19682 26358
rect 19755 26336 19800 26364
rect 17604 26330 17678 26336
rect 16776 26296 16804 26327
rect 17604 26296 17632 26330
rect 17770 26305 17776 26308
rect 15028 26268 16712 26296
rect 16776 26268 17632 26296
rect 14845 26259 14903 26265
rect 13725 26231 13783 26237
rect 13725 26197 13737 26231
rect 13771 26228 13783 26231
rect 16298 26228 16304 26240
rect 13771 26200 16304 26228
rect 13771 26197 13783 26200
rect 13725 26191 13783 26197
rect 16298 26188 16304 26200
rect 16356 26188 16362 26240
rect 16684 26228 16712 26268
rect 17764 26259 17776 26305
rect 17828 26296 17834 26308
rect 19334 26296 19340 26308
rect 17828 26268 17864 26296
rect 18524 26268 19340 26296
rect 17770 26256 17776 26259
rect 17828 26256 17834 26268
rect 18524 26228 18552 26268
rect 19334 26256 19340 26268
rect 19392 26256 19398 26308
rect 19654 26296 19682 26336
rect 19788 26327 19800 26336
rect 19794 26324 19800 26327
rect 19852 26324 19858 26376
rect 21082 26364 21088 26376
rect 20640 26336 21088 26364
rect 20640 26296 20668 26336
rect 21082 26324 21088 26336
rect 21140 26324 21146 26376
rect 21174 26324 21180 26376
rect 21232 26364 21238 26376
rect 22664 26364 22692 26404
rect 21232 26336 22692 26364
rect 22741 26367 22799 26373
rect 21232 26324 21238 26336
rect 22741 26333 22753 26367
rect 22787 26364 22799 26367
rect 23014 26364 23020 26376
rect 22787 26336 23020 26364
rect 22787 26333 22799 26336
rect 22741 26327 22799 26333
rect 19654 26268 20668 26296
rect 20714 26256 20720 26308
rect 20772 26296 20778 26308
rect 22094 26296 22100 26308
rect 20772 26268 22100 26296
rect 20772 26256 20778 26268
rect 22094 26256 22100 26268
rect 22152 26296 22158 26308
rect 22496 26299 22554 26305
rect 22496 26296 22508 26299
rect 22152 26268 22508 26296
rect 22152 26256 22158 26268
rect 22496 26265 22508 26268
rect 22542 26265 22554 26299
rect 22496 26259 22554 26265
rect 16684 26200 18552 26228
rect 18598 26188 18604 26240
rect 18656 26228 18662 26240
rect 18966 26228 18972 26240
rect 18656 26200 18972 26228
rect 18656 26188 18662 26200
rect 18966 26188 18972 26200
rect 19024 26188 19030 26240
rect 20162 26188 20168 26240
rect 20220 26228 20226 26240
rect 21361 26231 21419 26237
rect 21361 26228 21373 26231
rect 20220 26200 21373 26228
rect 20220 26188 20226 26200
rect 21361 26197 21373 26200
rect 21407 26197 21419 26231
rect 21361 26191 21419 26197
rect 22186 26188 22192 26240
rect 22244 26228 22250 26240
rect 22756 26228 22784 26327
rect 23014 26324 23020 26336
rect 23072 26324 23078 26376
rect 23382 26364 23388 26376
rect 23343 26336 23388 26364
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26364 23535 26367
rect 23584 26364 23612 26472
rect 23750 26460 23756 26472
rect 23808 26460 23814 26512
rect 24578 26500 24584 26512
rect 24539 26472 24584 26500
rect 24578 26460 24584 26472
rect 24636 26460 24642 26512
rect 26050 26392 26056 26444
rect 26108 26432 26114 26444
rect 26108 26404 26188 26432
rect 26108 26392 26114 26404
rect 23842 26364 23848 26376
rect 23523 26336 23612 26364
rect 23803 26336 23848 26364
rect 23523 26333 23535 26336
rect 23477 26327 23535 26333
rect 23842 26324 23848 26336
rect 23900 26324 23906 26376
rect 24394 26324 24400 26376
rect 24452 26364 24458 26376
rect 25961 26367 26019 26373
rect 25961 26364 25973 26367
rect 24452 26336 25973 26364
rect 24452 26324 24458 26336
rect 25961 26333 25973 26336
rect 26007 26333 26019 26367
rect 26160 26364 26188 26404
rect 26421 26367 26479 26373
rect 26421 26364 26433 26367
rect 26160 26336 26433 26364
rect 25961 26327 26019 26333
rect 26421 26333 26433 26336
rect 26467 26333 26479 26367
rect 26421 26327 26479 26333
rect 23569 26299 23627 26305
rect 23569 26296 23581 26299
rect 23124 26268 23581 26296
rect 23124 26240 23152 26268
rect 23569 26265 23581 26268
rect 23615 26265 23627 26299
rect 23569 26259 23627 26265
rect 23658 26256 23664 26308
rect 23716 26305 23722 26308
rect 23716 26299 23745 26305
rect 23733 26265 23745 26299
rect 25590 26296 25596 26308
rect 23716 26259 23745 26265
rect 23860 26268 25596 26296
rect 23716 26256 23722 26259
rect 22244 26200 22784 26228
rect 22244 26188 22250 26200
rect 23106 26188 23112 26240
rect 23164 26188 23170 26240
rect 23290 26188 23296 26240
rect 23348 26228 23354 26240
rect 23860 26228 23888 26268
rect 25590 26256 25596 26268
rect 25648 26256 25654 26308
rect 25716 26299 25774 26305
rect 25716 26265 25728 26299
rect 25762 26296 25774 26299
rect 26050 26296 26056 26308
rect 25762 26268 26056 26296
rect 25762 26265 25774 26268
rect 25716 26259 25774 26265
rect 26050 26256 26056 26268
rect 26108 26256 26114 26308
rect 26142 26256 26148 26308
rect 26200 26296 26206 26308
rect 26666 26299 26724 26305
rect 26666 26296 26678 26299
rect 26200 26268 26678 26296
rect 26200 26256 26206 26268
rect 26666 26265 26678 26268
rect 26712 26296 26724 26299
rect 27154 26296 27160 26308
rect 26712 26268 27160 26296
rect 26712 26265 26724 26268
rect 26666 26259 26724 26265
rect 27154 26256 27160 26268
rect 27212 26256 27218 26308
rect 23348 26200 23888 26228
rect 23348 26188 23354 26200
rect 23934 26188 23940 26240
rect 23992 26228 23998 26240
rect 24854 26228 24860 26240
rect 23992 26200 24860 26228
rect 23992 26188 23998 26200
rect 24854 26188 24860 26200
rect 24912 26188 24918 26240
rect 25038 26188 25044 26240
rect 25096 26228 25102 26240
rect 26234 26228 26240 26240
rect 25096 26200 26240 26228
rect 25096 26188 25102 26200
rect 26234 26188 26240 26200
rect 26292 26188 26298 26240
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 9674 25984 9680 26036
rect 9732 26024 9738 26036
rect 10410 26024 10416 26036
rect 9732 25996 10416 26024
rect 9732 25984 9738 25996
rect 10410 25984 10416 25996
rect 10468 25984 10474 26036
rect 12158 25984 12164 26036
rect 12216 26024 12222 26036
rect 12989 26027 13047 26033
rect 12989 26024 13001 26027
rect 12216 25996 13001 26024
rect 12216 25984 12222 25996
rect 12989 25993 13001 25996
rect 13035 26024 13047 26027
rect 14734 26024 14740 26036
rect 13035 25996 14740 26024
rect 13035 25993 13047 25996
rect 12989 25987 13047 25993
rect 14734 25984 14740 25996
rect 14792 25984 14798 26036
rect 15194 25984 15200 26036
rect 15252 26024 15258 26036
rect 15933 26027 15991 26033
rect 15933 26024 15945 26027
rect 15252 25996 15945 26024
rect 15252 25984 15258 25996
rect 15933 25993 15945 25996
rect 15979 25993 15991 26027
rect 15933 25987 15991 25993
rect 16666 25984 16672 26036
rect 16724 26024 16730 26036
rect 16724 25996 17724 26024
rect 16724 25984 16730 25996
rect 13538 25916 13544 25968
rect 13596 25956 13602 25968
rect 15473 25959 15531 25965
rect 13596 25928 15424 25956
rect 13596 25916 13602 25928
rect 10594 25848 10600 25900
rect 10652 25888 10658 25900
rect 14642 25888 14648 25900
rect 10652 25860 14648 25888
rect 10652 25848 10658 25860
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 14734 25848 14740 25900
rect 14792 25888 14798 25900
rect 15289 25891 15347 25897
rect 15289 25888 15301 25891
rect 14792 25860 15301 25888
rect 14792 25848 14798 25860
rect 15289 25857 15301 25860
rect 15335 25857 15347 25891
rect 15396 25888 15424 25928
rect 15473 25925 15485 25959
rect 15519 25956 15531 25959
rect 15838 25956 15844 25968
rect 15519 25928 15844 25956
rect 15519 25925 15531 25928
rect 15473 25919 15531 25925
rect 15838 25916 15844 25928
rect 15896 25916 15902 25968
rect 16101 25959 16159 25965
rect 16101 25956 16113 25959
rect 15948 25928 16113 25956
rect 15948 25888 15976 25928
rect 16101 25925 16113 25928
rect 16147 25956 16159 25959
rect 16206 25956 16212 25968
rect 16147 25928 16212 25956
rect 16147 25925 16159 25928
rect 16101 25919 16159 25925
rect 16206 25916 16212 25928
rect 16264 25916 16270 25968
rect 16301 25959 16359 25965
rect 16301 25925 16313 25959
rect 16347 25925 16359 25959
rect 16301 25919 16359 25925
rect 15396 25860 15976 25888
rect 15289 25851 15347 25857
rect 15304 25820 15332 25851
rect 15654 25820 15660 25832
rect 15304 25792 15660 25820
rect 15654 25780 15660 25792
rect 15712 25780 15718 25832
rect 16022 25780 16028 25832
rect 16080 25820 16086 25832
rect 16316 25820 16344 25919
rect 16758 25916 16764 25968
rect 16816 25956 16822 25968
rect 17221 25959 17279 25965
rect 17221 25956 17233 25959
rect 16816 25928 17233 25956
rect 16816 25916 16822 25928
rect 17221 25925 17233 25928
rect 17267 25925 17279 25959
rect 17221 25919 17279 25925
rect 17696 25956 17724 25996
rect 17770 25984 17776 26036
rect 17828 26024 17834 26036
rect 19610 26024 19616 26036
rect 17828 25996 19616 26024
rect 17828 25984 17834 25996
rect 19610 25984 19616 25996
rect 19668 25984 19674 26036
rect 19702 25984 19708 26036
rect 19760 26024 19766 26036
rect 19760 25996 21312 26024
rect 19760 25984 19766 25996
rect 18500 25959 18558 25965
rect 17696 25928 18460 25956
rect 17405 25891 17463 25897
rect 17405 25888 17417 25891
rect 17328 25860 17417 25888
rect 16080 25792 16344 25820
rect 16080 25780 16086 25792
rect 17218 25780 17224 25832
rect 17276 25820 17282 25832
rect 17328 25820 17356 25860
rect 17405 25857 17417 25860
rect 17451 25857 17463 25891
rect 17405 25851 17463 25857
rect 17494 25848 17500 25900
rect 17552 25888 17558 25900
rect 17696 25897 17724 25928
rect 17681 25891 17739 25897
rect 17552 25860 17597 25888
rect 17552 25848 17558 25860
rect 17681 25857 17693 25891
rect 17727 25857 17739 25891
rect 17681 25851 17739 25857
rect 17770 25848 17776 25900
rect 17828 25888 17834 25900
rect 18233 25891 18291 25897
rect 17828 25860 17873 25888
rect 17828 25848 17834 25860
rect 18233 25857 18245 25891
rect 18279 25888 18291 25891
rect 18322 25888 18328 25900
rect 18279 25860 18328 25888
rect 18279 25857 18291 25860
rect 18233 25851 18291 25857
rect 18322 25848 18328 25860
rect 18380 25848 18386 25900
rect 18432 25888 18460 25928
rect 18500 25925 18512 25959
rect 18546 25956 18558 25959
rect 19150 25956 19156 25968
rect 18546 25928 19156 25956
rect 18546 25925 18558 25928
rect 18500 25919 18558 25925
rect 19150 25916 19156 25928
rect 19208 25916 19214 25968
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 21186 25959 21244 25965
rect 21186 25956 21198 25959
rect 19392 25928 21198 25956
rect 19392 25916 19398 25928
rect 21186 25925 21198 25928
rect 21232 25925 21244 25959
rect 21284 25956 21312 25996
rect 21358 25984 21364 26036
rect 21416 26024 21422 26036
rect 23658 26024 23664 26036
rect 21416 25996 23664 26024
rect 21416 25984 21422 25996
rect 23658 25984 23664 25996
rect 23716 25984 23722 26036
rect 23842 25984 23848 26036
rect 23900 26024 23906 26036
rect 25685 26027 25743 26033
rect 25685 26024 25697 26027
rect 23900 25996 25697 26024
rect 23900 25984 23906 25996
rect 25685 25993 25697 25996
rect 25731 25993 25743 26027
rect 25685 25987 25743 25993
rect 26050 25984 26056 26036
rect 26108 26024 26114 26036
rect 26108 25996 27936 26024
rect 26108 25984 26114 25996
rect 24958 25959 25016 25965
rect 24958 25956 24970 25959
rect 21284 25928 24970 25956
rect 21186 25919 21244 25925
rect 24958 25925 24970 25928
rect 25004 25925 25016 25959
rect 26602 25956 26608 25968
rect 24958 25919 25016 25925
rect 25056 25928 26608 25956
rect 18966 25888 18972 25900
rect 18432 25860 18972 25888
rect 18966 25848 18972 25860
rect 19024 25848 19030 25900
rect 20162 25848 20168 25900
rect 20220 25888 20226 25900
rect 20346 25888 20352 25900
rect 20220 25860 20352 25888
rect 20220 25848 20226 25860
rect 20346 25848 20352 25860
rect 20404 25848 20410 25900
rect 20806 25848 20812 25900
rect 20864 25888 20870 25900
rect 21453 25891 21511 25897
rect 21453 25888 21465 25891
rect 20864 25860 21465 25888
rect 20864 25848 20870 25860
rect 21453 25857 21465 25860
rect 21499 25857 21511 25891
rect 21453 25851 21511 25857
rect 19978 25820 19984 25832
rect 17276 25792 17356 25820
rect 19536 25792 19984 25820
rect 17276 25780 17282 25792
rect 11149 25755 11207 25761
rect 11149 25721 11161 25755
rect 11195 25752 11207 25755
rect 12342 25752 12348 25764
rect 11195 25724 12348 25752
rect 11195 25721 11207 25724
rect 11149 25715 11207 25721
rect 12342 25712 12348 25724
rect 12400 25712 12406 25764
rect 14182 25752 14188 25764
rect 14143 25724 14188 25752
rect 14182 25712 14188 25724
rect 14240 25752 14246 25764
rect 14550 25752 14556 25764
rect 14240 25724 14556 25752
rect 14240 25712 14246 25724
rect 14550 25712 14556 25724
rect 14608 25712 14614 25764
rect 14642 25712 14648 25764
rect 14700 25752 14706 25764
rect 14700 25724 16160 25752
rect 14700 25712 14706 25724
rect 1578 25684 1584 25696
rect 1539 25656 1584 25684
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 11974 25684 11980 25696
rect 11935 25656 11980 25684
rect 11974 25644 11980 25656
rect 12032 25644 12038 25696
rect 12526 25684 12532 25696
rect 12487 25656 12532 25684
rect 12526 25644 12532 25656
rect 12584 25644 12590 25696
rect 13541 25687 13599 25693
rect 13541 25653 13553 25687
rect 13587 25684 13599 25687
rect 16022 25684 16028 25696
rect 13587 25656 16028 25684
rect 13587 25653 13599 25656
rect 13541 25647 13599 25653
rect 16022 25644 16028 25656
rect 16080 25644 16086 25696
rect 16132 25693 16160 25724
rect 16482 25712 16488 25764
rect 16540 25752 16546 25764
rect 17586 25752 17592 25764
rect 16540 25724 17592 25752
rect 16540 25712 16546 25724
rect 17586 25712 17592 25724
rect 17644 25712 17650 25764
rect 16117 25687 16175 25693
rect 16117 25653 16129 25687
rect 16163 25684 16175 25687
rect 16666 25684 16672 25696
rect 16163 25656 16672 25684
rect 16163 25653 16175 25656
rect 16117 25647 16175 25653
rect 16666 25644 16672 25656
rect 16724 25644 16730 25696
rect 17494 25644 17500 25696
rect 17552 25684 17558 25696
rect 19536 25684 19564 25792
rect 19978 25780 19984 25792
rect 20036 25780 20042 25832
rect 21468 25820 21496 25851
rect 21726 25848 21732 25900
rect 21784 25888 21790 25900
rect 22261 25891 22319 25897
rect 22261 25888 22273 25891
rect 21784 25860 22273 25888
rect 21784 25848 21790 25860
rect 22261 25857 22273 25860
rect 22307 25857 22319 25891
rect 22261 25851 22319 25857
rect 23658 25848 23664 25900
rect 23716 25888 23722 25900
rect 25056 25888 25084 25928
rect 25222 25888 25228 25900
rect 23716 25860 25084 25888
rect 25183 25860 25228 25888
rect 23716 25848 23722 25860
rect 25222 25848 25228 25860
rect 25280 25848 25286 25900
rect 25866 25888 25872 25900
rect 25827 25860 25872 25888
rect 25866 25848 25872 25860
rect 25924 25848 25930 25900
rect 26160 25897 26188 25928
rect 26602 25916 26608 25928
rect 26660 25916 26666 25968
rect 27154 25916 27160 25968
rect 27212 25956 27218 25968
rect 27908 25956 27936 25996
rect 27982 25984 27988 26036
rect 28040 26024 28046 26036
rect 28261 26027 28319 26033
rect 28261 26024 28273 26027
rect 28040 25996 28273 26024
rect 28040 25984 28046 25996
rect 28261 25993 28273 25996
rect 28307 25993 28319 26027
rect 28261 25987 28319 25993
rect 29454 25956 29460 25968
rect 27212 25928 27476 25956
rect 27908 25928 29460 25956
rect 27212 25916 27218 25928
rect 26145 25891 26203 25897
rect 26145 25857 26157 25891
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26878 25848 26884 25900
rect 26936 25888 26942 25900
rect 27448 25897 27476 25928
rect 29454 25916 29460 25928
rect 29512 25916 29518 25968
rect 27341 25891 27399 25897
rect 27341 25888 27353 25891
rect 26936 25860 27353 25888
rect 26936 25848 26942 25860
rect 27341 25857 27353 25860
rect 27387 25857 27399 25891
rect 27341 25851 27399 25857
rect 27433 25891 27491 25897
rect 27433 25857 27445 25891
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 27522 25848 27528 25900
rect 27580 25888 27586 25900
rect 27617 25891 27675 25897
rect 27617 25888 27629 25891
rect 27580 25860 27629 25888
rect 27580 25848 27586 25860
rect 27617 25857 27629 25860
rect 27663 25857 27675 25891
rect 27617 25851 27675 25857
rect 27709 25891 27767 25897
rect 27709 25857 27721 25891
rect 27755 25857 27767 25891
rect 27709 25851 27767 25857
rect 22002 25820 22008 25832
rect 21468 25792 22008 25820
rect 22002 25780 22008 25792
rect 22060 25780 22066 25832
rect 24118 25820 24124 25832
rect 23032 25792 24124 25820
rect 19613 25755 19671 25761
rect 19613 25721 19625 25755
rect 19659 25752 19671 25755
rect 20346 25752 20352 25764
rect 19659 25724 20352 25752
rect 19659 25721 19671 25724
rect 19613 25715 19671 25721
rect 20346 25712 20352 25724
rect 20404 25712 20410 25764
rect 20070 25684 20076 25696
rect 17552 25656 19564 25684
rect 20031 25656 20076 25684
rect 17552 25644 17558 25656
rect 20070 25644 20076 25656
rect 20128 25644 20134 25696
rect 20806 25644 20812 25696
rect 20864 25684 20870 25696
rect 21726 25684 21732 25696
rect 20864 25656 21732 25684
rect 20864 25644 20870 25656
rect 21726 25644 21732 25656
rect 21784 25644 21790 25696
rect 21818 25644 21824 25696
rect 21876 25684 21882 25696
rect 23032 25684 23060 25792
rect 24118 25780 24124 25792
rect 24176 25780 24182 25832
rect 26053 25823 26111 25829
rect 26053 25820 26065 25823
rect 25424 25792 26065 25820
rect 23106 25712 23112 25764
rect 23164 25752 23170 25764
rect 23845 25755 23903 25761
rect 23845 25752 23857 25755
rect 23164 25724 23857 25752
rect 23164 25712 23170 25724
rect 23845 25721 23857 25724
rect 23891 25721 23903 25755
rect 23845 25715 23903 25721
rect 23382 25684 23388 25696
rect 21876 25656 23060 25684
rect 23343 25656 23388 25684
rect 21876 25644 21882 25656
rect 23382 25644 23388 25656
rect 23440 25644 23446 25696
rect 23934 25644 23940 25696
rect 23992 25684 23998 25696
rect 25424 25684 25452 25792
rect 26053 25789 26065 25792
rect 26099 25789 26111 25823
rect 26053 25783 26111 25789
rect 26786 25780 26792 25832
rect 26844 25820 26850 25832
rect 27724 25820 27752 25851
rect 27798 25848 27804 25900
rect 27856 25888 27862 25900
rect 28169 25891 28227 25897
rect 28169 25888 28181 25891
rect 27856 25860 28181 25888
rect 27856 25848 27862 25860
rect 28169 25857 28181 25860
rect 28215 25857 28227 25891
rect 28350 25888 28356 25900
rect 28311 25860 28356 25888
rect 28169 25851 28227 25857
rect 28350 25848 28356 25860
rect 28408 25848 28414 25900
rect 26844 25792 27752 25820
rect 26844 25780 26850 25792
rect 25774 25712 25780 25764
rect 25832 25752 25838 25764
rect 25961 25755 26019 25761
rect 25961 25752 25973 25755
rect 25832 25724 25973 25752
rect 25832 25712 25838 25724
rect 25961 25721 25973 25724
rect 26007 25721 26019 25755
rect 27154 25752 27160 25764
rect 27115 25724 27160 25752
rect 25961 25715 26019 25721
rect 27154 25712 27160 25724
rect 27212 25712 27218 25764
rect 23992 25656 25452 25684
rect 23992 25644 23998 25656
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 12066 25480 12072 25492
rect 12027 25452 12072 25480
rect 12066 25440 12072 25452
rect 12124 25440 12130 25492
rect 12802 25440 12808 25492
rect 12860 25480 12866 25492
rect 13081 25483 13139 25489
rect 13081 25480 13093 25483
rect 12860 25452 13093 25480
rect 12860 25440 12866 25452
rect 13081 25449 13093 25452
rect 13127 25480 13139 25483
rect 13538 25480 13544 25492
rect 13127 25452 13544 25480
rect 13127 25449 13139 25452
rect 13081 25443 13139 25449
rect 13538 25440 13544 25452
rect 13596 25440 13602 25492
rect 13722 25440 13728 25492
rect 13780 25480 13786 25492
rect 16485 25483 16543 25489
rect 16485 25480 16497 25483
rect 13780 25452 16497 25480
rect 13780 25440 13786 25452
rect 16485 25449 16497 25452
rect 16531 25449 16543 25483
rect 16666 25480 16672 25492
rect 16627 25452 16672 25480
rect 16485 25443 16543 25449
rect 16666 25440 16672 25452
rect 16724 25440 16730 25492
rect 17630 25452 18276 25480
rect 11974 25372 11980 25424
rect 12032 25412 12038 25424
rect 14366 25412 14372 25424
rect 12032 25384 14372 25412
rect 12032 25372 12038 25384
rect 14366 25372 14372 25384
rect 14424 25412 14430 25424
rect 14734 25412 14740 25424
rect 14424 25384 14740 25412
rect 14424 25372 14430 25384
rect 14734 25372 14740 25384
rect 14792 25372 14798 25424
rect 15746 25412 15752 25424
rect 15707 25384 15752 25412
rect 15746 25372 15752 25384
rect 15804 25372 15810 25424
rect 17218 25372 17224 25424
rect 17276 25412 17282 25424
rect 17313 25415 17371 25421
rect 17313 25412 17325 25415
rect 17276 25384 17325 25412
rect 17276 25372 17282 25384
rect 17313 25381 17325 25384
rect 17359 25381 17371 25415
rect 17313 25375 17371 25381
rect 13446 25304 13452 25356
rect 13504 25344 13510 25356
rect 17630 25344 17658 25452
rect 13504 25316 17658 25344
rect 18248 25344 18276 25452
rect 18322 25440 18328 25492
rect 18380 25480 18386 25492
rect 18380 25452 18425 25480
rect 18380 25440 18386 25452
rect 19242 25440 19248 25492
rect 19300 25480 19306 25492
rect 19429 25483 19487 25489
rect 19429 25480 19441 25483
rect 19300 25452 19441 25480
rect 19300 25440 19306 25452
rect 19429 25449 19441 25452
rect 19475 25449 19487 25483
rect 20162 25480 20168 25492
rect 19429 25443 19487 25449
rect 19536 25452 20168 25480
rect 18690 25372 18696 25424
rect 18748 25412 18754 25424
rect 18966 25412 18972 25424
rect 18748 25384 18972 25412
rect 18748 25372 18754 25384
rect 18966 25372 18972 25384
rect 19024 25372 19030 25424
rect 19058 25372 19064 25424
rect 19116 25412 19122 25424
rect 19536 25412 19564 25452
rect 20162 25440 20168 25452
rect 20220 25440 20226 25492
rect 21082 25440 21088 25492
rect 21140 25480 21146 25492
rect 22738 25480 22744 25492
rect 21140 25452 22744 25480
rect 21140 25440 21146 25452
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 23106 25440 23112 25492
rect 23164 25480 23170 25492
rect 23164 25452 23520 25480
rect 23164 25440 23170 25452
rect 23492 25421 23520 25452
rect 23750 25440 23756 25492
rect 23808 25480 23814 25492
rect 24854 25480 24860 25492
rect 23808 25452 24860 25480
rect 23808 25440 23814 25452
rect 24854 25440 24860 25452
rect 24912 25440 24918 25492
rect 26970 25480 26976 25492
rect 24964 25452 26004 25480
rect 26931 25452 26976 25480
rect 19116 25384 19564 25412
rect 23477 25415 23535 25421
rect 19116 25372 19122 25384
rect 23477 25381 23489 25415
rect 23523 25381 23535 25415
rect 23477 25375 23535 25381
rect 19794 25344 19800 25356
rect 18248 25316 19800 25344
rect 13504 25304 13510 25316
rect 10778 25236 10784 25288
rect 10836 25276 10842 25288
rect 17218 25276 17224 25288
rect 10836 25248 17224 25276
rect 10836 25236 10842 25248
rect 17218 25236 17224 25248
rect 17276 25236 17282 25288
rect 17310 25236 17316 25288
rect 17368 25276 17374 25288
rect 17630 25285 17658 25316
rect 19794 25304 19800 25316
rect 19852 25304 19858 25356
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 24964 25344 24992 25452
rect 25976 25412 26004 25452
rect 26970 25440 26976 25452
rect 27028 25440 27034 25492
rect 28350 25412 28356 25424
rect 25976 25384 28356 25412
rect 28350 25372 28356 25384
rect 28408 25372 28414 25424
rect 24912 25316 24992 25344
rect 24912 25304 24918 25316
rect 26234 25304 26240 25356
rect 26292 25344 26298 25356
rect 27338 25344 27344 25356
rect 26292 25316 27344 25344
rect 26292 25304 26298 25316
rect 17497 25279 17555 25285
rect 17368 25270 17448 25276
rect 17497 25270 17509 25279
rect 17368 25248 17509 25270
rect 17368 25236 17374 25248
rect 17420 25245 17509 25248
rect 17543 25245 17555 25279
rect 17420 25242 17555 25245
rect 17497 25239 17555 25242
rect 17589 25279 17658 25285
rect 17589 25245 17601 25279
rect 17635 25245 17658 25279
rect 17589 25242 17658 25245
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25245 17831 25279
rect 17589 25239 17647 25242
rect 17773 25239 17831 25245
rect 15930 25208 15936 25220
rect 15856 25180 15936 25208
rect 12526 25100 12532 25152
rect 12584 25140 12590 25152
rect 13170 25140 13176 25152
rect 12584 25112 13176 25140
rect 12584 25100 12590 25112
rect 13170 25100 13176 25112
rect 13228 25140 13234 25152
rect 13725 25143 13783 25149
rect 13725 25140 13737 25143
rect 13228 25112 13737 25140
rect 13228 25100 13234 25112
rect 13725 25109 13737 25112
rect 13771 25140 13783 25143
rect 13998 25140 14004 25152
rect 13771 25112 14004 25140
rect 13771 25109 13783 25112
rect 13725 25103 13783 25109
rect 13998 25100 14004 25112
rect 14056 25100 14062 25152
rect 14734 25140 14740 25152
rect 14695 25112 14740 25140
rect 14734 25100 14740 25112
rect 14792 25100 14798 25152
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 15856 25140 15884 25180
rect 15930 25168 15936 25180
rect 15988 25168 15994 25220
rect 16206 25168 16212 25220
rect 16264 25208 16270 25220
rect 16637 25211 16695 25217
rect 16637 25208 16649 25211
rect 16264 25180 16649 25208
rect 16264 25168 16270 25180
rect 16637 25177 16649 25180
rect 16683 25177 16695 25211
rect 16637 25171 16695 25177
rect 16853 25211 16911 25217
rect 16853 25177 16865 25211
rect 16899 25177 16911 25211
rect 16853 25171 16911 25177
rect 16298 25140 16304 25152
rect 15243 25112 16304 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 16298 25100 16304 25112
rect 16356 25100 16362 25152
rect 16868 25140 16896 25171
rect 17678 25168 17684 25220
rect 17736 25208 17742 25220
rect 17788 25208 17816 25239
rect 17862 25236 17868 25288
rect 17920 25276 17926 25288
rect 17920 25248 17965 25276
rect 17920 25236 17926 25248
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 18509 25279 18567 25285
rect 18509 25276 18521 25279
rect 18288 25248 18521 25276
rect 18288 25236 18294 25248
rect 18509 25245 18521 25248
rect 18555 25245 18567 25279
rect 18601 25279 18659 25285
rect 18601 25266 18613 25279
rect 18647 25266 18659 25279
rect 18509 25239 18567 25245
rect 18598 25214 18604 25266
rect 18656 25214 18662 25266
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 18785 25279 18843 25285
rect 18785 25276 18797 25279
rect 18748 25248 18797 25276
rect 18748 25236 18754 25248
rect 18785 25245 18797 25248
rect 18831 25245 18843 25279
rect 18785 25239 18843 25245
rect 18877 25279 18935 25285
rect 18877 25245 18889 25279
rect 18923 25276 18935 25279
rect 18966 25276 18972 25288
rect 18923 25248 18972 25276
rect 18923 25245 18935 25248
rect 18877 25239 18935 25245
rect 17736 25180 17816 25208
rect 18800 25208 18828 25239
rect 18966 25236 18972 25248
rect 19024 25236 19030 25288
rect 19518 25236 19524 25288
rect 19576 25276 19582 25288
rect 20542 25279 20600 25285
rect 20542 25276 20554 25279
rect 19576 25248 20554 25276
rect 19576 25236 19582 25248
rect 20542 25245 20554 25248
rect 20588 25245 20600 25279
rect 20809 25279 20867 25285
rect 20809 25276 20821 25279
rect 20542 25239 20600 25245
rect 20640 25248 20821 25276
rect 19794 25208 19800 25220
rect 18800 25180 19800 25208
rect 17736 25168 17742 25180
rect 19794 25168 19800 25180
rect 19852 25168 19858 25220
rect 19978 25168 19984 25220
rect 20036 25208 20042 25220
rect 20640 25208 20668 25248
rect 20809 25245 20821 25248
rect 20855 25276 20867 25279
rect 21818 25276 21824 25288
rect 20855 25248 21824 25276
rect 20855 25245 20867 25248
rect 20809 25239 20867 25245
rect 21818 25236 21824 25248
rect 21876 25236 21882 25288
rect 22094 25236 22100 25288
rect 22152 25276 22158 25288
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 22152 25248 22661 25276
rect 22152 25236 22158 25248
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 22738 25236 22744 25288
rect 22796 25276 22802 25288
rect 23290 25276 23296 25288
rect 22796 25248 23296 25276
rect 22796 25236 22802 25248
rect 23290 25236 23296 25248
rect 23348 25236 23354 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25245 23443 25279
rect 23385 25239 23443 25245
rect 23569 25279 23627 25285
rect 23569 25245 23581 25279
rect 23615 25276 23627 25279
rect 23658 25276 23664 25288
rect 23615 25248 23664 25276
rect 23615 25245 23627 25248
rect 23569 25239 23627 25245
rect 20036 25180 20668 25208
rect 20036 25168 20042 25180
rect 20714 25168 20720 25220
rect 20772 25208 20778 25220
rect 22404 25211 22462 25217
rect 20772 25180 22094 25208
rect 20772 25168 20778 25180
rect 19058 25140 19064 25152
rect 16868 25112 19064 25140
rect 19058 25100 19064 25112
rect 19116 25100 19122 25152
rect 19426 25100 19432 25152
rect 19484 25140 19490 25152
rect 21269 25143 21327 25149
rect 21269 25140 21281 25143
rect 19484 25112 21281 25140
rect 19484 25100 19490 25112
rect 21269 25109 21281 25112
rect 21315 25109 21327 25143
rect 22066 25140 22094 25180
rect 22404 25177 22416 25211
rect 22450 25208 22462 25211
rect 23014 25208 23020 25220
rect 22450 25180 23020 25208
rect 22450 25177 22462 25180
rect 22404 25171 22462 25177
rect 23014 25168 23020 25180
rect 23072 25168 23078 25220
rect 23109 25143 23167 25149
rect 23109 25140 23121 25143
rect 22066 25112 23121 25140
rect 21269 25103 21327 25109
rect 23109 25109 23121 25112
rect 23155 25109 23167 25143
rect 23109 25103 23167 25109
rect 23290 25100 23296 25152
rect 23348 25140 23354 25152
rect 23400 25140 23428 25239
rect 23658 25236 23664 25248
rect 23716 25236 23722 25288
rect 24394 25236 24400 25288
rect 24452 25276 24458 25288
rect 25958 25276 25964 25288
rect 24452 25248 25964 25276
rect 24452 25236 24458 25248
rect 25958 25236 25964 25248
rect 26016 25236 26022 25288
rect 26528 25285 26556 25316
rect 27338 25304 27344 25316
rect 27396 25304 27402 25356
rect 27706 25344 27712 25356
rect 27448 25316 27712 25344
rect 26421 25279 26479 25285
rect 26421 25245 26433 25279
rect 26467 25245 26479 25279
rect 26421 25239 26479 25245
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25245 26571 25279
rect 26513 25239 26571 25245
rect 26697 25279 26755 25285
rect 26697 25245 26709 25279
rect 26743 25245 26755 25279
rect 26697 25239 26755 25245
rect 26789 25279 26847 25285
rect 26789 25245 26801 25279
rect 26835 25276 26847 25279
rect 27448 25276 27476 25316
rect 27706 25304 27712 25316
rect 27764 25304 27770 25356
rect 27614 25276 27620 25288
rect 26835 25248 27476 25276
rect 27575 25248 27620 25276
rect 26835 25245 26847 25248
rect 26789 25239 26847 25245
rect 25130 25168 25136 25220
rect 25188 25208 25194 25220
rect 25694 25211 25752 25217
rect 25694 25208 25706 25211
rect 25188 25180 25706 25208
rect 25188 25168 25194 25180
rect 25694 25177 25706 25180
rect 25740 25177 25752 25211
rect 26436 25208 26464 25239
rect 26602 25208 26608 25220
rect 26436 25180 26608 25208
rect 25694 25171 25752 25177
rect 26602 25168 26608 25180
rect 26660 25168 26666 25220
rect 23348 25112 23428 25140
rect 23348 25100 23354 25112
rect 23474 25100 23480 25152
rect 23532 25140 23538 25152
rect 24581 25143 24639 25149
rect 24581 25140 24593 25143
rect 23532 25112 24593 25140
rect 23532 25100 23538 25112
rect 24581 25109 24593 25112
rect 24627 25109 24639 25143
rect 24581 25103 24639 25109
rect 24946 25100 24952 25152
rect 25004 25140 25010 25152
rect 26712 25140 26740 25239
rect 27614 25236 27620 25248
rect 27672 25236 27678 25288
rect 27798 25236 27804 25288
rect 27856 25276 27862 25288
rect 27893 25279 27951 25285
rect 27893 25276 27905 25279
rect 27856 25248 27905 25276
rect 27856 25236 27862 25248
rect 27893 25245 27905 25248
rect 27939 25276 27951 25279
rect 27982 25276 27988 25288
rect 27939 25248 27988 25276
rect 27939 25245 27951 25248
rect 27893 25239 27951 25245
rect 27982 25236 27988 25248
rect 28040 25236 28046 25288
rect 27522 25208 27528 25220
rect 27448 25180 27528 25208
rect 25004 25112 26740 25140
rect 25004 25100 25010 25112
rect 27154 25100 27160 25152
rect 27212 25140 27218 25152
rect 27448 25149 27476 25180
rect 27522 25168 27528 25180
rect 27580 25168 27586 25220
rect 27433 25143 27491 25149
rect 27433 25140 27445 25143
rect 27212 25112 27445 25140
rect 27212 25100 27218 25112
rect 27433 25109 27445 25112
rect 27479 25109 27491 25143
rect 27798 25140 27804 25152
rect 27759 25112 27804 25140
rect 27433 25103 27491 25109
rect 27798 25100 27804 25112
rect 27856 25100 27862 25152
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 17218 24896 17224 24948
rect 17276 24936 17282 24948
rect 18233 24939 18291 24945
rect 17276 24908 18184 24936
rect 17276 24896 17282 24908
rect 13814 24828 13820 24880
rect 13872 24868 13878 24880
rect 14001 24871 14059 24877
rect 14001 24868 14013 24871
rect 13872 24840 14013 24868
rect 13872 24828 13878 24840
rect 14001 24837 14013 24840
rect 14047 24837 14059 24871
rect 16206 24868 16212 24880
rect 16167 24840 16212 24868
rect 14001 24831 14059 24837
rect 16206 24828 16212 24840
rect 16264 24868 16270 24880
rect 17465 24871 17523 24877
rect 17465 24868 17477 24871
rect 16264 24840 17477 24868
rect 16264 24828 16270 24840
rect 17465 24837 17477 24840
rect 17511 24837 17523 24871
rect 17465 24831 17523 24837
rect 17681 24871 17739 24877
rect 17681 24837 17693 24871
rect 17727 24868 17739 24871
rect 18046 24868 18052 24880
rect 17727 24840 18052 24868
rect 17727 24837 17739 24840
rect 17681 24831 17739 24837
rect 18046 24828 18052 24840
rect 18104 24828 18110 24880
rect 18156 24868 18184 24908
rect 18233 24905 18245 24939
rect 18279 24936 18291 24939
rect 18322 24936 18328 24948
rect 18279 24908 18328 24936
rect 18279 24905 18291 24908
rect 18233 24899 18291 24905
rect 18322 24896 18328 24908
rect 18380 24896 18386 24948
rect 19518 24896 19524 24948
rect 19576 24936 19582 24948
rect 21266 24936 21272 24948
rect 19576 24908 21272 24936
rect 19576 24896 19582 24908
rect 21266 24896 21272 24908
rect 21324 24896 21330 24948
rect 21453 24939 21511 24945
rect 21453 24905 21465 24939
rect 21499 24936 21511 24939
rect 25958 24936 25964 24948
rect 21499 24908 25964 24936
rect 21499 24905 21511 24908
rect 21453 24899 21511 24905
rect 25958 24896 25964 24908
rect 26016 24896 26022 24948
rect 26237 24939 26295 24945
rect 26237 24905 26249 24939
rect 26283 24936 26295 24939
rect 27062 24936 27068 24948
rect 26283 24908 27068 24936
rect 26283 24905 26295 24908
rect 26237 24899 26295 24905
rect 27062 24896 27068 24908
rect 27120 24896 27126 24948
rect 19702 24868 19708 24880
rect 18156 24840 18276 24868
rect 18248 24812 18276 24840
rect 19536 24840 19708 24868
rect 13354 24800 13360 24812
rect 13315 24772 13360 24800
rect 13354 24760 13360 24772
rect 13412 24760 13418 24812
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 13964 24772 15025 24800
rect 13964 24760 13970 24772
rect 15013 24769 15025 24772
rect 15059 24769 15071 24803
rect 15013 24763 15071 24769
rect 15028 24732 15056 24763
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 16298 24800 16304 24812
rect 15252 24772 16304 24800
rect 15252 24760 15258 24772
rect 16298 24760 16304 24772
rect 16356 24800 16362 24812
rect 18141 24803 18199 24809
rect 16356 24772 18000 24800
rect 18141 24790 18153 24803
rect 16356 24760 16362 24772
rect 17972 24732 18000 24772
rect 18064 24769 18153 24790
rect 18187 24769 18199 24803
rect 18064 24763 18199 24769
rect 18064 24762 18184 24763
rect 18064 24732 18092 24762
rect 18230 24760 18236 24812
rect 18288 24760 18294 24812
rect 18601 24804 18659 24809
rect 18601 24803 18828 24804
rect 18601 24769 18613 24803
rect 18647 24800 18828 24803
rect 18874 24800 18880 24812
rect 18647 24776 18880 24800
rect 18647 24772 18675 24776
rect 18800 24772 18880 24776
rect 18647 24769 18659 24772
rect 18601 24763 18659 24769
rect 18874 24760 18880 24772
rect 18932 24760 18938 24812
rect 19058 24800 19064 24812
rect 19019 24772 19064 24800
rect 19058 24760 19064 24772
rect 19116 24760 19122 24812
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24769 19303 24803
rect 19245 24763 19303 24769
rect 18417 24735 18475 24741
rect 15028 24704 17908 24732
rect 17972 24704 18276 24732
rect 14553 24667 14611 24673
rect 14553 24633 14565 24667
rect 14599 24664 14611 24667
rect 15194 24664 15200 24676
rect 14599 24636 15200 24664
rect 14599 24633 14611 24636
rect 14553 24627 14611 24633
rect 15194 24624 15200 24636
rect 15252 24624 15258 24676
rect 15378 24624 15384 24676
rect 15436 24664 15442 24676
rect 17313 24667 17371 24673
rect 17313 24664 17325 24667
rect 15436 24636 17325 24664
rect 15436 24624 15442 24636
rect 17313 24633 17325 24636
rect 17359 24633 17371 24667
rect 17313 24627 17371 24633
rect 15654 24596 15660 24608
rect 15615 24568 15660 24596
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 16666 24556 16672 24608
rect 16724 24596 16730 24608
rect 17218 24596 17224 24608
rect 16724 24568 17224 24596
rect 16724 24556 16730 24568
rect 17218 24556 17224 24568
rect 17276 24596 17282 24608
rect 17497 24599 17555 24605
rect 17497 24596 17509 24599
rect 17276 24568 17509 24596
rect 17276 24556 17282 24568
rect 17497 24565 17509 24568
rect 17543 24596 17555 24599
rect 17770 24596 17776 24608
rect 17543 24568 17776 24596
rect 17543 24565 17555 24568
rect 17497 24559 17555 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 17880 24596 17908 24704
rect 18248 24676 18276 24704
rect 18417 24701 18429 24735
rect 18463 24732 18475 24735
rect 18506 24732 18512 24744
rect 18463 24704 18512 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 18506 24692 18512 24704
rect 18564 24692 18570 24744
rect 18230 24624 18236 24676
rect 18288 24624 18294 24676
rect 18690 24624 18696 24676
rect 18748 24664 18754 24676
rect 19263 24664 19291 24763
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 19536 24809 19564 24840
rect 19702 24828 19708 24840
rect 19760 24868 19766 24880
rect 20318 24871 20376 24877
rect 19760 24840 20208 24868
rect 19760 24828 19766 24840
rect 19521 24803 19579 24809
rect 19392 24772 19437 24800
rect 19392 24760 19398 24772
rect 19521 24769 19533 24803
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 19623 24803 19681 24809
rect 19623 24769 19635 24803
rect 19669 24800 19681 24803
rect 20070 24800 20076 24812
rect 19669 24772 19932 24800
rect 20031 24772 20076 24800
rect 19669 24769 19681 24772
rect 19623 24763 19681 24769
rect 19904 24732 19932 24772
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20180 24800 20208 24840
rect 20318 24837 20330 24871
rect 20364 24868 20376 24871
rect 21358 24868 21364 24880
rect 20364 24840 21364 24868
rect 20364 24837 20376 24840
rect 20318 24831 20376 24837
rect 21358 24828 21364 24840
rect 21416 24828 21422 24880
rect 22462 24868 22468 24880
rect 22296 24840 22468 24868
rect 22296 24800 22324 24840
rect 22462 24828 22468 24840
rect 22520 24868 22526 24880
rect 22738 24868 22744 24880
rect 22520 24840 22744 24868
rect 22520 24828 22526 24840
rect 22738 24828 22744 24840
rect 22796 24828 22802 24880
rect 23198 24828 23204 24880
rect 23256 24868 23262 24880
rect 23256 24840 23428 24868
rect 23256 24828 23262 24840
rect 20180 24772 22324 24800
rect 22370 24760 22376 24812
rect 22428 24800 22434 24812
rect 23118 24803 23176 24809
rect 23118 24800 23130 24803
rect 22428 24772 23130 24800
rect 22428 24760 22434 24772
rect 23118 24769 23130 24772
rect 23164 24800 23176 24803
rect 23290 24800 23296 24812
rect 23164 24772 23296 24800
rect 23164 24769 23176 24772
rect 23118 24763 23176 24769
rect 23290 24760 23296 24772
rect 23348 24760 23354 24812
rect 23400 24809 23428 24840
rect 25590 24828 25596 24880
rect 25648 24868 25654 24880
rect 25648 24840 25912 24868
rect 25648 24828 25654 24840
rect 23385 24803 23443 24809
rect 23385 24769 23397 24803
rect 23431 24769 23443 24803
rect 23385 24763 23443 24769
rect 24946 24760 24952 24812
rect 25004 24809 25010 24812
rect 25004 24800 25016 24809
rect 25222 24800 25228 24812
rect 25004 24772 25049 24800
rect 25183 24772 25228 24800
rect 25004 24763 25016 24772
rect 25004 24760 25010 24763
rect 25222 24760 25228 24772
rect 25280 24760 25286 24812
rect 25884 24809 25912 24840
rect 26142 24828 26148 24880
rect 26200 24868 26206 24880
rect 26510 24868 26516 24880
rect 26200 24840 26516 24868
rect 26200 24828 26206 24840
rect 26510 24828 26516 24840
rect 26568 24828 26574 24880
rect 26694 24828 26700 24880
rect 26752 24868 26758 24880
rect 27309 24871 27367 24877
rect 27309 24868 27321 24871
rect 26752 24840 27321 24868
rect 26752 24828 26758 24840
rect 27309 24837 27321 24840
rect 27355 24837 27367 24871
rect 27522 24868 27528 24880
rect 27483 24840 27528 24868
rect 27309 24831 27367 24837
rect 27522 24828 27528 24840
rect 27580 24828 27586 24880
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24769 25835 24803
rect 25884 24803 25946 24809
rect 25884 24772 25900 24803
rect 25777 24763 25835 24769
rect 25888 24769 25900 24772
rect 25934 24769 25946 24803
rect 25888 24763 25946 24769
rect 26053 24803 26111 24809
rect 26053 24769 26065 24803
rect 26099 24800 26111 24803
rect 26878 24800 26884 24812
rect 26099 24772 26884 24800
rect 26099 24769 26111 24772
rect 26053 24763 26111 24769
rect 19904 24704 20116 24732
rect 19978 24664 19984 24676
rect 18748 24636 19984 24664
rect 18748 24624 18754 24636
rect 19978 24624 19984 24636
rect 20036 24624 20042 24676
rect 18322 24596 18328 24608
rect 17880 24568 18328 24596
rect 18322 24556 18328 24568
rect 18380 24596 18386 24608
rect 19334 24596 19340 24608
rect 18380 24568 19340 24596
rect 18380 24556 18386 24568
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 20088 24596 20116 24704
rect 25700 24664 25728 24763
rect 25792 24732 25820 24763
rect 26878 24760 26884 24772
rect 26936 24760 26942 24812
rect 27798 24760 27804 24812
rect 27856 24800 27862 24812
rect 27985 24803 28043 24809
rect 27985 24800 27997 24803
rect 27856 24772 27997 24800
rect 27856 24760 27862 24772
rect 27985 24769 27997 24772
rect 28031 24769 28043 24803
rect 27985 24763 28043 24769
rect 26970 24732 26976 24744
rect 25792 24704 26976 24732
rect 26970 24692 26976 24704
rect 27028 24692 27034 24744
rect 27430 24692 27436 24744
rect 27488 24692 27494 24744
rect 25958 24664 25964 24676
rect 21376 24636 22508 24664
rect 25700 24636 25964 24664
rect 21376 24596 21404 24636
rect 20088 24568 21404 24596
rect 21450 24556 21456 24608
rect 21508 24596 21514 24608
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21508 24568 22017 24596
rect 21508 24556 21514 24568
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22005 24559 22063 24565
rect 22186 24556 22192 24608
rect 22244 24596 22250 24608
rect 22370 24596 22376 24608
rect 22244 24568 22376 24596
rect 22244 24556 22250 24568
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 22480 24596 22508 24636
rect 25958 24624 25964 24636
rect 26016 24624 26022 24676
rect 26326 24624 26332 24676
rect 26384 24664 26390 24676
rect 27448 24664 27476 24692
rect 26384 24636 27476 24664
rect 26384 24624 26390 24636
rect 23198 24596 23204 24608
rect 22480 24568 23204 24596
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 23845 24599 23903 24605
rect 23845 24596 23857 24599
rect 23440 24568 23857 24596
rect 23440 24556 23446 24568
rect 23845 24565 23857 24568
rect 23891 24565 23903 24599
rect 23845 24559 23903 24565
rect 24578 24556 24584 24608
rect 24636 24596 24642 24608
rect 26050 24596 26056 24608
rect 24636 24568 26056 24596
rect 24636 24556 24642 24568
rect 26050 24556 26056 24568
rect 26108 24556 26114 24608
rect 27154 24596 27160 24608
rect 27115 24568 27160 24596
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 27246 24556 27252 24608
rect 27304 24596 27310 24608
rect 27341 24599 27399 24605
rect 27341 24596 27353 24599
rect 27304 24568 27353 24596
rect 27304 24556 27310 24568
rect 27341 24565 27353 24568
rect 27387 24565 27399 24599
rect 27341 24559 27399 24565
rect 27430 24556 27436 24608
rect 27488 24596 27494 24608
rect 27985 24599 28043 24605
rect 27985 24596 27997 24599
rect 27488 24568 27997 24596
rect 27488 24556 27494 24568
rect 27985 24565 27997 24568
rect 28031 24565 28043 24599
rect 27985 24559 28043 24565
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 14734 24352 14740 24404
rect 14792 24392 14798 24404
rect 15381 24395 15439 24401
rect 15381 24392 15393 24395
rect 14792 24364 15393 24392
rect 14792 24352 14798 24364
rect 15381 24361 15393 24364
rect 15427 24392 15439 24395
rect 15427 24364 16988 24392
rect 15427 24361 15439 24364
rect 15381 24355 15439 24361
rect 13262 24284 13268 24336
rect 13320 24324 13326 24336
rect 16758 24324 16764 24336
rect 13320 24296 16764 24324
rect 13320 24284 13326 24296
rect 16758 24284 16764 24296
rect 16816 24284 16822 24336
rect 13998 24216 14004 24268
rect 14056 24256 14062 24268
rect 14829 24259 14887 24265
rect 14829 24256 14841 24259
rect 14056 24228 14841 24256
rect 14056 24216 14062 24228
rect 14829 24225 14841 24228
rect 14875 24256 14887 24259
rect 16666 24256 16672 24268
rect 14875 24228 16672 24256
rect 14875 24225 14887 24228
rect 14829 24219 14887 24225
rect 16666 24216 16672 24228
rect 16724 24216 16730 24268
rect 16960 24256 16988 24364
rect 17126 24352 17132 24404
rect 17184 24392 17190 24404
rect 17865 24395 17923 24401
rect 17865 24392 17877 24395
rect 17184 24364 17877 24392
rect 17184 24352 17190 24364
rect 17865 24361 17877 24364
rect 17911 24361 17923 24395
rect 17865 24355 17923 24361
rect 17037 24327 17095 24333
rect 17037 24293 17049 24327
rect 17083 24324 17095 24327
rect 17218 24324 17224 24336
rect 17083 24296 17224 24324
rect 17083 24293 17095 24296
rect 17037 24287 17095 24293
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 17681 24327 17739 24333
rect 17681 24324 17693 24327
rect 17480 24296 17693 24324
rect 17310 24256 17316 24268
rect 16960 24228 17316 24256
rect 17310 24216 17316 24228
rect 17368 24216 17374 24268
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16206 24188 16212 24200
rect 15979 24160 16212 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 16206 24148 16212 24160
rect 16264 24188 16270 24200
rect 16485 24191 16543 24197
rect 16485 24188 16497 24191
rect 16264 24160 16497 24188
rect 16264 24148 16270 24160
rect 16485 24157 16497 24160
rect 16531 24188 16543 24191
rect 17218 24188 17224 24200
rect 16531 24160 17224 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 17218 24148 17224 24160
rect 17276 24148 17282 24200
rect 14274 24080 14280 24132
rect 14332 24120 14338 24132
rect 17480 24120 17508 24296
rect 17681 24293 17693 24296
rect 17727 24293 17739 24327
rect 17880 24324 17908 24355
rect 18598 24352 18604 24404
rect 18656 24392 18662 24404
rect 18693 24395 18751 24401
rect 18693 24392 18705 24395
rect 18656 24364 18705 24392
rect 18656 24352 18662 24364
rect 18693 24361 18705 24364
rect 18739 24361 18751 24395
rect 19613 24395 19671 24401
rect 19613 24392 19625 24395
rect 18693 24355 18751 24361
rect 18800 24364 19625 24392
rect 18800 24324 18828 24364
rect 19613 24361 19625 24364
rect 19659 24392 19671 24395
rect 19702 24392 19708 24404
rect 19659 24364 19708 24392
rect 19659 24361 19671 24364
rect 19613 24355 19671 24361
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 19797 24395 19855 24401
rect 19797 24361 19809 24395
rect 19843 24392 19855 24395
rect 23106 24392 23112 24404
rect 19843 24364 23112 24392
rect 19843 24361 19855 24364
rect 19797 24355 19855 24361
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 23566 24352 23572 24404
rect 23624 24392 23630 24404
rect 23661 24395 23719 24401
rect 23661 24392 23673 24395
rect 23624 24364 23673 24392
rect 23624 24352 23630 24364
rect 23661 24361 23673 24364
rect 23707 24361 23719 24395
rect 23661 24355 23719 24361
rect 24581 24395 24639 24401
rect 24581 24361 24593 24395
rect 24627 24392 24639 24395
rect 24854 24392 24860 24404
rect 24627 24364 24860 24392
rect 24627 24361 24639 24364
rect 24581 24355 24639 24361
rect 24854 24352 24860 24364
rect 24912 24352 24918 24404
rect 26605 24395 26663 24401
rect 26605 24392 26617 24395
rect 25056 24364 26617 24392
rect 17880 24296 18828 24324
rect 18877 24327 18935 24333
rect 17681 24287 17739 24293
rect 18877 24293 18889 24327
rect 18923 24293 18935 24327
rect 18877 24287 18935 24293
rect 18892 24256 18920 24287
rect 19058 24284 19064 24336
rect 19116 24324 19122 24336
rect 19886 24324 19892 24336
rect 19116 24296 19892 24324
rect 19116 24284 19122 24296
rect 19886 24284 19892 24296
rect 19944 24284 19950 24336
rect 20254 24324 20260 24336
rect 20215 24296 20260 24324
rect 20254 24284 20260 24296
rect 20312 24284 20318 24336
rect 20346 24284 20352 24336
rect 20404 24324 20410 24336
rect 21174 24324 21180 24336
rect 20404 24296 21180 24324
rect 20404 24284 20410 24296
rect 21174 24284 21180 24296
rect 21232 24284 21238 24336
rect 22649 24327 22707 24333
rect 22649 24293 22661 24327
rect 22695 24324 22707 24327
rect 22830 24324 22836 24336
rect 22695 24296 22836 24324
rect 22695 24293 22707 24296
rect 22649 24287 22707 24293
rect 22830 24284 22836 24296
rect 22888 24284 22894 24336
rect 22922 24284 22928 24336
rect 22980 24324 22986 24336
rect 25056 24324 25084 24364
rect 26605 24361 26617 24364
rect 26651 24361 26663 24395
rect 26786 24392 26792 24404
rect 26747 24364 26792 24392
rect 26605 24355 26663 24361
rect 26786 24352 26792 24364
rect 26844 24352 26850 24404
rect 27062 24352 27068 24404
rect 27120 24392 27126 24404
rect 27798 24392 27804 24404
rect 27120 24364 27804 24392
rect 27120 24352 27126 24364
rect 27798 24352 27804 24364
rect 27856 24352 27862 24404
rect 22980 24296 24348 24324
rect 22980 24284 22986 24296
rect 18892 24228 21404 24256
rect 19886 24188 19892 24200
rect 18432 24160 19892 24188
rect 18046 24129 18052 24132
rect 14332 24092 17508 24120
rect 18023 24123 18052 24129
rect 14332 24080 14338 24092
rect 18023 24089 18035 24123
rect 18104 24120 18110 24132
rect 18432 24120 18460 24160
rect 19886 24148 19892 24160
rect 19944 24148 19950 24200
rect 20070 24148 20076 24200
rect 20128 24188 20134 24200
rect 20433 24191 20491 24197
rect 20433 24188 20445 24191
rect 20128 24160 20445 24188
rect 20128 24148 20134 24160
rect 20433 24157 20445 24160
rect 20479 24157 20491 24191
rect 20433 24151 20491 24157
rect 20525 24191 20583 24197
rect 20525 24157 20537 24191
rect 20571 24188 20583 24191
rect 20714 24188 20720 24200
rect 20571 24157 20592 24188
rect 20675 24160 20720 24188
rect 20525 24151 20592 24157
rect 18104 24092 18460 24120
rect 18509 24123 18567 24129
rect 18023 24083 18052 24089
rect 18046 24080 18052 24083
rect 18104 24080 18110 24092
rect 18509 24089 18521 24123
rect 18555 24120 18567 24123
rect 19429 24123 19487 24129
rect 18555 24092 19389 24120
rect 18555 24089 18567 24092
rect 18509 24083 18567 24089
rect 16758 24012 16764 24064
rect 16816 24052 16822 24064
rect 17839 24055 17897 24061
rect 17839 24052 17851 24055
rect 16816 24024 17851 24052
rect 16816 24012 16822 24024
rect 17839 24021 17851 24024
rect 17885 24021 17897 24055
rect 17839 24015 17897 24021
rect 18709 24055 18767 24061
rect 18709 24021 18721 24055
rect 18755 24052 18767 24055
rect 19058 24052 19064 24064
rect 18755 24024 19064 24052
rect 18755 24021 18767 24024
rect 18709 24015 18767 24021
rect 19058 24012 19064 24024
rect 19116 24012 19122 24064
rect 19361 24052 19389 24092
rect 19429 24089 19441 24123
rect 19475 24120 19487 24123
rect 20162 24120 20168 24132
rect 19475 24092 20168 24120
rect 19475 24089 19487 24092
rect 19429 24083 19487 24089
rect 20162 24080 20168 24092
rect 20220 24080 20226 24132
rect 20564 24120 20592 24151
rect 20714 24148 20720 24160
rect 20772 24148 20778 24200
rect 20806 24148 20812 24200
rect 20864 24188 20870 24200
rect 21266 24188 21272 24200
rect 20864 24160 20909 24188
rect 21227 24160 21272 24188
rect 20864 24148 20870 24160
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 21376 24188 21404 24228
rect 23014 24216 23020 24268
rect 23072 24256 23078 24268
rect 23072 24228 23428 24256
rect 23072 24216 23078 24228
rect 23400 24197 23428 24228
rect 24320 24200 24348 24296
rect 24826 24296 25084 24324
rect 23109 24191 23167 24197
rect 23109 24188 23121 24191
rect 21376 24160 23121 24188
rect 23109 24157 23121 24160
rect 23155 24157 23167 24191
rect 23109 24151 23167 24157
rect 23201 24191 23259 24197
rect 23201 24157 23213 24191
rect 23247 24157 23259 24191
rect 23201 24151 23259 24157
rect 23385 24191 23443 24197
rect 23385 24157 23397 24191
rect 23431 24157 23443 24191
rect 23385 24151 23443 24157
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 23566 24188 23572 24200
rect 23523 24160 23572 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 20622 24120 20628 24132
rect 20564 24092 20628 24120
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 21174 24080 21180 24132
rect 21232 24120 21238 24132
rect 21514 24123 21572 24129
rect 21514 24120 21526 24123
rect 21232 24092 21526 24120
rect 21232 24080 21238 24092
rect 21514 24089 21526 24092
rect 21560 24089 21572 24123
rect 21514 24083 21572 24089
rect 21634 24080 21640 24132
rect 21692 24120 21698 24132
rect 23216 24120 23244 24151
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 24826 24188 24854 24296
rect 27982 24284 27988 24336
rect 28040 24324 28046 24336
rect 28077 24327 28135 24333
rect 28077 24324 28089 24327
rect 28040 24296 28089 24324
rect 28040 24284 28046 24296
rect 28077 24293 28089 24296
rect 28123 24293 28135 24327
rect 28077 24287 28135 24293
rect 24946 24216 24952 24268
rect 25004 24216 25010 24268
rect 24360 24160 24854 24188
rect 24964 24188 24992 24216
rect 25958 24188 25964 24200
rect 24964 24160 25820 24188
rect 25919 24160 25964 24188
rect 24360 24148 24366 24160
rect 21692 24092 24808 24120
rect 21692 24080 21698 24092
rect 19518 24052 19524 24064
rect 19361 24024 19524 24052
rect 19518 24012 19524 24024
rect 19576 24012 19582 24064
rect 19639 24055 19697 24061
rect 19639 24021 19651 24055
rect 19685 24052 19697 24055
rect 19794 24052 19800 24064
rect 19685 24024 19800 24052
rect 19685 24021 19697 24024
rect 19639 24015 19697 24021
rect 19794 24012 19800 24024
rect 19852 24012 19858 24064
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 23474 24052 23480 24064
rect 19944 24024 23480 24052
rect 19944 24012 19950 24024
rect 23474 24012 23480 24024
rect 23532 24012 23538 24064
rect 24780 24052 24808 24092
rect 25590 24080 25596 24132
rect 25648 24120 25654 24132
rect 25694 24123 25752 24129
rect 25694 24120 25706 24123
rect 25648 24092 25706 24120
rect 25648 24080 25654 24092
rect 25694 24089 25706 24092
rect 25740 24089 25752 24123
rect 25792 24120 25820 24160
rect 25958 24148 25964 24160
rect 26016 24148 26022 24200
rect 26326 24188 26332 24200
rect 26068 24160 26332 24188
rect 26068 24120 26096 24160
rect 26326 24148 26332 24160
rect 26384 24148 26390 24200
rect 27433 24191 27491 24197
rect 27433 24157 27445 24191
rect 27479 24188 27491 24191
rect 27522 24188 27528 24200
rect 27479 24160 27528 24188
rect 27479 24157 27491 24160
rect 27433 24151 27491 24157
rect 27522 24148 27528 24160
rect 27580 24148 27586 24200
rect 26418 24120 26424 24132
rect 25792 24092 26096 24120
rect 26379 24092 26424 24120
rect 25694 24083 25752 24089
rect 26418 24080 26424 24092
rect 26476 24080 26482 24132
rect 26510 24080 26516 24132
rect 26568 24120 26574 24132
rect 27249 24123 27307 24129
rect 27249 24120 27261 24123
rect 26568 24092 27261 24120
rect 26568 24080 26574 24092
rect 27249 24089 27261 24092
rect 27295 24089 27307 24123
rect 27249 24083 27307 24089
rect 27798 24080 27804 24132
rect 27856 24120 27862 24132
rect 28258 24120 28264 24132
rect 27856 24092 28264 24120
rect 27856 24080 27862 24092
rect 28258 24080 28264 24092
rect 28316 24080 28322 24132
rect 26234 24052 26240 24064
rect 24780 24024 26240 24052
rect 26234 24012 26240 24024
rect 26292 24012 26298 24064
rect 26326 24012 26332 24064
rect 26384 24052 26390 24064
rect 26621 24055 26679 24061
rect 26621 24052 26633 24055
rect 26384 24024 26633 24052
rect 26384 24012 26390 24024
rect 26621 24021 26633 24024
rect 26667 24021 26679 24055
rect 26621 24015 26679 24021
rect 26786 24012 26792 24064
rect 26844 24052 26850 24064
rect 27614 24052 27620 24064
rect 26844 24024 27620 24052
rect 26844 24012 26850 24024
rect 27614 24012 27620 24024
rect 27672 24012 27678 24064
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 15197 23851 15255 23857
rect 15197 23817 15209 23851
rect 15243 23848 15255 23851
rect 16390 23848 16396 23860
rect 15243 23820 16396 23848
rect 15243 23817 15255 23820
rect 15197 23811 15255 23817
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 17221 23851 17279 23857
rect 17221 23817 17233 23851
rect 17267 23848 17279 23851
rect 17310 23848 17316 23860
rect 17267 23820 17316 23848
rect 17267 23817 17279 23820
rect 17221 23811 17279 23817
rect 17310 23808 17316 23820
rect 17368 23848 17374 23860
rect 18690 23848 18696 23860
rect 17368 23820 18696 23848
rect 17368 23808 17374 23820
rect 18690 23808 18696 23820
rect 18748 23808 18754 23860
rect 19150 23808 19156 23860
rect 19208 23848 19214 23860
rect 20806 23848 20812 23860
rect 19208 23820 20812 23848
rect 19208 23808 19214 23820
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 23566 23848 23572 23860
rect 21100 23820 23572 23848
rect 12710 23740 12716 23792
rect 12768 23780 12774 23792
rect 17126 23780 17132 23792
rect 12768 23752 17132 23780
rect 12768 23740 12774 23752
rect 17126 23740 17132 23752
rect 17184 23780 17190 23792
rect 17865 23783 17923 23789
rect 17865 23780 17877 23783
rect 17184 23752 17877 23780
rect 17184 23740 17190 23752
rect 17865 23749 17877 23752
rect 17911 23749 17923 23783
rect 17865 23743 17923 23749
rect 17954 23740 17960 23792
rect 18012 23780 18018 23792
rect 18417 23783 18475 23789
rect 18417 23780 18429 23783
rect 18012 23752 18429 23780
rect 18012 23740 18018 23752
rect 18417 23749 18429 23752
rect 18463 23749 18475 23783
rect 18417 23743 18475 23749
rect 18601 23783 18659 23789
rect 18601 23749 18613 23783
rect 18647 23780 18659 23783
rect 18782 23780 18788 23792
rect 18647 23752 18788 23780
rect 18647 23749 18659 23752
rect 18601 23743 18659 23749
rect 18782 23740 18788 23752
rect 18840 23740 18846 23792
rect 19058 23740 19064 23792
rect 19116 23780 19122 23792
rect 19305 23783 19363 23789
rect 19305 23780 19317 23783
rect 19116 23752 19317 23780
rect 19116 23740 19122 23752
rect 19305 23749 19317 23752
rect 19351 23749 19363 23783
rect 19305 23743 19363 23749
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 19521 23783 19579 23789
rect 19521 23780 19533 23783
rect 19484 23752 19533 23780
rect 19484 23740 19490 23752
rect 19521 23749 19533 23752
rect 19567 23749 19579 23783
rect 19521 23743 19579 23749
rect 20073 23783 20131 23789
rect 20073 23749 20085 23783
rect 20119 23780 20131 23783
rect 20162 23780 20168 23792
rect 20119 23752 20168 23780
rect 20119 23749 20131 23752
rect 20073 23743 20131 23749
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 20346 23740 20352 23792
rect 20404 23780 20410 23792
rect 21100 23780 21128 23820
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 25498 23848 25504 23860
rect 24228 23820 25504 23848
rect 23842 23780 23848 23792
rect 20404 23752 21128 23780
rect 20404 23740 20410 23752
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 16209 23715 16267 23721
rect 16209 23712 16221 23715
rect 9824 23684 16221 23712
rect 9824 23672 9830 23684
rect 16209 23681 16221 23684
rect 16255 23712 16267 23715
rect 16666 23712 16672 23724
rect 16255 23684 16672 23712
rect 16255 23681 16267 23684
rect 16209 23675 16267 23681
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 16942 23672 16948 23724
rect 17000 23712 17006 23724
rect 19978 23712 19984 23724
rect 17000 23684 19840 23712
rect 19939 23684 19984 23712
rect 17000 23672 17006 23684
rect 14182 23604 14188 23656
rect 14240 23644 14246 23656
rect 15749 23647 15807 23653
rect 15749 23644 15761 23647
rect 14240 23616 15761 23644
rect 14240 23604 14246 23616
rect 15749 23613 15761 23616
rect 15795 23644 15807 23647
rect 19518 23644 19524 23656
rect 15795 23616 19524 23644
rect 15795 23613 15807 23616
rect 15749 23607 15807 23613
rect 19518 23604 19524 23616
rect 19576 23604 19582 23656
rect 19153 23579 19211 23585
rect 19153 23576 19165 23579
rect 17519 23548 19165 23576
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 16022 23468 16028 23520
rect 16080 23508 16086 23520
rect 17519 23508 17547 23548
rect 19153 23545 19165 23548
rect 19199 23545 19211 23579
rect 19812 23576 19840 23684
rect 19978 23672 19984 23684
rect 20036 23672 20042 23724
rect 20254 23712 20260 23724
rect 20215 23684 20260 23712
rect 20254 23672 20260 23684
rect 20312 23672 20318 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23712 20499 23715
rect 20622 23712 20628 23724
rect 20487 23684 20628 23712
rect 20487 23681 20499 23684
rect 20441 23675 20499 23681
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 20898 23672 20904 23724
rect 20956 23672 20962 23724
rect 21100 23721 21128 23752
rect 21836 23752 23848 23780
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 21174 23672 21180 23724
rect 21232 23712 21238 23724
rect 21358 23721 21364 23724
rect 21346 23715 21364 23721
rect 21232 23684 21277 23712
rect 21232 23672 21238 23684
rect 21346 23681 21358 23715
rect 21346 23675 21364 23681
rect 21358 23672 21364 23675
rect 21416 23672 21422 23724
rect 21450 23672 21456 23724
rect 21508 23712 21514 23724
rect 21836 23712 21864 23752
rect 23842 23740 23848 23752
rect 23900 23740 23906 23792
rect 21508 23684 21553 23712
rect 21652 23684 21864 23712
rect 21508 23672 21514 23684
rect 19886 23604 19892 23656
rect 19944 23644 19950 23656
rect 20916 23644 20944 23672
rect 21542 23644 21548 23656
rect 19944 23616 21548 23644
rect 19944 23604 19950 23616
rect 21542 23604 21548 23616
rect 21600 23604 21606 23656
rect 20901 23579 20959 23585
rect 19812 23548 20852 23576
rect 19153 23539 19211 23545
rect 16080 23480 17547 23508
rect 16080 23468 16086 23480
rect 17770 23468 17776 23520
rect 17828 23508 17834 23520
rect 17954 23508 17960 23520
rect 17828 23480 17960 23508
rect 17828 23468 17834 23480
rect 17954 23468 17960 23480
rect 18012 23508 18018 23520
rect 18598 23508 18604 23520
rect 18012 23480 18604 23508
rect 18012 23468 18018 23480
rect 18598 23468 18604 23480
rect 18656 23508 18662 23520
rect 19337 23511 19395 23517
rect 19337 23508 19349 23511
rect 18656 23480 19349 23508
rect 18656 23468 18662 23480
rect 19337 23477 19349 23480
rect 19383 23508 19395 23511
rect 19886 23508 19892 23520
rect 19383 23480 19892 23508
rect 19383 23477 19395 23480
rect 19337 23471 19395 23477
rect 19886 23468 19892 23480
rect 19944 23468 19950 23520
rect 20824 23508 20852 23548
rect 20901 23545 20913 23579
rect 20947 23576 20959 23579
rect 21652 23576 21680 23684
rect 21910 23672 21916 23724
rect 21968 23712 21974 23724
rect 22261 23715 22319 23721
rect 22261 23712 22273 23715
rect 21968 23684 22273 23712
rect 21968 23672 21974 23684
rect 22261 23681 22273 23684
rect 22307 23681 22319 23715
rect 22261 23675 22319 23681
rect 22554 23672 22560 23724
rect 22612 23712 22618 23724
rect 22612 23684 23060 23712
rect 22612 23672 22618 23684
rect 21726 23604 21732 23656
rect 21784 23644 21790 23656
rect 22002 23644 22008 23656
rect 21784 23616 22008 23644
rect 21784 23604 21790 23616
rect 22002 23604 22008 23616
rect 22060 23604 22066 23656
rect 23032 23644 23060 23684
rect 23474 23644 23480 23656
rect 23032 23616 23480 23644
rect 23474 23604 23480 23616
rect 23532 23604 23538 23656
rect 24228 23576 24256 23820
rect 25498 23808 25504 23820
rect 25556 23808 25562 23860
rect 25685 23851 25743 23857
rect 25685 23817 25697 23851
rect 25731 23848 25743 23851
rect 27522 23848 27528 23860
rect 25731 23820 27528 23848
rect 25731 23817 25743 23820
rect 25685 23811 25743 23817
rect 27522 23808 27528 23820
rect 27580 23808 27586 23860
rect 24854 23780 24860 23792
rect 24826 23740 24860 23780
rect 24912 23740 24918 23792
rect 24980 23783 25038 23789
rect 24980 23749 24992 23783
rect 25026 23780 25038 23783
rect 27430 23780 27436 23792
rect 25026 23752 27436 23780
rect 25026 23749 25038 23752
rect 24980 23743 25038 23749
rect 27430 23740 27436 23752
rect 27488 23740 27494 23792
rect 28166 23780 28172 23792
rect 27724 23752 28172 23780
rect 24578 23672 24584 23724
rect 24636 23712 24642 23724
rect 24826 23712 24854 23740
rect 25225 23715 25283 23721
rect 25225 23712 25237 23715
rect 24636 23684 25237 23712
rect 24636 23672 24642 23684
rect 25225 23681 25237 23684
rect 25271 23681 25283 23715
rect 25225 23675 25283 23681
rect 25869 23715 25927 23721
rect 25869 23681 25881 23715
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 26053 23715 26111 23721
rect 26053 23681 26065 23715
rect 26099 23712 26111 23715
rect 26234 23712 26240 23724
rect 26099 23684 26240 23712
rect 26099 23681 26111 23684
rect 26053 23675 26111 23681
rect 25884 23644 25912 23675
rect 26234 23672 26240 23684
rect 26292 23672 26298 23724
rect 26605 23715 26663 23721
rect 26605 23681 26617 23715
rect 26651 23712 26663 23715
rect 26970 23712 26976 23724
rect 26651 23684 26976 23712
rect 26651 23681 26663 23684
rect 26605 23675 26663 23681
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 27614 23672 27620 23724
rect 27672 23712 27678 23724
rect 27724 23721 27752 23752
rect 28166 23740 28172 23752
rect 28224 23740 28230 23792
rect 27709 23715 27767 23721
rect 27709 23712 27721 23715
rect 27672 23684 27721 23712
rect 27672 23672 27678 23684
rect 27709 23681 27721 23684
rect 27755 23681 27767 23715
rect 28350 23712 28356 23724
rect 28311 23684 28356 23712
rect 27709 23675 27767 23681
rect 28350 23672 28356 23684
rect 28408 23672 28414 23724
rect 28166 23644 28172 23656
rect 25884 23616 28172 23644
rect 28166 23604 28172 23616
rect 28224 23604 28230 23656
rect 27062 23576 27068 23588
rect 20947 23548 21680 23576
rect 23400 23548 24256 23576
rect 26436 23548 27068 23576
rect 20947 23545 20959 23548
rect 20901 23539 20959 23545
rect 23400 23517 23428 23548
rect 23385 23511 23443 23517
rect 23385 23508 23397 23511
rect 20824 23480 23397 23508
rect 23385 23477 23397 23480
rect 23431 23477 23443 23511
rect 23842 23508 23848 23520
rect 23755 23480 23848 23508
rect 23385 23471 23443 23477
rect 23842 23468 23848 23480
rect 23900 23508 23906 23520
rect 26436 23508 26464 23548
rect 27062 23536 27068 23548
rect 27120 23536 27126 23588
rect 23900 23480 26464 23508
rect 23900 23468 23906 23480
rect 26602 23468 26608 23520
rect 26660 23508 26666 23520
rect 27525 23511 27583 23517
rect 27525 23508 27537 23511
rect 26660 23480 27537 23508
rect 26660 23468 26666 23480
rect 27525 23477 27537 23480
rect 27571 23477 27583 23511
rect 27525 23471 27583 23477
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 16209 23307 16267 23313
rect 16209 23273 16221 23307
rect 16255 23304 16267 23307
rect 16298 23304 16304 23316
rect 16255 23276 16304 23304
rect 16255 23273 16267 23276
rect 16209 23267 16267 23273
rect 16298 23264 16304 23276
rect 16356 23264 16362 23316
rect 16758 23304 16764 23316
rect 16719 23276 16764 23304
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 17865 23307 17923 23313
rect 17865 23273 17877 23307
rect 17911 23304 17923 23307
rect 17954 23304 17960 23316
rect 17911 23276 17960 23304
rect 17911 23273 17923 23276
rect 17865 23267 17923 23273
rect 17954 23264 17960 23276
rect 18012 23264 18018 23316
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 19705 23307 19763 23313
rect 19705 23304 19717 23307
rect 19392 23276 19717 23304
rect 19392 23264 19398 23276
rect 19705 23273 19717 23276
rect 19751 23304 19763 23307
rect 20254 23304 20260 23316
rect 19751 23276 20260 23304
rect 19751 23273 19763 23276
rect 19705 23267 19763 23273
rect 20254 23264 20260 23276
rect 20312 23264 20318 23316
rect 20530 23313 20536 23316
rect 20524 23304 20536 23313
rect 20491 23276 20536 23304
rect 20524 23267 20536 23276
rect 20530 23264 20536 23267
rect 20588 23264 20594 23316
rect 20717 23307 20775 23313
rect 20717 23273 20729 23307
rect 20763 23304 20775 23307
rect 21818 23304 21824 23316
rect 20763 23276 21824 23304
rect 20763 23273 20775 23276
rect 20717 23267 20775 23273
rect 21818 23264 21824 23276
rect 21876 23264 21882 23316
rect 23750 23304 23756 23316
rect 22664 23276 23756 23304
rect 16776 23236 16804 23264
rect 18325 23239 18383 23245
rect 18325 23236 18337 23239
rect 16776 23208 18337 23236
rect 18325 23205 18337 23208
rect 18371 23236 18383 23239
rect 19794 23236 19800 23248
rect 18371 23208 19800 23236
rect 18371 23205 18383 23208
rect 18325 23199 18383 23205
rect 19794 23196 19800 23208
rect 19852 23236 19858 23248
rect 20162 23236 20168 23248
rect 19852 23208 20168 23236
rect 19852 23196 19858 23208
rect 20162 23196 20168 23208
rect 20220 23196 20226 23248
rect 20438 23196 20444 23248
rect 20496 23236 20502 23248
rect 22189 23239 22247 23245
rect 22189 23236 22201 23239
rect 20496 23208 22201 23236
rect 20496 23196 20502 23208
rect 22189 23205 22201 23208
rect 22235 23236 22247 23239
rect 22664 23236 22692 23276
rect 23750 23264 23756 23276
rect 23808 23264 23814 23316
rect 24118 23264 24124 23316
rect 24176 23304 24182 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 24176 23276 24777 23304
rect 24176 23264 24182 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 25038 23264 25044 23316
rect 25096 23304 25102 23316
rect 25222 23304 25228 23316
rect 25096 23276 25228 23304
rect 25096 23264 25102 23276
rect 25222 23264 25228 23276
rect 25280 23264 25286 23316
rect 25593 23307 25651 23313
rect 25593 23273 25605 23307
rect 25639 23304 25651 23307
rect 27154 23304 27160 23316
rect 25639 23276 27160 23304
rect 25639 23273 25651 23276
rect 25593 23267 25651 23273
rect 27154 23264 27160 23276
rect 27212 23264 27218 23316
rect 27706 23304 27712 23316
rect 27667 23276 27712 23304
rect 27706 23264 27712 23276
rect 27764 23264 27770 23316
rect 22235 23208 22692 23236
rect 22235 23205 22247 23208
rect 22189 23199 22247 23205
rect 25682 23196 25688 23248
rect 25740 23236 25746 23248
rect 25777 23239 25835 23245
rect 25777 23236 25789 23239
rect 25740 23208 25789 23236
rect 25740 23196 25746 23208
rect 25777 23205 25789 23208
rect 25823 23205 25835 23239
rect 25777 23199 25835 23205
rect 25866 23196 25872 23248
rect 25924 23236 25930 23248
rect 26421 23239 26479 23245
rect 26421 23236 26433 23239
rect 25924 23208 26433 23236
rect 25924 23196 25930 23208
rect 26421 23205 26433 23208
rect 26467 23236 26479 23239
rect 26786 23236 26792 23248
rect 26467 23208 26792 23236
rect 26467 23205 26479 23208
rect 26421 23199 26479 23205
rect 26786 23196 26792 23208
rect 26844 23196 26850 23248
rect 17586 23128 17592 23180
rect 17644 23168 17650 23180
rect 21177 23171 21235 23177
rect 21177 23168 21189 23171
rect 17644 23140 21189 23168
rect 17644 23128 17650 23140
rect 21177 23137 21189 23140
rect 21223 23137 21235 23171
rect 21177 23131 21235 23137
rect 21266 23128 21272 23180
rect 21324 23168 21330 23180
rect 21910 23168 21916 23180
rect 21324 23140 21916 23168
rect 21324 23128 21330 23140
rect 18046 23060 18052 23112
rect 18104 23100 18110 23112
rect 18104 23072 20392 23100
rect 18104 23060 18110 23072
rect 18138 22992 18144 23044
rect 18196 23032 18202 23044
rect 20364 23041 20392 23072
rect 20898 23060 20904 23112
rect 20956 23100 20962 23112
rect 21468 23109 21496 23140
rect 21910 23128 21916 23140
rect 21968 23128 21974 23180
rect 21361 23103 21419 23109
rect 21361 23100 21373 23103
rect 20956 23072 21373 23100
rect 20956 23060 20962 23072
rect 21192 23044 21220 23072
rect 21361 23069 21373 23072
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 21453 23103 21511 23109
rect 21453 23069 21465 23103
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 21637 23103 21695 23109
rect 21637 23069 21649 23103
rect 21683 23069 21695 23103
rect 21637 23063 21695 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22186 23100 22192 23112
rect 21775 23072 22192 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 19889 23035 19947 23041
rect 19889 23032 19901 23035
rect 18196 23004 19901 23032
rect 18196 22992 18202 23004
rect 19889 23001 19901 23004
rect 19935 23001 19947 23035
rect 19889 22995 19947 23001
rect 20349 23035 20407 23041
rect 20349 23001 20361 23035
rect 20395 23001 20407 23035
rect 20349 22995 20407 23001
rect 20714 22992 20720 23044
rect 20772 23032 20778 23044
rect 20772 23004 20944 23032
rect 20772 22992 20778 23004
rect 17310 22964 17316 22976
rect 17271 22936 17316 22964
rect 17310 22924 17316 22936
rect 17368 22924 17374 22976
rect 19518 22964 19524 22976
rect 19479 22936 19524 22964
rect 19518 22924 19524 22936
rect 19576 22924 19582 22976
rect 19689 22967 19747 22973
rect 19689 22933 19701 22967
rect 19735 22964 19747 22967
rect 19978 22964 19984 22976
rect 19735 22936 19984 22964
rect 19735 22933 19747 22936
rect 19689 22927 19747 22933
rect 19978 22924 19984 22936
rect 20036 22924 20042 22976
rect 20162 22924 20168 22976
rect 20220 22964 20226 22976
rect 20438 22964 20444 22976
rect 20220 22936 20444 22964
rect 20220 22924 20226 22936
rect 20438 22924 20444 22936
rect 20496 22964 20502 22976
rect 20549 22967 20607 22973
rect 20549 22964 20561 22967
rect 20496 22936 20561 22964
rect 20496 22924 20502 22936
rect 20549 22933 20561 22936
rect 20595 22964 20607 22967
rect 20806 22964 20812 22976
rect 20595 22936 20812 22964
rect 20595 22933 20607 22936
rect 20549 22927 20607 22933
rect 20806 22924 20812 22936
rect 20864 22924 20870 22976
rect 20916 22964 20944 23004
rect 21174 22992 21180 23044
rect 21232 22992 21238 23044
rect 21652 23032 21680 23063
rect 22186 23060 22192 23072
rect 22244 23060 22250 23112
rect 23569 23103 23627 23109
rect 23569 23069 23581 23103
rect 23615 23100 23627 23103
rect 23842 23100 23848 23112
rect 23615 23072 23848 23100
rect 23615 23069 23627 23072
rect 23569 23063 23627 23069
rect 23842 23060 23848 23072
rect 23900 23060 23906 23112
rect 26234 23100 26240 23112
rect 25148 23072 25737 23100
rect 26195 23072 26240 23100
rect 25148 23066 25176 23072
rect 21818 23032 21824 23044
rect 21652 23004 21824 23032
rect 21818 22992 21824 23004
rect 21876 22992 21882 23044
rect 23324 23035 23382 23041
rect 23324 23001 23336 23035
rect 23370 23032 23382 23035
rect 24486 23032 24492 23044
rect 23370 23004 24492 23032
rect 23370 23001 23382 23004
rect 23324 22995 23382 23001
rect 24486 22992 24492 23004
rect 24544 22992 24550 23044
rect 24581 23035 24639 23041
rect 24581 23001 24593 23035
rect 24627 23032 24639 23035
rect 24670 23032 24676 23044
rect 24627 23004 24676 23032
rect 24627 23001 24639 23004
rect 24581 22995 24639 23001
rect 24670 22992 24676 23004
rect 24728 22992 24734 23044
rect 24826 23038 25176 23066
rect 23106 22964 23112 22976
rect 20916 22936 23112 22964
rect 23106 22924 23112 22936
rect 23164 22924 23170 22976
rect 23198 22924 23204 22976
rect 23256 22964 23262 22976
rect 24826 22973 24854 23038
rect 25406 23032 25412 23044
rect 25367 23004 25412 23032
rect 25406 22992 25412 23004
rect 25464 22992 25470 23044
rect 25498 22992 25504 23044
rect 25556 23032 25562 23044
rect 25609 23035 25667 23041
rect 25609 23032 25621 23035
rect 25556 23004 25621 23032
rect 25556 22992 25562 23004
rect 25609 23001 25621 23004
rect 25655 23001 25667 23035
rect 25609 22995 25667 23001
rect 24791 22967 24854 22973
rect 24791 22964 24803 22967
rect 23256 22936 24803 22964
rect 23256 22924 23262 22936
rect 24791 22933 24803 22936
rect 24837 22936 24854 22967
rect 24837 22933 24849 22936
rect 24791 22927 24849 22933
rect 24946 22924 24952 22976
rect 25004 22964 25010 22976
rect 25709 22964 25737 23072
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 26421 23103 26479 23109
rect 26421 23069 26433 23103
rect 26467 23100 26479 23103
rect 26602 23100 26608 23112
rect 26467 23072 26608 23100
rect 26467 23069 26479 23072
rect 26421 23063 26479 23069
rect 26602 23060 26608 23072
rect 26660 23060 26666 23112
rect 27062 23100 27068 23112
rect 27023 23072 27068 23100
rect 27062 23060 27068 23072
rect 27120 23060 27126 23112
rect 28350 23100 28356 23112
rect 28311 23072 28356 23100
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 26418 22964 26424 22976
rect 25004 22936 25049 22964
rect 25709 22936 26424 22964
rect 25004 22924 25010 22936
rect 26418 22924 26424 22936
rect 26476 22924 26482 22976
rect 26878 22964 26884 22976
rect 26839 22936 26884 22964
rect 26878 22924 26884 22936
rect 26936 22924 26942 22976
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 16390 22720 16396 22772
rect 16448 22760 16454 22772
rect 16853 22763 16911 22769
rect 16853 22760 16865 22763
rect 16448 22732 16865 22760
rect 16448 22720 16454 22732
rect 16853 22729 16865 22732
rect 16899 22729 16911 22763
rect 16853 22723 16911 22729
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 18049 22763 18107 22769
rect 18049 22760 18061 22763
rect 17276 22732 18061 22760
rect 17276 22720 17282 22732
rect 18049 22729 18061 22732
rect 18095 22760 18107 22763
rect 18966 22760 18972 22772
rect 18095 22732 18972 22760
rect 18095 22729 18107 22732
rect 18049 22723 18107 22729
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 19061 22763 19119 22769
rect 19061 22729 19073 22763
rect 19107 22760 19119 22763
rect 19794 22760 19800 22772
rect 19107 22732 19656 22760
rect 19707 22732 19800 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19628 22692 19656 22732
rect 19794 22720 19800 22732
rect 19852 22760 19858 22772
rect 20254 22760 20260 22772
rect 19852 22732 20260 22760
rect 19852 22720 19858 22732
rect 20254 22720 20260 22732
rect 20312 22720 20318 22772
rect 20898 22720 20904 22772
rect 20956 22760 20962 22772
rect 21285 22763 21343 22769
rect 21285 22760 21297 22763
rect 20956 22732 21297 22760
rect 20956 22720 20962 22732
rect 21285 22729 21297 22732
rect 21331 22729 21343 22763
rect 21285 22723 21343 22729
rect 21453 22763 21511 22769
rect 21453 22729 21465 22763
rect 21499 22760 21511 22763
rect 22094 22760 22100 22772
rect 21499 22732 22100 22760
rect 21499 22729 21511 22732
rect 21453 22723 21511 22729
rect 22094 22720 22100 22732
rect 22152 22720 22158 22772
rect 22204 22732 22416 22760
rect 19886 22692 19892 22704
rect 19628 22664 19892 22692
rect 19886 22652 19892 22664
rect 19944 22652 19950 22704
rect 20438 22701 20444 22704
rect 20425 22695 20444 22701
rect 20425 22661 20437 22695
rect 20425 22655 20444 22661
rect 20438 22652 20444 22655
rect 20496 22652 20502 22704
rect 20625 22695 20683 22701
rect 20625 22661 20637 22695
rect 20671 22692 20683 22695
rect 20714 22692 20720 22704
rect 20671 22664 20720 22692
rect 20671 22661 20683 22664
rect 20625 22655 20683 22661
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 21082 22692 21088 22704
rect 21043 22664 21088 22692
rect 21082 22652 21088 22664
rect 21140 22652 21146 22704
rect 21818 22584 21824 22636
rect 21876 22624 21882 22636
rect 21995 22633 22053 22639
rect 21995 22630 22007 22633
rect 21928 22624 22007 22630
rect 21876 22602 22007 22624
rect 21876 22596 21956 22602
rect 21876 22584 21882 22596
rect 17494 22516 17500 22568
rect 17552 22556 17558 22568
rect 21928 22556 21956 22596
rect 21995 22599 22007 22602
rect 22041 22599 22053 22633
rect 21995 22593 22053 22599
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22624 22155 22627
rect 22204 22624 22232 22732
rect 22388 22692 22416 22732
rect 22462 22720 22468 22772
rect 22520 22760 22526 22772
rect 24210 22769 24216 22772
rect 24029 22763 24087 22769
rect 24029 22760 24041 22763
rect 22520 22732 24041 22760
rect 22520 22720 22526 22732
rect 24029 22729 24041 22732
rect 24075 22729 24087 22763
rect 24029 22723 24087 22729
rect 24197 22763 24216 22769
rect 24197 22729 24209 22763
rect 24268 22760 24274 22772
rect 25025 22763 25083 22769
rect 25025 22760 25037 22763
rect 24268 22732 25037 22760
rect 24197 22723 24216 22729
rect 24210 22720 24216 22723
rect 24268 22720 24274 22732
rect 25025 22729 25037 22732
rect 25071 22760 25083 22763
rect 25774 22760 25780 22772
rect 25071 22732 25452 22760
rect 25735 22732 25780 22760
rect 25071 22729 25083 22732
rect 25025 22723 25083 22729
rect 23106 22692 23112 22704
rect 22143 22596 22232 22624
rect 22278 22618 22284 22670
rect 22336 22633 22342 22670
rect 22388 22664 23112 22692
rect 23106 22652 23112 22664
rect 23164 22692 23170 22704
rect 23477 22695 23535 22701
rect 23477 22692 23489 22695
rect 23164 22664 23489 22692
rect 23164 22652 23170 22664
rect 23477 22661 23489 22664
rect 23523 22661 23535 22695
rect 23477 22655 23535 22661
rect 24302 22652 24308 22704
rect 24360 22692 24366 22704
rect 24397 22695 24455 22701
rect 24397 22692 24409 22695
rect 24360 22664 24409 22692
rect 24360 22652 24366 22664
rect 24397 22661 24409 22664
rect 24443 22661 24455 22695
rect 24397 22655 24455 22661
rect 25225 22695 25283 22701
rect 25225 22661 25237 22695
rect 25271 22661 25283 22695
rect 25424 22692 25452 22732
rect 25774 22720 25780 22732
rect 25832 22720 25838 22772
rect 26234 22720 26240 22772
rect 26292 22760 26298 22772
rect 26786 22760 26792 22772
rect 26292 22732 26792 22760
rect 26292 22720 26298 22732
rect 26786 22720 26792 22732
rect 26844 22720 26850 22772
rect 28166 22760 28172 22772
rect 28127 22732 28172 22760
rect 28166 22720 28172 22732
rect 28224 22720 28230 22772
rect 25498 22692 25504 22704
rect 25411 22664 25504 22692
rect 25225 22655 25283 22661
rect 22336 22618 22347 22633
rect 22143 22593 22155 22596
rect 22097 22587 22155 22593
rect 22289 22593 22301 22618
rect 22335 22593 22347 22618
rect 22289 22587 22347 22593
rect 22381 22627 22439 22633
rect 22381 22593 22393 22627
rect 22427 22624 22439 22627
rect 22830 22624 22836 22636
rect 22427 22596 22836 22624
rect 22427 22593 22439 22596
rect 22381 22587 22439 22593
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 23014 22584 23020 22636
rect 23072 22624 23078 22636
rect 23201 22627 23259 22633
rect 23072 22596 23117 22624
rect 23072 22584 23078 22596
rect 23201 22593 23213 22627
rect 23247 22593 23259 22627
rect 23566 22624 23572 22636
rect 23527 22596 23572 22624
rect 23201 22587 23259 22593
rect 22922 22556 22928 22568
rect 17552 22528 20383 22556
rect 21928 22528 22928 22556
rect 17552 22516 17558 22528
rect 15470 22448 15476 22500
rect 15528 22488 15534 22500
rect 20257 22491 20315 22497
rect 20257 22488 20269 22491
rect 15528 22460 20269 22488
rect 15528 22448 15534 22460
rect 20257 22457 20269 22460
rect 20303 22457 20315 22491
rect 20355 22488 20383 22528
rect 22922 22516 22928 22528
rect 22980 22516 22986 22568
rect 23216 22556 23244 22587
rect 23566 22584 23572 22596
rect 23624 22584 23630 22636
rect 23934 22584 23940 22636
rect 23992 22624 23998 22636
rect 25240 22624 25268 22655
rect 25498 22652 25504 22664
rect 25556 22692 25562 22704
rect 26694 22692 26700 22704
rect 25556 22664 26700 22692
rect 25556 22652 25562 22664
rect 26694 22652 26700 22664
rect 26752 22652 26758 22704
rect 23992 22596 25268 22624
rect 25961 22627 26019 22633
rect 23992 22584 23998 22596
rect 25961 22593 25973 22627
rect 26007 22624 26019 22627
rect 26878 22624 26884 22636
rect 26007 22596 26884 22624
rect 26007 22593 26019 22596
rect 25961 22587 26019 22593
rect 26878 22584 26884 22596
rect 26936 22584 26942 22636
rect 27709 22627 27767 22633
rect 27709 22593 27721 22627
rect 27755 22624 27767 22627
rect 27890 22624 27896 22636
rect 27755 22596 27896 22624
rect 27755 22593 27767 22596
rect 27709 22587 27767 22593
rect 27890 22584 27896 22596
rect 27948 22584 27954 22636
rect 28258 22584 28264 22636
rect 28316 22624 28322 22636
rect 28353 22627 28411 22633
rect 28353 22624 28365 22627
rect 28316 22596 28365 22624
rect 28316 22584 28322 22596
rect 28353 22593 28365 22596
rect 28399 22593 28411 22627
rect 28353 22587 28411 22593
rect 23842 22556 23848 22568
rect 23216 22528 23848 22556
rect 23842 22516 23848 22528
rect 23900 22516 23906 22568
rect 24946 22516 24952 22568
rect 25004 22556 25010 22568
rect 25590 22556 25596 22568
rect 25004 22528 25596 22556
rect 25004 22516 25010 22528
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 26605 22559 26663 22565
rect 26605 22525 26617 22559
rect 26651 22556 26663 22559
rect 28626 22556 28632 22568
rect 26651 22528 28632 22556
rect 26651 22525 26663 22528
rect 26605 22519 26663 22525
rect 28626 22516 28632 22528
rect 28684 22516 28690 22568
rect 24857 22491 24915 22497
rect 24857 22488 24869 22491
rect 20355 22460 24869 22488
rect 20257 22451 20315 22457
rect 24857 22457 24869 22460
rect 24903 22457 24915 22491
rect 24857 22451 24915 22457
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 17497 22423 17555 22429
rect 17497 22420 17509 22423
rect 16724 22392 17509 22420
rect 16724 22380 16730 22392
rect 17497 22389 17509 22392
rect 17543 22420 17555 22423
rect 20070 22420 20076 22432
rect 17543 22392 20076 22420
rect 17543 22389 17555 22392
rect 17497 22383 17555 22389
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 20438 22420 20444 22432
rect 20399 22392 20444 22420
rect 20438 22380 20444 22392
rect 20496 22380 20502 22432
rect 21269 22423 21327 22429
rect 21269 22389 21281 22423
rect 21315 22420 21327 22423
rect 21358 22420 21364 22432
rect 21315 22392 21364 22420
rect 21315 22389 21327 22392
rect 21269 22383 21327 22389
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 22278 22380 22284 22432
rect 22336 22420 22342 22432
rect 22557 22423 22615 22429
rect 22557 22420 22569 22423
rect 22336 22392 22569 22420
rect 22336 22380 22342 22392
rect 22557 22389 22569 22392
rect 22603 22389 22615 22423
rect 22557 22383 22615 22389
rect 24213 22423 24271 22429
rect 24213 22389 24225 22423
rect 24259 22420 24271 22423
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 24259 22392 25053 22420
rect 24259 22389 24271 22392
rect 24213 22383 24271 22389
rect 25041 22389 25053 22392
rect 25087 22420 25099 22423
rect 25774 22420 25780 22432
rect 25087 22392 25780 22420
rect 25087 22389 25099 22392
rect 25041 22383 25099 22389
rect 25774 22380 25780 22392
rect 25832 22420 25838 22432
rect 27154 22420 27160 22432
rect 25832 22392 27160 22420
rect 25832 22380 25838 22392
rect 27154 22380 27160 22392
rect 27212 22380 27218 22432
rect 27246 22380 27252 22432
rect 27304 22420 27310 22432
rect 29362 22420 29368 22432
rect 27304 22392 29368 22420
rect 27304 22380 27310 22392
rect 29362 22380 29368 22392
rect 29420 22380 29426 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 18877 22219 18935 22225
rect 18877 22185 18889 22219
rect 18923 22216 18935 22219
rect 20438 22216 20444 22228
rect 18923 22188 20444 22216
rect 18923 22185 18935 22188
rect 18877 22179 18935 22185
rect 20438 22176 20444 22188
rect 20496 22216 20502 22228
rect 22005 22219 22063 22225
rect 22005 22216 22017 22219
rect 20496 22188 22017 22216
rect 20496 22176 20502 22188
rect 22005 22185 22017 22188
rect 22051 22216 22063 22219
rect 22278 22216 22284 22228
rect 22051 22188 22284 22216
rect 22051 22185 22063 22188
rect 22005 22179 22063 22185
rect 22278 22176 22284 22188
rect 22336 22216 22342 22228
rect 22833 22219 22891 22225
rect 22833 22216 22845 22219
rect 22336 22188 22845 22216
rect 22336 22176 22342 22188
rect 22833 22185 22845 22188
rect 22879 22216 22891 22219
rect 22879 22188 22968 22216
rect 22879 22185 22891 22188
rect 22833 22179 22891 22185
rect 19705 22151 19763 22157
rect 19705 22117 19717 22151
rect 19751 22148 19763 22151
rect 19886 22148 19892 22160
rect 19751 22120 19892 22148
rect 19751 22117 19763 22120
rect 19705 22111 19763 22117
rect 19886 22108 19892 22120
rect 19944 22108 19950 22160
rect 19978 22108 19984 22160
rect 20036 22148 20042 22160
rect 20162 22148 20168 22160
rect 20036 22120 20168 22148
rect 20036 22108 20042 22120
rect 20162 22108 20168 22120
rect 20220 22108 20226 22160
rect 20254 22108 20260 22160
rect 20312 22148 20318 22160
rect 21085 22151 21143 22157
rect 21085 22148 21097 22151
rect 20312 22120 21097 22148
rect 20312 22108 20318 22120
rect 21085 22117 21097 22120
rect 21131 22148 21143 22151
rect 22940 22148 22968 22188
rect 23014 22176 23020 22228
rect 23072 22216 23078 22228
rect 23661 22219 23719 22225
rect 23661 22216 23673 22219
rect 23072 22188 23117 22216
rect 23166 22188 23673 22216
rect 23072 22176 23078 22188
rect 23166 22148 23194 22188
rect 23661 22185 23673 22188
rect 23707 22216 23719 22219
rect 24394 22216 24400 22228
rect 23707 22188 24400 22216
rect 23707 22185 23719 22188
rect 23661 22179 23719 22185
rect 24394 22176 24400 22188
rect 24452 22176 24458 22228
rect 25777 22219 25835 22225
rect 25777 22185 25789 22219
rect 25823 22216 25835 22219
rect 25866 22216 25872 22228
rect 25823 22188 25872 22216
rect 25823 22185 25835 22188
rect 25777 22179 25835 22185
rect 25866 22176 25872 22188
rect 25924 22176 25930 22228
rect 26142 22176 26148 22228
rect 26200 22216 26206 22228
rect 27065 22219 27123 22225
rect 27065 22216 27077 22219
rect 26200 22188 27077 22216
rect 26200 22176 26206 22188
rect 27065 22185 27077 22188
rect 27111 22185 27123 22219
rect 27065 22179 27123 22185
rect 27338 22176 27344 22228
rect 27396 22216 27402 22228
rect 27525 22219 27583 22225
rect 27525 22216 27537 22219
rect 27396 22188 27537 22216
rect 27396 22176 27402 22188
rect 27525 22185 27537 22188
rect 27571 22185 27583 22219
rect 27525 22179 27583 22185
rect 21131 22120 21486 22148
rect 22940 22120 23194 22148
rect 21131 22117 21143 22120
rect 21085 22111 21143 22117
rect 18325 22083 18383 22089
rect 18325 22049 18337 22083
rect 18371 22080 18383 22083
rect 19794 22080 19800 22092
rect 18371 22052 19800 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 19794 22040 19800 22052
rect 19852 22040 19858 22092
rect 19904 22080 19932 22108
rect 21358 22080 21364 22092
rect 19904 22052 21364 22080
rect 21358 22040 21364 22052
rect 21416 22040 21422 22092
rect 21458 22080 21486 22120
rect 23382 22108 23388 22160
rect 23440 22148 23446 22160
rect 23477 22151 23535 22157
rect 23477 22148 23489 22151
rect 23440 22120 23489 22148
rect 23440 22108 23446 22120
rect 23477 22117 23489 22120
rect 23523 22117 23535 22151
rect 23477 22111 23535 22117
rect 26421 22151 26479 22157
rect 26421 22117 26433 22151
rect 26467 22148 26479 22151
rect 28534 22148 28540 22160
rect 26467 22120 28540 22148
rect 26467 22117 26479 22120
rect 26421 22111 26479 22117
rect 28534 22108 28540 22120
rect 28592 22108 28598 22160
rect 24118 22080 24124 22092
rect 21458 22052 24124 22080
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 15930 21972 15936 22024
rect 15988 22012 15994 22024
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 15988 21984 17785 22012
rect 15988 21972 15994 21984
rect 17773 21981 17785 21984
rect 17819 22012 17831 22015
rect 20254 22012 20260 22024
rect 17819 21984 20260 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 21266 22012 21272 22024
rect 21227 21984 21272 22012
rect 21266 21972 21272 21984
rect 21324 21972 21330 22024
rect 24765 22015 24823 22021
rect 22004 21984 22784 22012
rect 17402 21904 17408 21956
rect 17460 21944 17466 21956
rect 17460 21916 19748 21944
rect 17460 21904 17466 21916
rect 19720 21876 19748 21916
rect 20806 21904 20812 21956
rect 20864 21944 20870 21956
rect 22004 21953 22032 21984
rect 21989 21947 22047 21953
rect 21989 21944 22001 21947
rect 20864 21916 22001 21944
rect 20864 21904 20870 21916
rect 21989 21913 22001 21916
rect 22035 21913 22047 21947
rect 21989 21907 22047 21913
rect 22189 21947 22247 21953
rect 22189 21913 22201 21947
rect 22235 21944 22247 21947
rect 22462 21944 22468 21956
rect 22235 21916 22468 21944
rect 22235 21913 22247 21916
rect 22189 21907 22247 21913
rect 22462 21904 22468 21916
rect 22520 21904 22526 21956
rect 22646 21944 22652 21956
rect 22607 21916 22652 21944
rect 22646 21904 22652 21916
rect 22704 21904 22710 21956
rect 22756 21944 22784 21984
rect 24765 21981 24777 22015
rect 24811 22012 24823 22015
rect 27338 22012 27344 22024
rect 24811 21984 27344 22012
rect 24811 21981 24823 21984
rect 24765 21975 24823 21981
rect 27338 21972 27344 21984
rect 27396 21972 27402 22024
rect 27522 21972 27528 22024
rect 27580 22012 27586 22024
rect 27706 22012 27712 22024
rect 27580 21984 27712 22012
rect 27580 21972 27586 21984
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 28350 22012 28356 22024
rect 28311 21984 28356 22012
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 22756 21916 22876 21944
rect 21821 21879 21879 21885
rect 21821 21876 21833 21879
rect 19720 21848 21833 21876
rect 21821 21845 21833 21848
rect 21867 21845 21879 21879
rect 21821 21839 21879 21845
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 22738 21876 22744 21888
rect 22428 21848 22744 21876
rect 22428 21836 22434 21848
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 22848 21885 22876 21916
rect 23014 21904 23020 21956
rect 23072 21944 23078 21956
rect 23845 21947 23903 21953
rect 23845 21944 23857 21947
rect 23072 21916 23857 21944
rect 23072 21904 23078 21916
rect 23845 21913 23857 21916
rect 23891 21913 23903 21947
rect 23845 21907 23903 21913
rect 22848 21879 22917 21885
rect 22848 21848 22871 21879
rect 22859 21845 22871 21848
rect 22905 21876 22917 21879
rect 23382 21876 23388 21888
rect 22905 21848 23388 21876
rect 22905 21845 22917 21848
rect 22859 21839 22917 21845
rect 23382 21836 23388 21848
rect 23440 21876 23446 21888
rect 23635 21879 23693 21885
rect 23635 21876 23647 21879
rect 23440 21848 23647 21876
rect 23440 21836 23446 21848
rect 23635 21845 23647 21848
rect 23681 21876 23693 21879
rect 24486 21876 24492 21888
rect 23681 21848 24492 21876
rect 23681 21845 23693 21848
rect 23635 21839 23693 21845
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 24670 21876 24676 21888
rect 24631 21848 24676 21876
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 19337 21675 19395 21681
rect 19337 21641 19349 21675
rect 19383 21672 19395 21675
rect 19426 21672 19432 21684
rect 19383 21644 19432 21672
rect 19383 21641 19395 21644
rect 19337 21635 19395 21641
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 21450 21632 21456 21684
rect 21508 21672 21514 21684
rect 22097 21675 22155 21681
rect 22097 21672 22109 21675
rect 21508 21644 22109 21672
rect 21508 21632 21514 21644
rect 22097 21641 22109 21644
rect 22143 21641 22155 21675
rect 22097 21635 22155 21641
rect 23845 21675 23903 21681
rect 23845 21641 23857 21675
rect 23891 21672 23903 21675
rect 24394 21672 24400 21684
rect 23891 21644 24400 21672
rect 23891 21641 23903 21644
rect 23845 21635 23903 21641
rect 24394 21632 24400 21644
rect 24452 21632 24458 21684
rect 25958 21632 25964 21684
rect 26016 21672 26022 21684
rect 26421 21675 26479 21681
rect 26421 21672 26433 21675
rect 26016 21644 26433 21672
rect 26016 21632 26022 21644
rect 26421 21641 26433 21644
rect 26467 21641 26479 21675
rect 26421 21635 26479 21641
rect 18690 21564 18696 21616
rect 18748 21604 18754 21616
rect 21174 21604 21180 21616
rect 18748 21576 21180 21604
rect 18748 21564 18754 21576
rect 21174 21564 21180 21576
rect 21232 21564 21238 21616
rect 21266 21564 21272 21616
rect 21324 21604 21330 21616
rect 22249 21607 22307 21613
rect 22249 21604 22261 21607
rect 21324 21576 22261 21604
rect 21324 21564 21330 21576
rect 22249 21573 22261 21576
rect 22295 21573 22307 21607
rect 22462 21604 22468 21616
rect 22423 21576 22468 21604
rect 22249 21567 22307 21573
rect 22462 21564 22468 21576
rect 22520 21564 22526 21616
rect 23290 21604 23296 21616
rect 23063 21573 23121 21579
rect 23251 21576 23296 21604
rect 23063 21539 23075 21573
rect 23109 21570 23121 21573
rect 23109 21539 23136 21570
rect 23290 21564 23296 21576
rect 23348 21564 23354 21616
rect 23400 21576 23888 21604
rect 23063 21536 23136 21539
rect 23400 21536 23428 21576
rect 23750 21536 23756 21548
rect 23063 21533 23428 21536
rect 23108 21508 23428 21533
rect 23711 21508 23756 21536
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 1578 21468 1584 21480
rect 1539 21440 1584 21468
rect 1578 21428 1584 21440
rect 1636 21428 1642 21480
rect 12342 21428 12348 21480
rect 12400 21468 12406 21480
rect 23860 21468 23888 21576
rect 24486 21564 24492 21616
rect 24544 21604 24550 21616
rect 25130 21604 25136 21616
rect 24544 21576 25136 21604
rect 24544 21564 24550 21576
rect 25130 21564 25136 21576
rect 25188 21604 25194 21616
rect 25685 21607 25743 21613
rect 25685 21604 25697 21607
rect 25188 21576 25697 21604
rect 25188 21564 25194 21576
rect 25685 21573 25697 21576
rect 25731 21604 25743 21607
rect 26142 21604 26148 21616
rect 25731 21576 26148 21604
rect 25731 21573 25743 21576
rect 25685 21567 25743 21573
rect 26142 21564 26148 21576
rect 26200 21604 26206 21616
rect 26326 21604 26332 21616
rect 26200 21576 26332 21604
rect 26200 21564 26206 21576
rect 26326 21564 26332 21576
rect 26384 21564 26390 21616
rect 27246 21604 27252 21616
rect 26620 21576 27252 21604
rect 24026 21496 24032 21548
rect 24084 21536 24090 21548
rect 26620 21545 26648 21576
rect 27246 21564 27252 21576
rect 27304 21564 27310 21616
rect 24397 21539 24455 21545
rect 24397 21536 24409 21539
rect 24084 21508 24409 21536
rect 24084 21496 24090 21508
rect 24397 21505 24409 21508
rect 24443 21505 24455 21539
rect 24397 21499 24455 21505
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21505 26663 21539
rect 26605 21499 26663 21505
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21536 27215 21539
rect 28074 21536 28080 21548
rect 27203 21508 28080 21536
rect 27203 21505 27215 21508
rect 27157 21499 27215 21505
rect 28074 21496 28080 21508
rect 28132 21496 28138 21548
rect 24210 21468 24216 21480
rect 12400 21440 22324 21468
rect 23860 21440 24216 21468
rect 12400 21428 12406 21440
rect 19058 21360 19064 21412
rect 19116 21400 19122 21412
rect 19797 21403 19855 21409
rect 19797 21400 19809 21403
rect 19116 21372 19809 21400
rect 19116 21360 19122 21372
rect 19797 21369 19809 21372
rect 19843 21369 19855 21403
rect 19797 21363 19855 21369
rect 18782 21332 18788 21344
rect 18743 21304 18788 21332
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 19812 21332 19840 21363
rect 20438 21360 20444 21412
rect 20496 21400 20502 21412
rect 20717 21403 20775 21409
rect 20717 21400 20729 21403
rect 20496 21372 20729 21400
rect 20496 21360 20502 21372
rect 20717 21369 20729 21372
rect 20763 21369 20775 21403
rect 22296 21400 22324 21440
rect 24210 21428 24216 21440
rect 24268 21428 24274 21480
rect 22296 21372 23152 21400
rect 20717 21363 20775 21369
rect 23124 21344 23152 21372
rect 20898 21332 20904 21344
rect 19812 21304 20904 21332
rect 20898 21292 20904 21304
rect 20956 21332 20962 21344
rect 21358 21332 21364 21344
rect 20956 21304 21364 21332
rect 20956 21292 20962 21304
rect 21358 21292 21364 21304
rect 21416 21292 21422 21344
rect 21450 21292 21456 21344
rect 21508 21332 21514 21344
rect 22281 21335 22339 21341
rect 22281 21332 22293 21335
rect 21508 21304 22293 21332
rect 21508 21292 21514 21304
rect 22281 21301 22293 21304
rect 22327 21332 22339 21335
rect 22370 21332 22376 21344
rect 22327 21304 22376 21332
rect 22327 21301 22339 21304
rect 22281 21295 22339 21301
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 22646 21292 22652 21344
rect 22704 21332 22710 21344
rect 22925 21335 22983 21341
rect 22925 21332 22937 21335
rect 22704 21304 22937 21332
rect 22704 21292 22710 21304
rect 22925 21301 22937 21304
rect 22971 21301 22983 21335
rect 23106 21332 23112 21344
rect 23067 21304 23112 21332
rect 22925 21295 22983 21301
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 28350 21332 28356 21344
rect 28311 21304 28356 21332
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 19889 21131 19947 21137
rect 19889 21097 19901 21131
rect 19935 21128 19947 21131
rect 20346 21128 20352 21140
rect 19935 21100 20352 21128
rect 19935 21097 19947 21100
rect 19889 21091 19947 21097
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 20438 21088 20444 21140
rect 20496 21128 20502 21140
rect 20496 21100 20541 21128
rect 20496 21088 20502 21100
rect 20806 21088 20812 21140
rect 20864 21128 20870 21140
rect 20901 21131 20959 21137
rect 20901 21128 20913 21131
rect 20864 21100 20913 21128
rect 20864 21088 20870 21100
rect 20901 21097 20913 21100
rect 20947 21097 20959 21131
rect 20901 21091 20959 21097
rect 21358 21088 21364 21140
rect 21416 21128 21422 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 21416 21100 21465 21128
rect 21416 21088 21422 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 21453 21091 21511 21097
rect 23109 21131 23167 21137
rect 23109 21097 23121 21131
rect 23155 21128 23167 21131
rect 24854 21128 24860 21140
rect 23155 21100 24860 21128
rect 23155 21097 23167 21100
rect 23109 21091 23167 21097
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 25130 21128 25136 21140
rect 25091 21100 25136 21128
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 25774 21128 25780 21140
rect 25735 21100 25780 21128
rect 25774 21088 25780 21100
rect 25832 21128 25838 21140
rect 26237 21131 26295 21137
rect 26237 21128 26249 21131
rect 25832 21100 26249 21128
rect 25832 21088 25838 21100
rect 26237 21097 26249 21100
rect 26283 21128 26295 21131
rect 26326 21128 26332 21140
rect 26283 21100 26332 21128
rect 26283 21097 26295 21100
rect 26237 21091 26295 21097
rect 26326 21088 26332 21100
rect 26384 21088 26390 21140
rect 28353 21131 28411 21137
rect 28353 21097 28365 21131
rect 28399 21128 28411 21131
rect 29178 21128 29184 21140
rect 28399 21100 29184 21128
rect 28399 21097 28411 21100
rect 28353 21091 28411 21097
rect 29178 21088 29184 21100
rect 29236 21088 29242 21140
rect 18782 21020 18788 21072
rect 18840 21060 18846 21072
rect 19518 21060 19524 21072
rect 18840 21032 19524 21060
rect 18840 21020 18846 21032
rect 19518 21020 19524 21032
rect 19576 21060 19582 21072
rect 21082 21060 21088 21072
rect 19576 21032 21088 21060
rect 19576 21020 19582 21032
rect 21082 21020 21088 21032
rect 21140 21020 21146 21072
rect 22370 21020 22376 21072
rect 22428 21060 22434 21072
rect 23750 21060 23756 21072
rect 22428 21032 23756 21060
rect 22428 21020 22434 21032
rect 23750 21020 23756 21032
rect 23808 21020 23814 21072
rect 24210 21020 24216 21072
rect 24268 21060 24274 21072
rect 24581 21063 24639 21069
rect 24581 21060 24593 21063
rect 24268 21032 24593 21060
rect 24268 21020 24274 21032
rect 24581 21029 24593 21032
rect 24627 21060 24639 21063
rect 24762 21060 24768 21072
rect 24627 21032 24768 21060
rect 24627 21029 24639 21032
rect 24581 21023 24639 21029
rect 24762 21020 24768 21032
rect 24820 21020 24826 21072
rect 24670 20992 24676 21004
rect 22066 20964 24676 20992
rect 20530 20884 20536 20936
rect 20588 20924 20594 20936
rect 22066 20924 22094 20964
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 24854 20952 24860 21004
rect 24912 20992 24918 21004
rect 25792 20992 25820 21088
rect 27709 21063 27767 21069
rect 27709 21029 27721 21063
rect 27755 21060 27767 21063
rect 28442 21060 28448 21072
rect 27755 21032 28448 21060
rect 27755 21029 27767 21032
rect 27709 21023 27767 21029
rect 28442 21020 28448 21032
rect 28500 21020 28506 21072
rect 24912 20964 25820 20992
rect 27065 20995 27123 21001
rect 24912 20952 24918 20964
rect 27065 20961 27077 20995
rect 27111 20992 27123 20995
rect 29270 20992 29276 21004
rect 27111 20964 29276 20992
rect 27111 20961 27123 20964
rect 27065 20955 27123 20961
rect 29270 20952 29276 20964
rect 29328 20952 29334 21004
rect 20588 20896 22094 20924
rect 22373 20927 22431 20933
rect 20588 20884 20594 20896
rect 22373 20893 22385 20927
rect 22419 20924 22431 20927
rect 22646 20924 22652 20936
rect 22419 20896 22652 20924
rect 22419 20893 22431 20896
rect 22373 20887 22431 20893
rect 22646 20884 22652 20896
rect 22704 20924 22710 20936
rect 23014 20924 23020 20936
rect 22704 20896 23020 20924
rect 22704 20884 22710 20896
rect 23014 20884 23020 20896
rect 23072 20884 23078 20936
rect 23201 20927 23259 20933
rect 23201 20893 23213 20927
rect 23247 20924 23259 20927
rect 24578 20924 24584 20936
rect 23247 20896 24584 20924
rect 23247 20893 23259 20896
rect 23201 20887 23259 20893
rect 24578 20884 24584 20896
rect 24636 20884 24642 20936
rect 22554 20856 22560 20868
rect 22515 20828 22560 20856
rect 22554 20816 22560 20828
rect 22612 20816 22618 20868
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 19978 20584 19984 20596
rect 19939 20556 19984 20584
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 20990 20584 20996 20596
rect 20951 20556 20996 20584
rect 20990 20544 20996 20556
rect 21048 20544 21054 20596
rect 22097 20587 22155 20593
rect 22097 20553 22109 20587
rect 22143 20584 22155 20587
rect 22462 20584 22468 20596
rect 22143 20556 22468 20584
rect 22143 20553 22155 20556
rect 22097 20547 22155 20553
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 22646 20584 22652 20596
rect 22607 20556 22652 20584
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 23201 20587 23259 20593
rect 23201 20584 23213 20587
rect 22980 20556 23213 20584
rect 22980 20544 22986 20556
rect 23201 20553 23213 20556
rect 23247 20553 23259 20587
rect 23201 20547 23259 20553
rect 24762 20544 24768 20596
rect 24820 20584 24826 20596
rect 26053 20587 26111 20593
rect 24820 20556 24992 20584
rect 24820 20544 24826 20556
rect 20254 20476 20260 20528
rect 20312 20516 20318 20528
rect 22370 20516 22376 20528
rect 20312 20488 22376 20516
rect 20312 20476 20318 20488
rect 22370 20476 22376 20488
rect 22428 20476 22434 20528
rect 23106 20476 23112 20528
rect 23164 20516 23170 20528
rect 23845 20519 23903 20525
rect 23845 20516 23857 20519
rect 23164 20488 23857 20516
rect 23164 20476 23170 20488
rect 23845 20485 23857 20488
rect 23891 20516 23903 20519
rect 24854 20516 24860 20528
rect 23891 20488 24860 20516
rect 23891 20485 23903 20488
rect 23845 20479 23903 20485
rect 24854 20476 24860 20488
rect 24912 20476 24918 20528
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 20128 20420 20545 20448
rect 20128 20408 20134 20420
rect 20533 20417 20545 20420
rect 20579 20448 20591 20451
rect 22830 20448 22836 20460
rect 20579 20420 22836 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 22830 20408 22836 20420
rect 22888 20448 22894 20460
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 22888 20420 24317 20448
rect 22888 20408 22894 20420
rect 24305 20417 24317 20420
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 24964 20253 24992 20556
rect 26053 20553 26065 20587
rect 26099 20584 26111 20587
rect 26418 20584 26424 20596
rect 26099 20556 26424 20584
rect 26099 20553 26111 20556
rect 26053 20547 26111 20553
rect 26418 20544 26424 20556
rect 26476 20544 26482 20596
rect 27246 20584 27252 20596
rect 27207 20556 27252 20584
rect 27246 20544 27252 20556
rect 27304 20544 27310 20596
rect 28169 20587 28227 20593
rect 28169 20553 28181 20587
rect 28215 20584 28227 20587
rect 29454 20584 29460 20596
rect 28215 20556 29460 20584
rect 28215 20553 28227 20556
rect 28169 20547 28227 20553
rect 29454 20544 29460 20556
rect 29512 20544 29518 20596
rect 28350 20448 28356 20460
rect 28311 20420 28356 20448
rect 28350 20408 28356 20420
rect 28408 20408 28414 20460
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20244 25007 20247
rect 25501 20247 25559 20253
rect 25501 20244 25513 20247
rect 24995 20216 25513 20244
rect 24995 20213 25007 20216
rect 24949 20207 25007 20213
rect 25501 20213 25513 20216
rect 25547 20244 25559 20247
rect 25958 20244 25964 20256
rect 25547 20216 25964 20244
rect 25547 20213 25559 20216
rect 25501 20207 25559 20213
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 26326 20204 26332 20256
rect 26384 20244 26390 20256
rect 26605 20247 26663 20253
rect 26605 20244 26617 20247
rect 26384 20216 26617 20244
rect 26384 20204 26390 20216
rect 26605 20213 26617 20216
rect 26651 20244 26663 20247
rect 26970 20244 26976 20256
rect 26651 20216 26976 20244
rect 26651 20213 26663 20216
rect 26605 20207 26663 20213
rect 26970 20204 26976 20216
rect 27028 20204 27034 20256
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 20622 20040 20628 20052
rect 20583 20012 20628 20040
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 21634 20040 21640 20052
rect 21595 20012 21640 20040
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 22278 20040 22284 20052
rect 22239 20012 22284 20040
rect 22278 20000 22284 20012
rect 22336 20040 22342 20052
rect 23109 20043 23167 20049
rect 23109 20040 23121 20043
rect 22336 20012 23121 20040
rect 22336 20000 22342 20012
rect 23109 20009 23121 20012
rect 23155 20040 23167 20043
rect 23661 20043 23719 20049
rect 23661 20040 23673 20043
rect 23155 20012 23673 20040
rect 23155 20009 23167 20012
rect 23109 20003 23167 20009
rect 23661 20009 23673 20012
rect 23707 20040 23719 20043
rect 23750 20040 23756 20052
rect 23707 20012 23756 20040
rect 23707 20009 23719 20012
rect 23661 20003 23719 20009
rect 23750 20000 23756 20012
rect 23808 20000 23814 20052
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 25133 20043 25191 20049
rect 25133 20040 25145 20043
rect 24176 20012 25145 20040
rect 24176 20000 24182 20012
rect 25133 20009 25145 20012
rect 25179 20009 25191 20043
rect 25133 20003 25191 20009
rect 27157 20043 27215 20049
rect 27157 20009 27169 20043
rect 27203 20040 27215 20043
rect 27522 20040 27528 20052
rect 27203 20012 27528 20040
rect 27203 20009 27215 20012
rect 27157 20003 27215 20009
rect 27522 20000 27528 20012
rect 27580 20000 27586 20052
rect 27709 20043 27767 20049
rect 27709 20009 27721 20043
rect 27755 20040 27767 20043
rect 28350 20040 28356 20052
rect 27755 20012 28356 20040
rect 27755 20009 27767 20012
rect 27709 20003 27767 20009
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 20640 19972 20668 20000
rect 24581 19975 24639 19981
rect 24581 19972 24593 19975
rect 20640 19944 24593 19972
rect 24581 19941 24593 19944
rect 24627 19972 24639 19975
rect 25774 19972 25780 19984
rect 24627 19944 25780 19972
rect 24627 19941 24639 19944
rect 24581 19935 24639 19941
rect 25774 19932 25780 19944
rect 25832 19932 25838 19984
rect 21177 19907 21235 19913
rect 21177 19873 21189 19907
rect 21223 19904 21235 19907
rect 22646 19904 22652 19916
rect 21223 19876 22652 19904
rect 21223 19873 21235 19876
rect 21177 19867 21235 19873
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 28350 19836 28356 19848
rect 28311 19808 28356 19836
rect 28350 19796 28356 19808
rect 28408 19796 28414 19848
rect 25777 19703 25835 19709
rect 25777 19669 25789 19703
rect 25823 19700 25835 19703
rect 25958 19700 25964 19712
rect 25823 19672 25964 19700
rect 25823 19669 25835 19672
rect 25777 19663 25835 19669
rect 25958 19660 25964 19672
rect 26016 19660 26022 19712
rect 26234 19660 26240 19712
rect 26292 19700 26298 19712
rect 26329 19703 26387 19709
rect 26329 19700 26341 19703
rect 26292 19672 26341 19700
rect 26292 19660 26298 19672
rect 26329 19669 26341 19672
rect 26375 19700 26387 19703
rect 27154 19700 27160 19712
rect 26375 19672 27160 19700
rect 26375 19669 26387 19672
rect 26329 19663 26387 19669
rect 27154 19660 27160 19672
rect 27212 19660 27218 19712
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 21634 19456 21640 19508
rect 21692 19496 21698 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21692 19468 22017 19496
rect 21692 19456 21698 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22020 19224 22048 19459
rect 22646 19456 22652 19508
rect 22704 19496 22710 19508
rect 22833 19499 22891 19505
rect 22833 19496 22845 19499
rect 22704 19468 22845 19496
rect 22704 19456 22710 19468
rect 22833 19465 22845 19468
rect 22879 19465 22891 19499
rect 22833 19459 22891 19465
rect 23477 19499 23535 19505
rect 23477 19465 23489 19499
rect 23523 19496 23535 19499
rect 23658 19496 23664 19508
rect 23523 19468 23664 19496
rect 23523 19465 23535 19468
rect 23477 19459 23535 19465
rect 23658 19456 23664 19468
rect 23716 19456 23722 19508
rect 26142 19496 26148 19508
rect 26103 19468 26148 19496
rect 26142 19456 26148 19468
rect 26200 19456 26206 19508
rect 27709 19499 27767 19505
rect 27709 19465 27721 19499
rect 27755 19496 27767 19499
rect 28258 19496 28264 19508
rect 27755 19468 28264 19496
rect 27755 19465 27767 19468
rect 27709 19459 27767 19465
rect 28258 19456 28264 19468
rect 28316 19456 28322 19508
rect 25133 19431 25191 19437
rect 25133 19428 25145 19431
rect 24826 19400 25145 19428
rect 24029 19295 24087 19301
rect 24029 19261 24041 19295
rect 24075 19292 24087 19295
rect 24826 19292 24854 19400
rect 25133 19397 25145 19400
rect 25179 19428 25191 19431
rect 26050 19428 26056 19440
rect 25179 19400 26056 19428
rect 25179 19397 25191 19400
rect 25133 19391 25191 19397
rect 26050 19388 26056 19400
rect 26108 19388 26114 19440
rect 24075 19264 24854 19292
rect 24075 19261 24087 19264
rect 24029 19255 24087 19261
rect 24581 19227 24639 19233
rect 24581 19224 24593 19227
rect 22020 19196 24593 19224
rect 24581 19193 24593 19196
rect 24627 19224 24639 19227
rect 24854 19224 24860 19236
rect 24627 19196 24860 19224
rect 24627 19193 24639 19196
rect 24581 19187 24639 19193
rect 24854 19184 24860 19196
rect 24912 19184 24918 19236
rect 28350 19156 28356 19168
rect 28311 19128 28356 19156
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 23566 18952 23572 18964
rect 23527 18924 23572 18952
rect 23566 18912 23572 18924
rect 23624 18912 23630 18964
rect 24857 18955 24915 18961
rect 24857 18921 24869 18955
rect 24903 18952 24915 18955
rect 24946 18952 24952 18964
rect 24903 18924 24952 18952
rect 24903 18921 24915 18924
rect 24857 18915 24915 18921
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 23750 18844 23756 18896
rect 23808 18884 23814 18896
rect 26237 18887 26295 18893
rect 26237 18884 26249 18887
rect 23808 18856 26249 18884
rect 23808 18844 23814 18856
rect 26237 18853 26249 18856
rect 26283 18853 26295 18887
rect 26237 18847 26295 18853
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 28077 18819 28135 18825
rect 28077 18816 28089 18819
rect 23624 18788 28089 18816
rect 23624 18776 23630 18788
rect 28077 18785 28089 18788
rect 28123 18785 28135 18819
rect 28077 18779 28135 18785
rect 28350 18748 28356 18760
rect 28311 18720 28356 18748
rect 28350 18708 28356 18720
rect 28408 18708 28414 18760
rect 22370 18612 22376 18624
rect 22331 18584 22376 18612
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 22462 18572 22468 18624
rect 22520 18612 22526 18624
rect 23017 18615 23075 18621
rect 23017 18612 23029 18615
rect 22520 18584 23029 18612
rect 22520 18572 22526 18584
rect 23017 18581 23029 18584
rect 23063 18612 23075 18615
rect 25409 18615 25467 18621
rect 25409 18612 25421 18615
rect 23063 18584 25421 18612
rect 23063 18581 23075 18584
rect 23017 18575 23075 18581
rect 25409 18581 25421 18584
rect 25455 18612 25467 18615
rect 25682 18612 25688 18624
rect 25455 18584 25688 18612
rect 25455 18581 25467 18584
rect 25409 18575 25467 18581
rect 25682 18572 25688 18584
rect 25740 18572 25746 18624
rect 26878 18612 26884 18624
rect 26839 18584 26884 18612
rect 26878 18572 26884 18584
rect 26936 18572 26942 18624
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 25038 18408 25044 18420
rect 23716 18380 25044 18408
rect 23716 18368 23722 18380
rect 25038 18368 25044 18380
rect 25096 18408 25102 18420
rect 25869 18411 25927 18417
rect 25869 18408 25881 18411
rect 25096 18380 25881 18408
rect 25096 18368 25102 18380
rect 25869 18377 25881 18380
rect 25915 18377 25927 18411
rect 26510 18408 26516 18420
rect 26471 18380 26516 18408
rect 25869 18371 25927 18377
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 27614 18368 27620 18420
rect 27672 18408 27678 18420
rect 27709 18411 27767 18417
rect 27709 18408 27721 18411
rect 27672 18380 27721 18408
rect 27672 18368 27678 18380
rect 27709 18377 27721 18380
rect 27755 18377 27767 18411
rect 27709 18371 27767 18377
rect 21082 18300 21088 18352
rect 21140 18340 21146 18352
rect 23753 18343 23811 18349
rect 23753 18340 23765 18343
rect 21140 18312 23765 18340
rect 21140 18300 21146 18312
rect 23753 18309 23765 18312
rect 23799 18309 23811 18343
rect 23753 18303 23811 18309
rect 25958 18300 25964 18352
rect 26016 18340 26022 18352
rect 27157 18343 27215 18349
rect 27157 18340 27169 18343
rect 26016 18312 27169 18340
rect 26016 18300 26022 18312
rect 27157 18309 27169 18312
rect 27203 18309 27215 18343
rect 28350 18340 28356 18352
rect 28311 18312 28356 18340
rect 27157 18303 27215 18309
rect 28350 18300 28356 18312
rect 28408 18300 28414 18352
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 24854 18028 24860 18080
rect 24912 18068 24918 18080
rect 25409 18071 25467 18077
rect 24912 18040 24957 18068
rect 24912 18028 24918 18040
rect 25409 18037 25421 18071
rect 25455 18068 25467 18071
rect 25682 18068 25688 18080
rect 25455 18040 25688 18068
rect 25455 18037 25467 18040
rect 25409 18031 25467 18037
rect 25682 18028 25688 18040
rect 25740 18028 25746 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 22738 17824 22744 17876
rect 22796 17864 22802 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 22796 17836 24593 17864
rect 22796 17824 22802 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 25590 17864 25596 17876
rect 25551 17836 25596 17864
rect 24581 17827 24639 17833
rect 24596 17796 24624 17827
rect 25590 17824 25596 17836
rect 25648 17824 25654 17876
rect 25774 17824 25780 17876
rect 25832 17864 25838 17876
rect 26237 17867 26295 17873
rect 26237 17864 26249 17867
rect 25832 17836 26249 17864
rect 25832 17824 25838 17836
rect 26237 17833 26249 17836
rect 26283 17833 26295 17867
rect 26970 17864 26976 17876
rect 26931 17836 26976 17864
rect 26237 17827 26295 17833
rect 26970 17824 26976 17836
rect 27028 17824 27034 17876
rect 27709 17867 27767 17873
rect 27709 17833 27721 17867
rect 27755 17864 27767 17867
rect 27798 17864 27804 17876
rect 27755 17836 27804 17864
rect 27755 17833 27767 17836
rect 27709 17827 27767 17833
rect 27798 17824 27804 17836
rect 27856 17824 27862 17876
rect 25498 17796 25504 17808
rect 24596 17768 25504 17796
rect 25498 17756 25504 17768
rect 25556 17756 25562 17808
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 28350 17660 28356 17672
rect 28311 17632 28356 17660
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 25038 17320 25044 17332
rect 24999 17292 25044 17320
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 25498 17320 25504 17332
rect 25459 17292 25504 17320
rect 25498 17280 25504 17292
rect 25556 17280 25562 17332
rect 27154 17320 27160 17332
rect 27115 17292 27160 17320
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 23566 17212 23572 17264
rect 23624 17252 23630 17264
rect 26053 17255 26111 17261
rect 26053 17252 26065 17255
rect 23624 17224 26065 17252
rect 23624 17212 23630 17224
rect 26053 17221 26065 17224
rect 26099 17221 26111 17255
rect 26053 17215 26111 17221
rect 28350 16980 28356 16992
rect 28311 16952 28356 16980
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 26237 16779 26295 16785
rect 26237 16776 26249 16779
rect 24912 16748 26249 16776
rect 24912 16736 24918 16748
rect 26237 16745 26249 16748
rect 26283 16745 26295 16779
rect 26237 16739 26295 16745
rect 26878 16736 26884 16788
rect 26936 16776 26942 16788
rect 27801 16779 27859 16785
rect 27801 16776 27813 16779
rect 26936 16748 27813 16776
rect 26936 16736 26942 16748
rect 27801 16745 27813 16748
rect 27847 16745 27859 16779
rect 27801 16739 27859 16745
rect 25682 16668 25688 16720
rect 25740 16708 25746 16720
rect 26973 16711 27031 16717
rect 26973 16708 26985 16711
rect 25740 16680 26985 16708
rect 25740 16668 25746 16680
rect 26973 16677 26985 16680
rect 27019 16677 27031 16711
rect 26973 16671 27031 16677
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 22370 16192 22376 16244
rect 22428 16232 22434 16244
rect 27617 16235 27675 16241
rect 27617 16232 27629 16235
rect 22428 16204 27629 16232
rect 22428 16192 22434 16204
rect 27617 16201 27629 16204
rect 27663 16201 27675 16235
rect 27617 16195 27675 16201
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 28350 15892 28356 15904
rect 28311 15864 28356 15892
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 28350 14872 28356 14884
rect 28311 14844 28356 14872
rect 28350 14832 28356 14844
rect 28408 14832 28414 14884
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 28350 13716 28356 13728
rect 28311 13688 28356 13716
rect 28350 13676 28356 13688
rect 28408 13676 28414 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 28350 13308 28356 13320
rect 28311 13280 28356 13308
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 28350 11540 28356 11552
rect 28311 11512 28356 11540
rect 28350 11500 28356 11512
rect 28408 11500 28414 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 28350 11132 28356 11144
rect 28311 11104 28356 11132
rect 28350 11092 28356 11104
rect 28408 11092 28414 11144
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 28350 9432 28356 9444
rect 28311 9404 28356 9432
rect 28350 9392 28356 9404
rect 28408 9392 28414 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 28350 9092 28356 9104
rect 28311 9064 28356 9092
rect 28350 9052 28356 9064
rect 28408 9052 28414 9104
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 28350 7868 28356 7880
rect 28311 7840 28356 7868
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 28350 6780 28356 6792
rect 28311 6752 28356 6780
rect 28350 6740 28356 6752
rect 28408 6740 28414 6792
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 28350 5692 28356 5704
rect 28311 5664 28356 5692
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 28350 5012 28356 5024
rect 28311 4984 28356 5012
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 28350 3652 28356 3664
rect 28311 3624 28356 3652
rect 28350 3612 28356 3624
rect 28408 3612 28414 3664
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 28350 2836 28356 2848
rect 28311 2808 28356 2836
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
<< via1 >>
rect 11796 32172 11848 32224
rect 14924 32172 14976 32224
rect 20260 32036 20312 32088
rect 21548 32036 21600 32088
rect 8392 31900 8444 31952
rect 26884 31900 26936 31952
rect 14004 31832 14056 31884
rect 18696 31832 18748 31884
rect 11704 31764 11756 31816
rect 8576 31696 8628 31748
rect 13820 31696 13872 31748
rect 16580 31696 16632 31748
rect 18788 31696 18840 31748
rect 13728 31628 13780 31680
rect 18512 31628 18564 31680
rect 19984 31696 20036 31748
rect 21640 31696 21692 31748
rect 22652 31628 22704 31680
rect 22744 31628 22796 31680
rect 28356 31628 28408 31680
rect 7896 31526 7948 31578
rect 7960 31526 8012 31578
rect 8024 31526 8076 31578
rect 8088 31526 8140 31578
rect 8152 31526 8204 31578
rect 14842 31526 14894 31578
rect 14906 31526 14958 31578
rect 14970 31526 15022 31578
rect 15034 31526 15086 31578
rect 15098 31526 15150 31578
rect 21788 31526 21840 31578
rect 21852 31526 21904 31578
rect 21916 31526 21968 31578
rect 21980 31526 22032 31578
rect 22044 31526 22096 31578
rect 28734 31526 28786 31578
rect 28798 31526 28850 31578
rect 28862 31526 28914 31578
rect 28926 31526 28978 31578
rect 28990 31526 29042 31578
rect 1676 31424 1728 31476
rect 4988 31424 5040 31476
rect 8300 31424 8352 31476
rect 11612 31424 11664 31476
rect 11796 31467 11848 31476
rect 11796 31433 11805 31467
rect 11805 31433 11839 31467
rect 11839 31433 11848 31467
rect 11796 31424 11848 31433
rect 8484 31356 8536 31408
rect 9864 31356 9916 31408
rect 3884 31288 3936 31340
rect 5356 31331 5408 31340
rect 5356 31297 5365 31331
rect 5365 31297 5399 31331
rect 5399 31297 5408 31331
rect 5356 31288 5408 31297
rect 7196 31288 7248 31340
rect 8576 31331 8628 31340
rect 8576 31297 8585 31331
rect 8585 31297 8619 31331
rect 8619 31297 8628 31331
rect 8576 31288 8628 31297
rect 572 31220 624 31272
rect 11152 31331 11204 31340
rect 11152 31297 11161 31331
rect 11161 31297 11195 31331
rect 11195 31297 11204 31331
rect 11980 31331 12032 31340
rect 11152 31288 11204 31297
rect 11980 31297 11989 31331
rect 11989 31297 12023 31331
rect 12023 31297 12032 31331
rect 11980 31288 12032 31297
rect 13544 31424 13596 31476
rect 19156 31424 19208 31476
rect 15568 31356 15620 31408
rect 13268 31331 13320 31340
rect 13268 31297 13277 31331
rect 13277 31297 13311 31331
rect 13311 31297 13320 31331
rect 13268 31288 13320 31297
rect 13360 31331 13412 31340
rect 13360 31297 13369 31331
rect 13369 31297 13403 31331
rect 13403 31297 13412 31331
rect 13360 31288 13412 31297
rect 13728 31263 13780 31272
rect 13728 31229 13737 31263
rect 13737 31229 13771 31263
rect 13771 31229 13780 31263
rect 13728 31220 13780 31229
rect 5816 31084 5868 31136
rect 6184 31084 6236 31136
rect 7656 31084 7708 31136
rect 10140 31084 10192 31136
rect 12164 31084 12216 31136
rect 12716 31084 12768 31136
rect 13912 31084 13964 31136
rect 15476 31288 15528 31340
rect 16764 31288 16816 31340
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 18144 31356 18196 31408
rect 18880 31288 18932 31340
rect 19524 31288 19576 31340
rect 23204 31424 23256 31476
rect 28172 31467 28224 31476
rect 28172 31433 28181 31467
rect 28181 31433 28215 31467
rect 28215 31433 28224 31467
rect 28172 31424 28224 31433
rect 20628 31356 20680 31408
rect 21088 31356 21140 31408
rect 21180 31399 21232 31408
rect 21180 31365 21198 31399
rect 21198 31365 21232 31399
rect 21180 31356 21232 31365
rect 21364 31356 21416 31408
rect 16488 31220 16540 31272
rect 18512 31220 18564 31272
rect 20812 31288 20864 31340
rect 20904 31288 20956 31340
rect 21548 31288 21600 31340
rect 24860 31331 24912 31340
rect 24860 31297 24894 31331
rect 24894 31297 24912 31331
rect 24860 31288 24912 31297
rect 26700 31288 26752 31340
rect 27252 31331 27304 31340
rect 27252 31297 27261 31331
rect 27261 31297 27295 31331
rect 27295 31297 27304 31331
rect 27252 31288 27304 31297
rect 22100 31220 22152 31272
rect 23940 31220 23992 31272
rect 24492 31220 24544 31272
rect 26148 31220 26200 31272
rect 27896 31288 27948 31340
rect 28356 31331 28408 31340
rect 28356 31297 28365 31331
rect 28365 31297 28399 31331
rect 28399 31297 28408 31331
rect 28356 31288 28408 31297
rect 16948 31084 17000 31136
rect 21916 31152 21968 31204
rect 19248 31084 19300 31136
rect 19432 31127 19484 31136
rect 19432 31093 19441 31127
rect 19441 31093 19475 31127
rect 19475 31093 19484 31127
rect 19432 31084 19484 31093
rect 19892 31084 19944 31136
rect 20536 31084 20588 31136
rect 20720 31084 20772 31136
rect 23848 31127 23900 31136
rect 23848 31093 23857 31127
rect 23857 31093 23891 31127
rect 23891 31093 23900 31127
rect 25964 31127 26016 31136
rect 23848 31084 23900 31093
rect 25964 31093 25973 31127
rect 25973 31093 26007 31127
rect 26007 31093 26016 31127
rect 25964 31084 26016 31093
rect 26424 31127 26476 31136
rect 26424 31093 26433 31127
rect 26433 31093 26467 31127
rect 26467 31093 26476 31127
rect 26424 31084 26476 31093
rect 4423 30982 4475 31034
rect 4487 30982 4539 31034
rect 4551 30982 4603 31034
rect 4615 30982 4667 31034
rect 4679 30982 4731 31034
rect 11369 30982 11421 31034
rect 11433 30982 11485 31034
rect 11497 30982 11549 31034
rect 11561 30982 11613 31034
rect 11625 30982 11677 31034
rect 18315 30982 18367 31034
rect 18379 30982 18431 31034
rect 18443 30982 18495 31034
rect 18507 30982 18559 31034
rect 18571 30982 18623 31034
rect 25261 30982 25313 31034
rect 25325 30982 25377 31034
rect 25389 30982 25441 31034
rect 25453 30982 25505 31034
rect 25517 30982 25569 31034
rect 6184 30923 6236 30932
rect 6184 30889 6193 30923
rect 6193 30889 6227 30923
rect 6227 30889 6236 30923
rect 6184 30880 6236 30889
rect 7748 30880 7800 30932
rect 8484 30880 8536 30932
rect 8668 30812 8720 30864
rect 7104 30744 7156 30796
rect 11244 30880 11296 30932
rect 11796 30923 11848 30932
rect 11796 30889 11805 30923
rect 11805 30889 11839 30923
rect 11839 30889 11848 30923
rect 11796 30880 11848 30889
rect 12440 30880 12492 30932
rect 13268 30880 13320 30932
rect 17500 30855 17552 30864
rect 17500 30821 17509 30855
rect 17509 30821 17543 30855
rect 17543 30821 17552 30855
rect 17500 30812 17552 30821
rect 18972 30880 19024 30932
rect 20352 30880 20404 30932
rect 20628 30923 20680 30932
rect 20628 30889 20637 30923
rect 20637 30889 20671 30923
rect 20671 30889 20680 30923
rect 20628 30880 20680 30889
rect 21732 30880 21784 30932
rect 25964 30880 26016 30932
rect 20260 30812 20312 30864
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 11704 30744 11756 30796
rect 11888 30744 11940 30796
rect 8392 30719 8444 30728
rect 8392 30685 8401 30719
rect 8401 30685 8435 30719
rect 8435 30685 8444 30719
rect 8392 30676 8444 30685
rect 9312 30676 9364 30728
rect 12440 30744 12492 30796
rect 8484 30608 8536 30660
rect 3424 30583 3476 30592
rect 3424 30549 3433 30583
rect 3433 30549 3467 30583
rect 3467 30549 3476 30583
rect 3424 30540 3476 30549
rect 4804 30540 4856 30592
rect 5724 30583 5776 30592
rect 5724 30549 5733 30583
rect 5733 30549 5767 30583
rect 5767 30549 5776 30583
rect 5724 30540 5776 30549
rect 7380 30583 7432 30592
rect 7380 30549 7389 30583
rect 7389 30549 7423 30583
rect 7423 30549 7432 30583
rect 7380 30540 7432 30549
rect 10048 30608 10100 30660
rect 11152 30608 11204 30660
rect 12348 30676 12400 30728
rect 13176 30719 13228 30728
rect 13176 30685 13185 30719
rect 13185 30685 13219 30719
rect 13219 30685 13228 30719
rect 13176 30676 13228 30685
rect 13268 30719 13320 30728
rect 13268 30685 13277 30719
rect 13277 30685 13311 30719
rect 13311 30685 13320 30719
rect 13452 30719 13504 30728
rect 13268 30676 13320 30685
rect 13452 30685 13461 30719
rect 13461 30685 13495 30719
rect 13495 30685 13504 30719
rect 13452 30676 13504 30685
rect 8668 30540 8720 30592
rect 11060 30540 11112 30592
rect 12072 30608 12124 30660
rect 14004 30676 14056 30728
rect 14556 30676 14608 30728
rect 15108 30719 15160 30728
rect 15108 30685 15117 30719
rect 15117 30685 15151 30719
rect 15151 30685 15160 30719
rect 15108 30676 15160 30685
rect 15292 30676 15344 30728
rect 17316 30744 17368 30796
rect 18880 30787 18932 30796
rect 18880 30753 18889 30787
rect 18889 30753 18923 30787
rect 18923 30753 18932 30787
rect 18880 30744 18932 30753
rect 17684 30676 17736 30728
rect 16304 30608 16356 30660
rect 18236 30676 18288 30728
rect 19064 30676 19116 30728
rect 19892 30744 19944 30796
rect 20168 30744 20220 30796
rect 20352 30719 20404 30728
rect 17960 30608 18012 30660
rect 19616 30608 19668 30660
rect 11980 30540 12032 30592
rect 13636 30540 13688 30592
rect 14648 30583 14700 30592
rect 14648 30549 14657 30583
rect 14657 30549 14691 30583
rect 14691 30549 14700 30583
rect 14648 30540 14700 30549
rect 15660 30583 15712 30592
rect 15660 30549 15669 30583
rect 15669 30549 15703 30583
rect 15703 30549 15712 30583
rect 15660 30540 15712 30549
rect 17868 30540 17920 30592
rect 20352 30685 20361 30719
rect 20361 30685 20395 30719
rect 20395 30685 20404 30719
rect 20352 30676 20404 30685
rect 20536 30744 20588 30796
rect 22100 30744 22152 30796
rect 21180 30676 21232 30728
rect 20076 30608 20128 30660
rect 20260 30651 20312 30660
rect 20260 30617 20269 30651
rect 20269 30617 20303 30651
rect 20303 30617 20312 30651
rect 20260 30608 20312 30617
rect 20536 30608 20588 30660
rect 21916 30676 21968 30728
rect 22652 30676 22704 30728
rect 23480 30719 23532 30728
rect 23480 30685 23489 30719
rect 23489 30685 23523 30719
rect 23523 30685 23532 30719
rect 23480 30676 23532 30685
rect 23756 30719 23808 30728
rect 23756 30685 23765 30719
rect 23765 30685 23799 30719
rect 23799 30685 23808 30719
rect 23756 30676 23808 30685
rect 23940 30676 23992 30728
rect 25964 30719 26016 30728
rect 25964 30685 25973 30719
rect 25973 30685 26007 30719
rect 26007 30685 26016 30719
rect 25964 30676 26016 30685
rect 28080 30676 28132 30728
rect 21640 30608 21692 30660
rect 21732 30608 21784 30660
rect 21548 30540 21600 30592
rect 22652 30540 22704 30592
rect 23480 30540 23532 30592
rect 24308 30540 24360 30592
rect 24584 30583 24636 30592
rect 24584 30549 24593 30583
rect 24593 30549 24627 30583
rect 24627 30549 24636 30583
rect 24584 30540 24636 30549
rect 25044 30540 25096 30592
rect 26424 30583 26476 30592
rect 26424 30549 26433 30583
rect 26433 30549 26467 30583
rect 26467 30549 26476 30583
rect 26424 30540 26476 30549
rect 28264 30583 28316 30592
rect 28264 30549 28273 30583
rect 28273 30549 28307 30583
rect 28307 30549 28316 30583
rect 28264 30540 28316 30549
rect 7896 30438 7948 30490
rect 7960 30438 8012 30490
rect 8024 30438 8076 30490
rect 8088 30438 8140 30490
rect 8152 30438 8204 30490
rect 14842 30438 14894 30490
rect 14906 30438 14958 30490
rect 14970 30438 15022 30490
rect 15034 30438 15086 30490
rect 15098 30438 15150 30490
rect 21788 30438 21840 30490
rect 21852 30438 21904 30490
rect 21916 30438 21968 30490
rect 21980 30438 22032 30490
rect 22044 30438 22096 30490
rect 28734 30438 28786 30490
rect 28798 30438 28850 30490
rect 28862 30438 28914 30490
rect 28926 30438 28978 30490
rect 28990 30438 29042 30490
rect 3424 30336 3476 30388
rect 6552 30379 6604 30388
rect 6552 30345 6561 30379
rect 6561 30345 6595 30379
rect 6595 30345 6604 30379
rect 6552 30336 6604 30345
rect 9956 30336 10008 30388
rect 10140 30336 10192 30388
rect 16396 30336 16448 30388
rect 17040 30336 17092 30388
rect 17316 30336 17368 30388
rect 24584 30336 24636 30388
rect 5724 30268 5776 30320
rect 7104 30311 7156 30320
rect 7104 30277 7113 30311
rect 7113 30277 7147 30311
rect 7147 30277 7156 30311
rect 7104 30268 7156 30277
rect 7656 30268 7708 30320
rect 8944 30268 8996 30320
rect 10600 30268 10652 30320
rect 9404 30243 9456 30252
rect 9404 30209 9413 30243
rect 9413 30209 9447 30243
rect 9447 30209 9456 30243
rect 9404 30200 9456 30209
rect 10876 30268 10928 30320
rect 11152 30268 11204 30320
rect 5540 30132 5592 30184
rect 8576 30132 8628 30184
rect 10508 30132 10560 30184
rect 11704 30200 11756 30252
rect 12256 30243 12308 30252
rect 12256 30209 12265 30243
rect 12265 30209 12299 30243
rect 12299 30209 12308 30243
rect 12256 30200 12308 30209
rect 12900 30268 12952 30320
rect 10784 30132 10836 30184
rect 12624 30243 12676 30252
rect 12624 30209 12633 30243
rect 12633 30209 12667 30243
rect 12667 30209 12676 30243
rect 12624 30200 12676 30209
rect 14372 30268 14424 30320
rect 14648 30268 14700 30320
rect 20628 30268 20680 30320
rect 13360 30243 13412 30252
rect 13360 30209 13394 30243
rect 13394 30209 13412 30243
rect 13360 30200 13412 30209
rect 9772 30064 9824 30116
rect 9956 30064 10008 30116
rect 10324 30064 10376 30116
rect 11152 30107 11204 30116
rect 6828 29996 6880 30048
rect 8300 29996 8352 30048
rect 9588 30039 9640 30048
rect 9588 30005 9597 30039
rect 9597 30005 9631 30039
rect 9631 30005 9640 30039
rect 9588 29996 9640 30005
rect 10140 30039 10192 30048
rect 10140 30005 10149 30039
rect 10149 30005 10183 30039
rect 10183 30005 10192 30039
rect 11152 30073 11161 30107
rect 11161 30073 11195 30107
rect 11195 30073 11204 30107
rect 11152 30064 11204 30073
rect 12808 30064 12860 30116
rect 10140 29996 10192 30005
rect 10600 29996 10652 30048
rect 10968 30039 11020 30048
rect 10968 30005 10977 30039
rect 10977 30005 11011 30039
rect 11011 30005 11020 30039
rect 10968 29996 11020 30005
rect 12072 30039 12124 30048
rect 12072 30005 12081 30039
rect 12081 30005 12115 30039
rect 12115 30005 12124 30039
rect 12072 29996 12124 30005
rect 12164 29996 12216 30048
rect 15752 30200 15804 30252
rect 16028 30243 16080 30252
rect 16028 30209 16057 30243
rect 16057 30209 16080 30243
rect 16028 30200 16080 30209
rect 16948 30200 17000 30252
rect 14464 30107 14516 30116
rect 14464 30073 14473 30107
rect 14473 30073 14507 30107
rect 14507 30073 14516 30107
rect 16856 30132 16908 30184
rect 17224 30132 17276 30184
rect 17500 30243 17552 30252
rect 17500 30209 17509 30243
rect 17509 30209 17543 30243
rect 17543 30209 17552 30243
rect 17500 30200 17552 30209
rect 14464 30064 14516 30073
rect 14832 29996 14884 30048
rect 16488 30064 16540 30116
rect 18604 30132 18656 30184
rect 19708 30200 19760 30252
rect 20352 30243 20404 30252
rect 20352 30209 20386 30243
rect 20386 30209 20404 30243
rect 20352 30200 20404 30209
rect 23848 30268 23900 30320
rect 24216 30268 24268 30320
rect 25044 30336 25096 30388
rect 25228 30379 25280 30388
rect 25228 30345 25237 30379
rect 25237 30345 25271 30379
rect 25271 30345 25280 30379
rect 25228 30336 25280 30345
rect 27160 30379 27212 30388
rect 27160 30345 27169 30379
rect 27169 30345 27203 30379
rect 27203 30345 27212 30379
rect 27160 30336 27212 30345
rect 27344 30336 27396 30388
rect 27528 30336 27580 30388
rect 19800 30132 19852 30184
rect 15660 29996 15712 30048
rect 15936 29996 15988 30048
rect 18052 29996 18104 30048
rect 18144 29996 18196 30048
rect 18328 29996 18380 30048
rect 22284 30243 22336 30252
rect 22284 30209 22318 30243
rect 22318 30209 22336 30243
rect 22284 30200 22336 30209
rect 21180 30132 21232 30184
rect 21272 30064 21324 30116
rect 21180 29996 21232 30048
rect 26608 30200 26660 30252
rect 26976 30200 27028 30252
rect 27528 30243 27580 30252
rect 27528 30209 27537 30243
rect 27537 30209 27571 30243
rect 27571 30209 27580 30243
rect 27528 30200 27580 30209
rect 23848 30175 23900 30184
rect 23848 30141 23857 30175
rect 23857 30141 23891 30175
rect 23891 30141 23900 30175
rect 23848 30132 23900 30141
rect 26700 30132 26752 30184
rect 25688 30064 25740 30116
rect 23388 30039 23440 30048
rect 23388 30005 23397 30039
rect 23397 30005 23431 30039
rect 23431 30005 23440 30039
rect 23388 29996 23440 30005
rect 25044 29996 25096 30048
rect 4423 29894 4475 29946
rect 4487 29894 4539 29946
rect 4551 29894 4603 29946
rect 4615 29894 4667 29946
rect 4679 29894 4731 29946
rect 11369 29894 11421 29946
rect 11433 29894 11485 29946
rect 11497 29894 11549 29946
rect 11561 29894 11613 29946
rect 11625 29894 11677 29946
rect 18315 29894 18367 29946
rect 18379 29894 18431 29946
rect 18443 29894 18495 29946
rect 18507 29894 18559 29946
rect 18571 29894 18623 29946
rect 25261 29894 25313 29946
rect 25325 29894 25377 29946
rect 25389 29894 25441 29946
rect 25453 29894 25505 29946
rect 25517 29894 25569 29946
rect 5540 29792 5592 29844
rect 5816 29792 5868 29844
rect 8300 29792 8352 29844
rect 8484 29835 8536 29844
rect 8484 29801 8493 29835
rect 8493 29801 8527 29835
rect 8527 29801 8536 29835
rect 8484 29792 8536 29801
rect 9634 29792 9686 29844
rect 12532 29792 12584 29844
rect 12624 29792 12676 29844
rect 14280 29792 14332 29844
rect 4804 29656 4856 29708
rect 11060 29724 11112 29776
rect 11612 29724 11664 29776
rect 1584 29631 1636 29640
rect 1584 29597 1593 29631
rect 1593 29597 1627 29631
rect 1627 29597 1636 29631
rect 1584 29588 1636 29597
rect 5724 29588 5776 29640
rect 10140 29588 10192 29640
rect 9588 29563 9640 29572
rect 5264 29495 5316 29504
rect 5264 29461 5273 29495
rect 5273 29461 5307 29495
rect 5307 29461 5316 29495
rect 5264 29452 5316 29461
rect 6920 29495 6972 29504
rect 6920 29461 6929 29495
rect 6929 29461 6963 29495
rect 6963 29461 6972 29495
rect 6920 29452 6972 29461
rect 9588 29529 9597 29563
rect 9597 29529 9631 29563
rect 9631 29529 9640 29563
rect 9588 29520 9640 29529
rect 10508 29656 10560 29708
rect 10784 29656 10836 29708
rect 11336 29699 11388 29708
rect 11336 29665 11345 29699
rect 11345 29665 11379 29699
rect 11379 29665 11388 29699
rect 11336 29656 11388 29665
rect 13452 29724 13504 29776
rect 13728 29767 13780 29776
rect 13728 29733 13737 29767
rect 13737 29733 13771 29767
rect 13771 29733 13780 29767
rect 13728 29724 13780 29733
rect 15568 29792 15620 29844
rect 15292 29724 15344 29776
rect 10416 29631 10468 29640
rect 10416 29597 10425 29631
rect 10425 29597 10459 29631
rect 10459 29597 10468 29631
rect 10416 29588 10468 29597
rect 10876 29631 10928 29640
rect 10876 29597 10885 29631
rect 10885 29597 10919 29631
rect 10919 29597 10928 29631
rect 10876 29588 10928 29597
rect 11060 29588 11112 29640
rect 10784 29520 10836 29572
rect 9956 29452 10008 29504
rect 10324 29452 10376 29504
rect 10600 29495 10652 29504
rect 10600 29461 10609 29495
rect 10609 29461 10643 29495
rect 10643 29461 10652 29495
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 12164 29588 12216 29640
rect 12440 29520 12492 29572
rect 12992 29520 13044 29572
rect 15568 29656 15620 29708
rect 15844 29792 15896 29844
rect 16396 29792 16448 29844
rect 20444 29792 20496 29844
rect 17040 29767 17092 29776
rect 17040 29733 17049 29767
rect 17049 29733 17083 29767
rect 17083 29733 17092 29767
rect 17040 29724 17092 29733
rect 18788 29724 18840 29776
rect 17316 29656 17368 29708
rect 18696 29656 18748 29708
rect 19432 29656 19484 29708
rect 19616 29656 19668 29708
rect 21272 29724 21324 29776
rect 20812 29656 20864 29708
rect 15016 29631 15068 29640
rect 15016 29597 15025 29631
rect 15025 29597 15059 29631
rect 15059 29597 15068 29631
rect 15016 29588 15068 29597
rect 15384 29588 15436 29640
rect 16488 29588 16540 29640
rect 17408 29588 17460 29640
rect 18052 29588 18104 29640
rect 19708 29588 19760 29640
rect 19892 29588 19944 29640
rect 21088 29588 21140 29640
rect 22376 29631 22428 29640
rect 22376 29597 22385 29631
rect 22385 29597 22419 29631
rect 22419 29597 22428 29631
rect 22376 29588 22428 29597
rect 14004 29520 14056 29572
rect 14832 29520 14884 29572
rect 15752 29520 15804 29572
rect 18144 29520 18196 29572
rect 18328 29520 18380 29572
rect 20168 29520 20220 29572
rect 20444 29520 20496 29572
rect 10600 29452 10652 29461
rect 14648 29452 14700 29504
rect 16948 29452 17000 29504
rect 17960 29452 18012 29504
rect 18512 29452 18564 29504
rect 18696 29452 18748 29504
rect 21088 29452 21140 29504
rect 23388 29724 23440 29776
rect 22928 29588 22980 29640
rect 24124 29588 24176 29640
rect 23848 29520 23900 29572
rect 25964 29588 26016 29640
rect 28264 29588 28316 29640
rect 28632 29588 28684 29640
rect 25136 29520 25188 29572
rect 24676 29452 24728 29504
rect 25044 29452 25096 29504
rect 27988 29452 28040 29504
rect 7896 29350 7948 29402
rect 7960 29350 8012 29402
rect 8024 29350 8076 29402
rect 8088 29350 8140 29402
rect 8152 29350 8204 29402
rect 14842 29350 14894 29402
rect 14906 29350 14958 29402
rect 14970 29350 15022 29402
rect 15034 29350 15086 29402
rect 15098 29350 15150 29402
rect 21788 29350 21840 29402
rect 21852 29350 21904 29402
rect 21916 29350 21968 29402
rect 21980 29350 22032 29402
rect 22044 29350 22096 29402
rect 28734 29350 28786 29402
rect 28798 29350 28850 29402
rect 28862 29350 28914 29402
rect 28926 29350 28978 29402
rect 28990 29350 29042 29402
rect 5264 29248 5316 29300
rect 6920 29248 6972 29300
rect 8484 29291 8536 29300
rect 8484 29257 8493 29291
rect 8493 29257 8527 29291
rect 8527 29257 8536 29291
rect 8484 29248 8536 29257
rect 8760 29248 8812 29300
rect 9864 29248 9916 29300
rect 9496 29180 9548 29232
rect 10692 29180 10744 29232
rect 16580 29248 16632 29300
rect 9864 29112 9916 29164
rect 10508 29112 10560 29164
rect 12164 29180 12216 29232
rect 12256 29155 12308 29164
rect 12256 29121 12265 29155
rect 12265 29121 12299 29155
rect 12299 29121 12308 29155
rect 12256 29112 12308 29121
rect 12440 29155 12492 29164
rect 12440 29121 12464 29155
rect 12464 29121 12492 29155
rect 12440 29112 12492 29121
rect 12624 29155 12676 29164
rect 12624 29121 12633 29155
rect 12633 29121 12667 29155
rect 12667 29121 12676 29155
rect 13544 29180 13596 29232
rect 15016 29180 15068 29232
rect 12624 29112 12676 29121
rect 14464 29112 14516 29164
rect 15384 29180 15436 29232
rect 15476 29180 15528 29232
rect 14740 29044 14792 29096
rect 15752 29112 15804 29164
rect 16764 29180 16816 29232
rect 18880 29248 18932 29300
rect 20444 29248 20496 29300
rect 20720 29180 20772 29232
rect 17316 29155 17368 29164
rect 17316 29121 17325 29155
rect 17325 29121 17359 29155
rect 17359 29121 17368 29155
rect 17316 29112 17368 29121
rect 17500 29155 17552 29164
rect 17500 29121 17509 29155
rect 17509 29121 17543 29155
rect 17543 29121 17552 29155
rect 17500 29112 17552 29121
rect 17960 29112 18012 29164
rect 16948 29044 17000 29096
rect 18052 29044 18104 29096
rect 18788 29112 18840 29164
rect 18880 29112 18932 29164
rect 21088 29248 21140 29300
rect 21272 29248 21324 29300
rect 25136 29248 25188 29300
rect 26884 29248 26936 29300
rect 20996 29180 21048 29232
rect 24768 29180 24820 29232
rect 23112 29155 23164 29164
rect 23112 29121 23130 29155
rect 23130 29121 23164 29155
rect 23112 29112 23164 29121
rect 22376 29044 22428 29096
rect 23388 29087 23440 29096
rect 23388 29053 23397 29087
rect 23397 29053 23431 29087
rect 23431 29053 23440 29087
rect 23848 29087 23900 29096
rect 23388 29044 23440 29053
rect 23848 29053 23857 29087
rect 23857 29053 23891 29087
rect 23891 29053 23900 29087
rect 23848 29044 23900 29053
rect 8944 29019 8996 29028
rect 8944 28985 8953 29019
rect 8953 28985 8987 29019
rect 8987 28985 8996 29019
rect 8944 28976 8996 28985
rect 8760 28908 8812 28960
rect 9220 28908 9272 28960
rect 11060 28976 11112 29028
rect 12992 28976 13044 29028
rect 13084 28976 13136 29028
rect 10600 28908 10652 28960
rect 10968 28951 11020 28960
rect 10968 28917 10977 28951
rect 10977 28917 11011 28951
rect 11011 28917 11020 28951
rect 10968 28908 11020 28917
rect 11244 28908 11296 28960
rect 14464 28951 14516 28960
rect 14464 28917 14473 28951
rect 14473 28917 14507 28951
rect 14507 28917 14516 28951
rect 16764 28976 16816 29028
rect 14464 28908 14516 28917
rect 16396 28908 16448 28960
rect 16488 28908 16540 28960
rect 20352 28976 20404 29028
rect 21640 28976 21692 29028
rect 19432 28908 19484 28960
rect 19616 28951 19668 28960
rect 19616 28917 19625 28951
rect 19625 28917 19659 28951
rect 19659 28917 19668 28951
rect 19616 28908 19668 28917
rect 19892 28908 19944 28960
rect 20260 28908 20312 28960
rect 20444 28908 20496 28960
rect 23848 28908 23900 28960
rect 27160 29112 27212 29164
rect 27528 29155 27580 29164
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 27620 29155 27672 29164
rect 27620 29121 27655 29155
rect 27655 29121 27672 29155
rect 27620 29112 27672 29121
rect 27804 29155 27856 29164
rect 27804 29121 27813 29155
rect 27813 29121 27847 29155
rect 27847 29121 27856 29155
rect 27804 29112 27856 29121
rect 25964 29087 26016 29096
rect 24952 28976 25004 29028
rect 25964 29053 25973 29087
rect 25973 29053 26007 29087
rect 26007 29053 26016 29087
rect 25964 29044 26016 29053
rect 26700 28976 26752 29028
rect 26884 28976 26936 29028
rect 28356 28951 28408 28960
rect 28356 28917 28365 28951
rect 28365 28917 28399 28951
rect 28399 28917 28408 28951
rect 28356 28908 28408 28917
rect 28632 28908 28684 28960
rect 4423 28806 4475 28858
rect 4487 28806 4539 28858
rect 4551 28806 4603 28858
rect 4615 28806 4667 28858
rect 4679 28806 4731 28858
rect 11369 28806 11421 28858
rect 11433 28806 11485 28858
rect 11497 28806 11549 28858
rect 11561 28806 11613 28858
rect 11625 28806 11677 28858
rect 18315 28806 18367 28858
rect 18379 28806 18431 28858
rect 18443 28806 18495 28858
rect 18507 28806 18559 28858
rect 18571 28806 18623 28858
rect 25261 28806 25313 28858
rect 25325 28806 25377 28858
rect 25389 28806 25441 28858
rect 25453 28806 25505 28858
rect 25517 28806 25569 28858
rect 8392 28704 8444 28756
rect 8668 28704 8720 28756
rect 9496 28704 9548 28756
rect 11060 28704 11112 28756
rect 11152 28704 11204 28756
rect 11612 28747 11664 28756
rect 11612 28713 11621 28747
rect 11621 28713 11655 28747
rect 11655 28713 11664 28747
rect 11612 28704 11664 28713
rect 13176 28704 13228 28756
rect 20076 28704 20128 28756
rect 20260 28704 20312 28756
rect 23664 28704 23716 28756
rect 23848 28704 23900 28756
rect 25504 28704 25556 28756
rect 7104 28636 7156 28688
rect 7748 28636 7800 28688
rect 12164 28636 12216 28688
rect 9496 28568 9548 28620
rect 11244 28568 11296 28620
rect 14556 28636 14608 28688
rect 15016 28636 15068 28688
rect 15476 28636 15528 28688
rect 16764 28636 16816 28688
rect 1584 28543 1636 28552
rect 1584 28509 1593 28543
rect 1593 28509 1627 28543
rect 1627 28509 1636 28543
rect 1584 28500 1636 28509
rect 8944 28500 8996 28552
rect 10140 28543 10192 28552
rect 10140 28509 10149 28543
rect 10149 28509 10183 28543
rect 10183 28509 10192 28543
rect 10140 28500 10192 28509
rect 10416 28500 10468 28552
rect 12348 28500 12400 28552
rect 12532 28543 12584 28552
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 13820 28568 13872 28620
rect 9680 28432 9732 28484
rect 11428 28475 11480 28484
rect 11428 28441 11437 28475
rect 11437 28441 11471 28475
rect 11471 28441 11480 28475
rect 11428 28432 11480 28441
rect 11796 28432 11848 28484
rect 13728 28543 13780 28552
rect 13728 28509 13737 28543
rect 13737 28509 13771 28543
rect 13771 28509 13780 28543
rect 13728 28500 13780 28509
rect 14556 28500 14608 28552
rect 15292 28568 15344 28620
rect 16672 28568 16724 28620
rect 17776 28568 17828 28620
rect 19432 28636 19484 28688
rect 20812 28636 20864 28688
rect 22376 28636 22428 28688
rect 15108 28543 15160 28552
rect 15108 28509 15117 28543
rect 15117 28509 15151 28543
rect 15151 28509 15160 28543
rect 11888 28364 11940 28416
rect 13084 28364 13136 28416
rect 13268 28364 13320 28416
rect 14004 28432 14056 28484
rect 15108 28500 15160 28509
rect 15384 28500 15436 28552
rect 19340 28568 19392 28620
rect 20444 28611 20496 28620
rect 20444 28577 20453 28611
rect 20453 28577 20487 28611
rect 20487 28577 20496 28611
rect 20444 28568 20496 28577
rect 17592 28432 17644 28484
rect 17776 28432 17828 28484
rect 18512 28432 18564 28484
rect 22376 28543 22428 28552
rect 22376 28509 22385 28543
rect 22385 28509 22419 28543
rect 22419 28509 22428 28543
rect 22376 28500 22428 28509
rect 16120 28364 16172 28416
rect 16304 28364 16356 28416
rect 19248 28432 19300 28484
rect 22008 28432 22060 28484
rect 22284 28432 22336 28484
rect 23112 28611 23164 28620
rect 23112 28577 23121 28611
rect 23121 28577 23155 28611
rect 23155 28577 23164 28611
rect 23112 28568 23164 28577
rect 22928 28500 22980 28552
rect 24400 28568 24452 28620
rect 24676 28500 24728 28552
rect 25412 28500 25464 28552
rect 26516 28432 26568 28484
rect 18788 28364 18840 28416
rect 20168 28407 20220 28416
rect 20168 28373 20177 28407
rect 20177 28373 20211 28407
rect 20211 28373 20220 28407
rect 20168 28364 20220 28373
rect 20444 28364 20496 28416
rect 21088 28364 21140 28416
rect 24952 28364 25004 28416
rect 25228 28364 25280 28416
rect 25596 28364 25648 28416
rect 26148 28364 26200 28416
rect 27804 28407 27856 28416
rect 27804 28373 27813 28407
rect 27813 28373 27847 28407
rect 27847 28373 27856 28407
rect 27804 28364 27856 28373
rect 28356 28407 28408 28416
rect 28356 28373 28365 28407
rect 28365 28373 28399 28407
rect 28399 28373 28408 28407
rect 28356 28364 28408 28373
rect 7896 28262 7948 28314
rect 7960 28262 8012 28314
rect 8024 28262 8076 28314
rect 8088 28262 8140 28314
rect 8152 28262 8204 28314
rect 14842 28262 14894 28314
rect 14906 28262 14958 28314
rect 14970 28262 15022 28314
rect 15034 28262 15086 28314
rect 15098 28262 15150 28314
rect 21788 28262 21840 28314
rect 21852 28262 21904 28314
rect 21916 28262 21968 28314
rect 21980 28262 22032 28314
rect 22044 28262 22096 28314
rect 28734 28262 28786 28314
rect 28798 28262 28850 28314
rect 28862 28262 28914 28314
rect 28926 28262 28978 28314
rect 28990 28262 29042 28314
rect 9312 28160 9364 28212
rect 10048 28203 10100 28212
rect 10048 28169 10057 28203
rect 10057 28169 10091 28203
rect 10091 28169 10100 28203
rect 10048 28160 10100 28169
rect 10140 28160 10192 28212
rect 10508 28203 10560 28212
rect 10508 28169 10517 28203
rect 10517 28169 10551 28203
rect 10551 28169 10560 28203
rect 10508 28160 10560 28169
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 11796 28160 11848 28212
rect 13084 28203 13136 28212
rect 7380 28092 7432 28144
rect 9220 28092 9272 28144
rect 10324 28092 10376 28144
rect 11888 28092 11940 28144
rect 13084 28169 13093 28203
rect 13093 28169 13127 28203
rect 13127 28169 13136 28203
rect 13084 28160 13136 28169
rect 17684 28160 17736 28212
rect 18236 28203 18288 28212
rect 18236 28169 18245 28203
rect 18245 28169 18279 28203
rect 18279 28169 18288 28203
rect 18236 28160 18288 28169
rect 19064 28160 19116 28212
rect 12348 28135 12400 28144
rect 12348 28101 12373 28135
rect 12373 28101 12400 28135
rect 12348 28092 12400 28101
rect 14648 28092 14700 28144
rect 16304 28092 16356 28144
rect 12532 28024 12584 28076
rect 12992 28067 13044 28076
rect 12992 28033 13001 28067
rect 13001 28033 13035 28067
rect 13035 28033 13044 28067
rect 12992 28024 13044 28033
rect 6828 27956 6880 28008
rect 11796 27956 11848 28008
rect 11980 27956 12032 28008
rect 12256 27956 12308 28008
rect 13268 27999 13320 28008
rect 13268 27965 13277 27999
rect 13277 27965 13311 27999
rect 13311 27965 13320 27999
rect 13268 27956 13320 27965
rect 13544 27956 13596 28008
rect 11612 27888 11664 27940
rect 14740 28024 14792 28076
rect 16028 28024 16080 28076
rect 17684 28024 17736 28076
rect 17776 28067 17828 28076
rect 17776 28033 17785 28067
rect 17785 28033 17819 28067
rect 17819 28033 17828 28067
rect 17776 28024 17828 28033
rect 19064 28024 19116 28076
rect 19248 28092 19300 28144
rect 27804 28160 27856 28212
rect 19524 28092 19576 28144
rect 19984 28092 20036 28144
rect 20812 28092 20864 28144
rect 21180 28135 21232 28144
rect 21180 28101 21198 28135
rect 21198 28101 21232 28135
rect 21180 28092 21232 28101
rect 21732 28092 21784 28144
rect 22744 28092 22796 28144
rect 20260 28024 20312 28076
rect 14464 27956 14516 28008
rect 14648 27956 14700 28008
rect 16120 27956 16172 28008
rect 17040 27956 17092 28008
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 8484 27820 8536 27872
rect 10416 27820 10468 27872
rect 10600 27820 10652 27872
rect 12256 27820 12308 27872
rect 13912 27888 13964 27940
rect 14096 27888 14148 27940
rect 14556 27888 14608 27940
rect 14832 27888 14884 27940
rect 13084 27820 13136 27872
rect 14924 27820 14976 27872
rect 15936 27820 15988 27872
rect 17040 27820 17092 27872
rect 17500 27956 17552 28008
rect 17960 27956 18012 28008
rect 19708 27956 19760 28008
rect 19984 27956 20036 28008
rect 21548 28024 21600 28076
rect 23296 28024 23348 28076
rect 23756 28024 23808 28076
rect 24492 28092 24544 28144
rect 26332 28092 26384 28144
rect 26884 28092 26936 28144
rect 27988 28092 28040 28144
rect 27344 28067 27396 28076
rect 27344 28033 27353 28067
rect 27353 28033 27387 28067
rect 27387 28033 27396 28067
rect 27344 28024 27396 28033
rect 27620 28067 27672 28076
rect 27620 28033 27629 28067
rect 27629 28033 27663 28067
rect 27663 28033 27672 28067
rect 27620 28024 27672 28033
rect 27804 28024 27856 28076
rect 22376 27956 22428 28008
rect 23388 27999 23440 28008
rect 23388 27965 23397 27999
rect 23397 27965 23431 27999
rect 23431 27965 23440 27999
rect 23388 27956 23440 27965
rect 23848 27999 23900 28008
rect 23848 27965 23857 27999
rect 23857 27965 23891 27999
rect 23891 27965 23900 27999
rect 23848 27956 23900 27965
rect 24952 27956 25004 28008
rect 17592 27888 17644 27940
rect 18604 27820 18656 27872
rect 20076 27863 20128 27872
rect 20076 27829 20085 27863
rect 20085 27829 20119 27863
rect 20119 27829 20128 27863
rect 20076 27820 20128 27829
rect 20812 27820 20864 27872
rect 21548 27820 21600 27872
rect 22376 27820 22428 27872
rect 25228 27931 25280 27940
rect 25228 27897 25237 27931
rect 25237 27897 25271 27931
rect 25271 27897 25280 27931
rect 25228 27888 25280 27897
rect 25504 27956 25556 28008
rect 26148 27956 26200 28008
rect 26792 27888 26844 27940
rect 27436 27931 27488 27940
rect 27436 27897 27445 27931
rect 27445 27897 27479 27931
rect 27479 27897 27488 27931
rect 27436 27888 27488 27897
rect 23848 27820 23900 27872
rect 25044 27820 25096 27872
rect 25320 27820 25372 27872
rect 26056 27820 26108 27872
rect 26424 27820 26476 27872
rect 28264 27863 28316 27872
rect 28264 27829 28273 27863
rect 28273 27829 28307 27863
rect 28307 27829 28316 27863
rect 28264 27820 28316 27829
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 7748 27616 7800 27668
rect 8484 27659 8536 27668
rect 8484 27625 8493 27659
rect 8493 27625 8527 27659
rect 8527 27625 8536 27659
rect 8484 27616 8536 27625
rect 9220 27616 9272 27668
rect 12164 27659 12216 27668
rect 9680 27548 9732 27600
rect 10324 27548 10376 27600
rect 10508 27548 10560 27600
rect 11704 27548 11756 27600
rect 12164 27625 12173 27659
rect 12173 27625 12207 27659
rect 12207 27625 12216 27659
rect 12164 27616 12216 27625
rect 12256 27616 12308 27668
rect 12808 27548 12860 27600
rect 14740 27616 14792 27668
rect 14372 27548 14424 27600
rect 15936 27616 15988 27668
rect 16028 27616 16080 27668
rect 16304 27616 16356 27668
rect 23848 27616 23900 27668
rect 24860 27616 24912 27668
rect 25688 27616 25740 27668
rect 25872 27616 25924 27668
rect 26056 27616 26108 27668
rect 27896 27616 27948 27668
rect 17132 27548 17184 27600
rect 17684 27548 17736 27600
rect 19064 27548 19116 27600
rect 19892 27548 19944 27600
rect 11336 27480 11388 27532
rect 13544 27480 13596 27532
rect 13820 27480 13872 27532
rect 14556 27480 14608 27532
rect 14832 27480 14884 27532
rect 9680 27344 9732 27396
rect 12900 27344 12952 27396
rect 13360 27387 13412 27396
rect 13360 27353 13369 27387
rect 13369 27353 13403 27387
rect 13403 27353 13412 27387
rect 13360 27344 13412 27353
rect 8300 27276 8352 27328
rect 10692 27276 10744 27328
rect 11336 27276 11388 27328
rect 13544 27319 13596 27328
rect 14924 27455 14976 27464
rect 14924 27421 14933 27455
rect 14933 27421 14967 27455
rect 14967 27421 14976 27455
rect 14924 27412 14976 27421
rect 16028 27480 16080 27532
rect 15292 27412 15344 27464
rect 17500 27412 17552 27464
rect 19340 27480 19392 27532
rect 19524 27412 19576 27464
rect 19708 27412 19760 27464
rect 20168 27455 20220 27464
rect 20168 27421 20177 27455
rect 20177 27421 20211 27455
rect 20211 27421 20220 27455
rect 20168 27412 20220 27421
rect 20996 27548 21048 27600
rect 22560 27548 22612 27600
rect 20628 27455 20680 27464
rect 20628 27421 20637 27455
rect 20637 27421 20671 27455
rect 20671 27421 20680 27455
rect 20628 27412 20680 27421
rect 20720 27412 20772 27464
rect 22376 27412 22428 27464
rect 23572 27548 23624 27600
rect 23020 27412 23072 27464
rect 23296 27412 23348 27464
rect 23940 27412 23992 27464
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 26056 27412 26108 27464
rect 13820 27344 13872 27396
rect 16120 27344 16172 27396
rect 16948 27344 17000 27396
rect 17132 27344 17184 27396
rect 13544 27285 13569 27319
rect 13569 27285 13596 27319
rect 13544 27276 13596 27285
rect 14188 27276 14240 27328
rect 16672 27276 16724 27328
rect 19064 27344 19116 27396
rect 19708 27276 19760 27328
rect 21732 27276 21784 27328
rect 22652 27344 22704 27396
rect 23388 27344 23440 27396
rect 25044 27344 25096 27396
rect 26792 27344 26844 27396
rect 27068 27344 27120 27396
rect 27896 27344 27948 27396
rect 23572 27276 23624 27328
rect 27344 27276 27396 27328
rect 27528 27276 27580 27328
rect 28356 27319 28408 27328
rect 28356 27285 28365 27319
rect 28365 27285 28399 27319
rect 28399 27285 28408 27319
rect 28356 27276 28408 27285
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 9496 27115 9548 27124
rect 9496 27081 9505 27115
rect 9505 27081 9539 27115
rect 9539 27081 9548 27115
rect 9496 27072 9548 27081
rect 9680 27072 9732 27124
rect 10600 27115 10652 27124
rect 10600 27081 10609 27115
rect 10609 27081 10643 27115
rect 10643 27081 10652 27115
rect 10600 27072 10652 27081
rect 11152 27115 11204 27124
rect 11152 27081 11161 27115
rect 11161 27081 11195 27115
rect 11195 27081 11204 27115
rect 11152 27072 11204 27081
rect 11888 27072 11940 27124
rect 12624 27072 12676 27124
rect 14740 27072 14792 27124
rect 15476 27072 15528 27124
rect 16488 27072 16540 27124
rect 17868 27072 17920 27124
rect 12348 27004 12400 27056
rect 14372 27047 14424 27056
rect 14372 27013 14381 27047
rect 14381 27013 14415 27047
rect 14415 27013 14424 27047
rect 14372 27004 14424 27013
rect 15568 27004 15620 27056
rect 21364 27072 21416 27124
rect 12992 26936 13044 26988
rect 8576 26868 8628 26920
rect 13636 26936 13688 26988
rect 13820 26936 13872 26988
rect 14832 26979 14884 26988
rect 14832 26945 14841 26979
rect 14841 26945 14875 26979
rect 14875 26945 14884 26979
rect 14832 26936 14884 26945
rect 15292 26979 15344 26988
rect 13912 26868 13964 26920
rect 15292 26945 15301 26979
rect 15301 26945 15335 26979
rect 15335 26945 15344 26979
rect 15292 26936 15344 26945
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 18328 27004 18380 27056
rect 18696 27004 18748 27056
rect 19248 27004 19300 27056
rect 19616 27004 19668 27056
rect 16120 26936 16172 26945
rect 17684 26936 17736 26988
rect 20352 26979 20404 26988
rect 20352 26945 20386 26979
rect 20386 26945 20404 26979
rect 20352 26936 20404 26945
rect 20536 27004 20588 27056
rect 22284 27072 22336 27124
rect 23848 27115 23900 27124
rect 23848 27081 23857 27115
rect 23857 27081 23891 27115
rect 23891 27081 23900 27115
rect 23848 27072 23900 27081
rect 24124 27072 24176 27124
rect 25044 27072 25096 27124
rect 25136 27072 25188 27124
rect 25872 27072 25924 27124
rect 22284 26979 22336 26988
rect 22284 26945 22318 26979
rect 22318 26945 22336 26979
rect 22284 26936 22336 26945
rect 24584 26936 24636 26988
rect 25596 26936 25648 26988
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 16764 26868 16816 26920
rect 17408 26911 17460 26920
rect 17408 26877 17417 26911
rect 17417 26877 17451 26911
rect 17451 26877 17460 26911
rect 17408 26868 17460 26877
rect 19248 26868 19300 26920
rect 19340 26868 19392 26920
rect 19984 26868 20036 26920
rect 22008 26911 22060 26920
rect 22008 26877 22017 26911
rect 22017 26877 22051 26911
rect 22051 26877 22060 26911
rect 22008 26868 22060 26877
rect 25228 26911 25280 26920
rect 25228 26877 25237 26911
rect 25237 26877 25271 26911
rect 25271 26877 25280 26911
rect 25228 26868 25280 26877
rect 25688 26868 25740 26920
rect 26608 26936 26660 26988
rect 27252 26936 27304 26988
rect 27528 26936 27580 26988
rect 27620 26979 27672 26988
rect 27620 26945 27629 26979
rect 27629 26945 27663 26979
rect 27663 26945 27672 26979
rect 27620 26936 27672 26945
rect 28080 26936 28132 26988
rect 26424 26868 26476 26920
rect 27160 26868 27212 26920
rect 15752 26800 15804 26852
rect 9772 26732 9824 26784
rect 13360 26775 13412 26784
rect 13360 26741 13369 26775
rect 13369 26741 13403 26775
rect 13403 26741 13412 26775
rect 13360 26732 13412 26741
rect 14188 26775 14240 26784
rect 14188 26741 14197 26775
rect 14197 26741 14231 26775
rect 14231 26741 14240 26775
rect 14188 26732 14240 26741
rect 14556 26732 14608 26784
rect 15568 26732 15620 26784
rect 16304 26800 16356 26852
rect 16120 26732 16172 26784
rect 16764 26732 16816 26784
rect 19800 26732 19852 26784
rect 19984 26732 20036 26784
rect 21732 26800 21784 26852
rect 23020 26800 23072 26852
rect 23940 26800 23992 26852
rect 25504 26800 25556 26852
rect 26608 26800 26660 26852
rect 27528 26843 27580 26852
rect 27528 26809 27537 26843
rect 27537 26809 27571 26843
rect 27571 26809 27580 26843
rect 27528 26800 27580 26809
rect 21272 26732 21324 26784
rect 22284 26732 22336 26784
rect 23664 26732 23716 26784
rect 25044 26732 25096 26784
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 10600 26528 10652 26580
rect 10692 26528 10744 26580
rect 12072 26571 12124 26580
rect 12072 26537 12081 26571
rect 12081 26537 12115 26571
rect 12115 26537 12124 26571
rect 12072 26528 12124 26537
rect 12348 26528 12400 26580
rect 11152 26460 11204 26512
rect 12348 26392 12400 26444
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 9864 26324 9916 26333
rect 12624 26435 12676 26444
rect 12624 26401 12633 26435
rect 12633 26401 12667 26435
rect 12667 26401 12676 26435
rect 14188 26528 14240 26580
rect 14372 26460 14424 26512
rect 14648 26460 14700 26512
rect 15660 26460 15712 26512
rect 12624 26392 12676 26401
rect 13360 26392 13412 26444
rect 11888 26256 11940 26308
rect 13912 26256 13964 26308
rect 14648 26299 14700 26308
rect 14648 26265 14657 26299
rect 14657 26265 14691 26299
rect 14691 26265 14700 26299
rect 14648 26256 14700 26265
rect 15108 26324 15160 26376
rect 15568 26367 15620 26376
rect 15568 26333 15577 26367
rect 15577 26333 15611 26367
rect 15611 26333 15620 26367
rect 23388 26528 23440 26580
rect 16120 26460 16172 26512
rect 16488 26460 16540 26512
rect 16580 26460 16632 26512
rect 17132 26460 17184 26512
rect 18696 26460 18748 26512
rect 20812 26460 20864 26512
rect 20996 26460 21048 26512
rect 23204 26503 23256 26512
rect 23204 26469 23213 26503
rect 23213 26469 23247 26503
rect 23247 26469 23256 26503
rect 23204 26460 23256 26469
rect 17500 26435 17552 26444
rect 15568 26324 15620 26333
rect 16120 26324 16172 26376
rect 16672 26324 16724 26376
rect 17500 26401 17509 26435
rect 17509 26401 17543 26435
rect 17543 26401 17552 26435
rect 17500 26392 17552 26401
rect 18512 26392 18564 26444
rect 19524 26435 19576 26444
rect 19524 26401 19533 26435
rect 19533 26401 19567 26435
rect 19567 26401 19576 26435
rect 19524 26392 19576 26401
rect 28356 26571 28408 26580
rect 28356 26537 28365 26571
rect 28365 26537 28399 26571
rect 28399 26537 28408 26571
rect 28356 26528 28408 26537
rect 19800 26367 19852 26376
rect 16304 26188 16356 26240
rect 17776 26299 17828 26308
rect 17776 26265 17810 26299
rect 17810 26265 17828 26299
rect 17776 26256 17828 26265
rect 19340 26256 19392 26308
rect 19800 26333 19834 26367
rect 19834 26333 19852 26367
rect 19800 26324 19852 26333
rect 21088 26324 21140 26376
rect 21180 26324 21232 26376
rect 20720 26256 20772 26308
rect 22100 26256 22152 26308
rect 18604 26188 18656 26240
rect 18972 26188 19024 26240
rect 20168 26188 20220 26240
rect 22192 26188 22244 26240
rect 23020 26324 23072 26376
rect 23388 26367 23440 26376
rect 23388 26333 23397 26367
rect 23397 26333 23431 26367
rect 23431 26333 23440 26367
rect 23388 26324 23440 26333
rect 23756 26460 23808 26512
rect 24584 26503 24636 26512
rect 24584 26469 24593 26503
rect 24593 26469 24627 26503
rect 24627 26469 24636 26503
rect 24584 26460 24636 26469
rect 26056 26392 26108 26444
rect 23848 26367 23900 26376
rect 23848 26333 23857 26367
rect 23857 26333 23891 26367
rect 23891 26333 23900 26367
rect 23848 26324 23900 26333
rect 24400 26324 24452 26376
rect 23664 26299 23716 26308
rect 23664 26265 23699 26299
rect 23699 26265 23716 26299
rect 23664 26256 23716 26265
rect 23112 26188 23164 26240
rect 23296 26188 23348 26240
rect 25596 26256 25648 26308
rect 26056 26256 26108 26308
rect 26148 26256 26200 26308
rect 27160 26256 27212 26308
rect 23940 26188 23992 26240
rect 24860 26188 24912 26240
rect 25044 26188 25096 26240
rect 26240 26188 26292 26240
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 9680 25984 9732 26036
rect 10416 26027 10468 26036
rect 10416 25993 10425 26027
rect 10425 25993 10459 26027
rect 10459 25993 10468 26027
rect 10416 25984 10468 25993
rect 12164 25984 12216 26036
rect 14740 25984 14792 26036
rect 15200 25984 15252 26036
rect 16672 25984 16724 26036
rect 13544 25916 13596 25968
rect 10600 25848 10652 25900
rect 14648 25891 14700 25900
rect 14648 25857 14657 25891
rect 14657 25857 14691 25891
rect 14691 25857 14700 25891
rect 14648 25848 14700 25857
rect 14740 25848 14792 25900
rect 15844 25916 15896 25968
rect 16212 25916 16264 25968
rect 15660 25780 15712 25832
rect 16028 25780 16080 25832
rect 16764 25916 16816 25968
rect 17776 25984 17828 26036
rect 19616 25984 19668 26036
rect 19708 25984 19760 26036
rect 17224 25780 17276 25832
rect 17500 25891 17552 25900
rect 17500 25857 17509 25891
rect 17509 25857 17543 25891
rect 17543 25857 17552 25891
rect 17500 25848 17552 25857
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 18328 25848 18380 25900
rect 19156 25916 19208 25968
rect 19340 25916 19392 25968
rect 21364 25984 21416 26036
rect 23664 25984 23716 26036
rect 23848 25984 23900 26036
rect 26056 25984 26108 26036
rect 18972 25848 19024 25900
rect 20168 25848 20220 25900
rect 20352 25848 20404 25900
rect 20812 25848 20864 25900
rect 12348 25712 12400 25764
rect 14188 25755 14240 25764
rect 14188 25721 14197 25755
rect 14197 25721 14231 25755
rect 14231 25721 14240 25755
rect 14188 25712 14240 25721
rect 14556 25712 14608 25764
rect 14648 25712 14700 25764
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 11980 25687 12032 25696
rect 11980 25653 11989 25687
rect 11989 25653 12023 25687
rect 12023 25653 12032 25687
rect 11980 25644 12032 25653
rect 12532 25687 12584 25696
rect 12532 25653 12541 25687
rect 12541 25653 12575 25687
rect 12575 25653 12584 25687
rect 12532 25644 12584 25653
rect 16028 25644 16080 25696
rect 16488 25712 16540 25764
rect 17592 25712 17644 25764
rect 16672 25644 16724 25696
rect 17500 25644 17552 25696
rect 19984 25780 20036 25832
rect 21732 25848 21784 25900
rect 23664 25848 23716 25900
rect 25228 25891 25280 25900
rect 25228 25857 25237 25891
rect 25237 25857 25271 25891
rect 25271 25857 25280 25891
rect 25228 25848 25280 25857
rect 25872 25891 25924 25900
rect 25872 25857 25881 25891
rect 25881 25857 25915 25891
rect 25915 25857 25924 25891
rect 25872 25848 25924 25857
rect 26608 25916 26660 25968
rect 27160 25916 27212 25968
rect 27988 25984 28040 26036
rect 26884 25848 26936 25900
rect 29460 25916 29512 25968
rect 27528 25848 27580 25900
rect 22008 25823 22060 25832
rect 22008 25789 22017 25823
rect 22017 25789 22051 25823
rect 22051 25789 22060 25823
rect 22008 25780 22060 25789
rect 20352 25712 20404 25764
rect 20076 25687 20128 25696
rect 20076 25653 20085 25687
rect 20085 25653 20119 25687
rect 20119 25653 20128 25687
rect 20076 25644 20128 25653
rect 20812 25644 20864 25696
rect 21732 25644 21784 25696
rect 21824 25644 21876 25696
rect 24124 25780 24176 25832
rect 23112 25712 23164 25764
rect 23388 25687 23440 25696
rect 23388 25653 23397 25687
rect 23397 25653 23431 25687
rect 23431 25653 23440 25687
rect 23388 25644 23440 25653
rect 23940 25644 23992 25696
rect 26792 25780 26844 25832
rect 27804 25848 27856 25900
rect 28356 25891 28408 25900
rect 28356 25857 28365 25891
rect 28365 25857 28399 25891
rect 28399 25857 28408 25891
rect 28356 25848 28408 25857
rect 25780 25712 25832 25764
rect 27160 25755 27212 25764
rect 27160 25721 27169 25755
rect 27169 25721 27203 25755
rect 27203 25721 27212 25755
rect 27160 25712 27212 25721
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 12072 25483 12124 25492
rect 12072 25449 12081 25483
rect 12081 25449 12115 25483
rect 12115 25449 12124 25483
rect 12072 25440 12124 25449
rect 12808 25440 12860 25492
rect 13544 25440 13596 25492
rect 13728 25440 13780 25492
rect 16672 25483 16724 25492
rect 16672 25449 16681 25483
rect 16681 25449 16715 25483
rect 16715 25449 16724 25483
rect 16672 25440 16724 25449
rect 11980 25372 12032 25424
rect 14372 25372 14424 25424
rect 14740 25372 14792 25424
rect 15752 25415 15804 25424
rect 15752 25381 15761 25415
rect 15761 25381 15795 25415
rect 15795 25381 15804 25415
rect 15752 25372 15804 25381
rect 17224 25372 17276 25424
rect 13452 25304 13504 25356
rect 18328 25483 18380 25492
rect 18328 25449 18337 25483
rect 18337 25449 18371 25483
rect 18371 25449 18380 25483
rect 18328 25440 18380 25449
rect 19248 25440 19300 25492
rect 18696 25372 18748 25424
rect 18972 25372 19024 25424
rect 19064 25372 19116 25424
rect 20168 25440 20220 25492
rect 21088 25440 21140 25492
rect 22744 25440 22796 25492
rect 23112 25440 23164 25492
rect 23756 25440 23808 25492
rect 24860 25440 24912 25492
rect 26976 25483 27028 25492
rect 10784 25236 10836 25288
rect 17224 25236 17276 25288
rect 17316 25236 17368 25288
rect 19800 25304 19852 25356
rect 24860 25304 24912 25356
rect 26976 25449 26985 25483
rect 26985 25449 27019 25483
rect 27019 25449 27028 25483
rect 26976 25440 27028 25449
rect 28356 25372 28408 25424
rect 26240 25304 26292 25356
rect 15936 25211 15988 25220
rect 12532 25100 12584 25152
rect 13176 25100 13228 25152
rect 14004 25100 14056 25152
rect 14740 25143 14792 25152
rect 14740 25109 14749 25143
rect 14749 25109 14783 25143
rect 14783 25109 14792 25143
rect 14740 25100 14792 25109
rect 15936 25177 15945 25211
rect 15945 25177 15979 25211
rect 15979 25177 15988 25211
rect 15936 25168 15988 25177
rect 16212 25168 16264 25220
rect 16304 25100 16356 25152
rect 17684 25168 17736 25220
rect 17868 25279 17920 25288
rect 17868 25245 17877 25279
rect 17877 25245 17911 25279
rect 17911 25245 17920 25279
rect 17868 25236 17920 25245
rect 18236 25236 18288 25288
rect 18604 25245 18613 25266
rect 18613 25245 18647 25266
rect 18647 25245 18656 25266
rect 18604 25214 18656 25245
rect 18696 25236 18748 25288
rect 18972 25236 19024 25288
rect 19524 25236 19576 25288
rect 19800 25168 19852 25220
rect 19984 25168 20036 25220
rect 21824 25236 21876 25288
rect 22100 25236 22152 25288
rect 22744 25236 22796 25288
rect 23296 25279 23348 25288
rect 23296 25245 23305 25279
rect 23305 25245 23339 25279
rect 23339 25245 23348 25279
rect 23296 25236 23348 25245
rect 20720 25168 20772 25220
rect 19064 25100 19116 25152
rect 19432 25100 19484 25152
rect 23020 25168 23072 25220
rect 23296 25100 23348 25152
rect 23664 25236 23716 25288
rect 24400 25236 24452 25288
rect 25964 25279 26016 25288
rect 25964 25245 25973 25279
rect 25973 25245 26007 25279
rect 26007 25245 26016 25279
rect 25964 25236 26016 25245
rect 27344 25304 27396 25356
rect 27712 25304 27764 25356
rect 27620 25279 27672 25288
rect 25136 25168 25188 25220
rect 26608 25168 26660 25220
rect 23480 25100 23532 25152
rect 24952 25100 25004 25152
rect 27620 25245 27629 25279
rect 27629 25245 27663 25279
rect 27663 25245 27672 25279
rect 27620 25236 27672 25245
rect 27804 25236 27856 25288
rect 27988 25236 28040 25288
rect 27160 25100 27212 25152
rect 27528 25168 27580 25220
rect 27804 25143 27856 25152
rect 27804 25109 27813 25143
rect 27813 25109 27847 25143
rect 27847 25109 27856 25143
rect 27804 25100 27856 25109
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 17224 24896 17276 24948
rect 13820 24828 13872 24880
rect 16212 24871 16264 24880
rect 16212 24837 16221 24871
rect 16221 24837 16255 24871
rect 16255 24837 16264 24871
rect 16212 24828 16264 24837
rect 18052 24828 18104 24880
rect 18328 24896 18380 24948
rect 19524 24896 19576 24948
rect 21272 24896 21324 24948
rect 25964 24896 26016 24948
rect 27068 24896 27120 24948
rect 13360 24803 13412 24812
rect 13360 24769 13369 24803
rect 13369 24769 13403 24803
rect 13403 24769 13412 24803
rect 13360 24760 13412 24769
rect 13912 24760 13964 24812
rect 15200 24760 15252 24812
rect 16304 24760 16356 24812
rect 18236 24760 18288 24812
rect 18880 24760 18932 24812
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 15200 24624 15252 24676
rect 15384 24624 15436 24676
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 16672 24556 16724 24608
rect 17224 24556 17276 24608
rect 17776 24556 17828 24608
rect 18512 24692 18564 24744
rect 18236 24624 18288 24676
rect 18696 24624 18748 24676
rect 19340 24803 19392 24812
rect 19340 24769 19349 24803
rect 19349 24769 19383 24803
rect 19383 24769 19392 24803
rect 19708 24828 19760 24880
rect 19340 24760 19392 24769
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 21364 24828 21416 24880
rect 22468 24828 22520 24880
rect 22744 24828 22796 24880
rect 23204 24828 23256 24880
rect 22376 24760 22428 24812
rect 23296 24760 23348 24812
rect 25596 24828 25648 24880
rect 24952 24803 25004 24812
rect 24952 24769 24970 24803
rect 24970 24769 25004 24803
rect 25228 24803 25280 24812
rect 24952 24760 25004 24769
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 26148 24828 26200 24880
rect 26516 24828 26568 24880
rect 26700 24828 26752 24880
rect 27528 24871 27580 24880
rect 27528 24837 27537 24871
rect 27537 24837 27571 24871
rect 27571 24837 27580 24871
rect 27528 24828 27580 24837
rect 19984 24624 20036 24676
rect 18328 24556 18380 24608
rect 19340 24556 19392 24608
rect 26884 24760 26936 24812
rect 27804 24760 27856 24812
rect 26976 24692 27028 24744
rect 27436 24692 27488 24744
rect 21456 24556 21508 24608
rect 22192 24556 22244 24608
rect 22376 24556 22428 24608
rect 25964 24624 26016 24676
rect 26332 24624 26384 24676
rect 23204 24556 23256 24608
rect 23388 24556 23440 24608
rect 24584 24556 24636 24608
rect 26056 24556 26108 24608
rect 27160 24599 27212 24608
rect 27160 24565 27169 24599
rect 27169 24565 27203 24599
rect 27203 24565 27212 24599
rect 27160 24556 27212 24565
rect 27252 24556 27304 24608
rect 27436 24556 27488 24608
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 14740 24352 14792 24404
rect 13268 24284 13320 24336
rect 16764 24284 16816 24336
rect 14004 24216 14056 24268
rect 16672 24216 16724 24268
rect 17132 24352 17184 24404
rect 17224 24284 17276 24336
rect 17316 24216 17368 24268
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 16212 24148 16264 24200
rect 17224 24148 17276 24200
rect 14280 24080 14332 24132
rect 18604 24352 18656 24404
rect 19708 24352 19760 24404
rect 23112 24352 23164 24404
rect 23572 24352 23624 24404
rect 24860 24352 24912 24404
rect 19064 24284 19116 24336
rect 19892 24284 19944 24336
rect 20260 24327 20312 24336
rect 20260 24293 20269 24327
rect 20269 24293 20303 24327
rect 20303 24293 20312 24327
rect 20260 24284 20312 24293
rect 20352 24284 20404 24336
rect 21180 24284 21232 24336
rect 22836 24284 22888 24336
rect 22928 24284 22980 24336
rect 26792 24395 26844 24404
rect 26792 24361 26801 24395
rect 26801 24361 26835 24395
rect 26835 24361 26844 24395
rect 26792 24352 26844 24361
rect 27068 24352 27120 24404
rect 27804 24352 27856 24404
rect 18052 24123 18104 24132
rect 18052 24089 18069 24123
rect 18069 24089 18104 24123
rect 19892 24148 19944 24200
rect 20076 24148 20128 24200
rect 20720 24191 20772 24200
rect 18052 24080 18104 24089
rect 16764 24012 16816 24064
rect 19064 24012 19116 24064
rect 20168 24080 20220 24132
rect 20720 24157 20729 24191
rect 20729 24157 20763 24191
rect 20763 24157 20772 24191
rect 20720 24148 20772 24157
rect 20812 24191 20864 24200
rect 20812 24157 20821 24191
rect 20821 24157 20855 24191
rect 20855 24157 20864 24191
rect 21272 24191 21324 24200
rect 20812 24148 20864 24157
rect 21272 24157 21281 24191
rect 21281 24157 21315 24191
rect 21315 24157 21324 24191
rect 21272 24148 21324 24157
rect 23020 24216 23072 24268
rect 20628 24080 20680 24132
rect 21180 24080 21232 24132
rect 21640 24080 21692 24132
rect 23572 24148 23624 24200
rect 24308 24148 24360 24200
rect 27988 24284 28040 24336
rect 24952 24216 25004 24268
rect 25964 24191 26016 24200
rect 19524 24012 19576 24064
rect 19800 24012 19852 24064
rect 19892 24012 19944 24064
rect 23480 24012 23532 24064
rect 25596 24080 25648 24132
rect 25964 24157 25973 24191
rect 25973 24157 26007 24191
rect 26007 24157 26016 24191
rect 25964 24148 26016 24157
rect 26332 24148 26384 24200
rect 27528 24148 27580 24200
rect 26424 24123 26476 24132
rect 26424 24089 26433 24123
rect 26433 24089 26467 24123
rect 26467 24089 26476 24123
rect 26424 24080 26476 24089
rect 26516 24080 26568 24132
rect 27804 24080 27856 24132
rect 28264 24123 28316 24132
rect 28264 24089 28273 24123
rect 28273 24089 28307 24123
rect 28307 24089 28316 24123
rect 28264 24080 28316 24089
rect 26240 24012 26292 24064
rect 26332 24012 26384 24064
rect 26792 24012 26844 24064
rect 27620 24012 27672 24064
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 16396 23808 16448 23860
rect 17316 23808 17368 23860
rect 18696 23808 18748 23860
rect 19156 23808 19208 23860
rect 20812 23808 20864 23860
rect 12716 23740 12768 23792
rect 17132 23740 17184 23792
rect 17960 23740 18012 23792
rect 18788 23740 18840 23792
rect 19064 23740 19116 23792
rect 19432 23740 19484 23792
rect 20168 23740 20220 23792
rect 20352 23740 20404 23792
rect 23572 23808 23624 23860
rect 9772 23672 9824 23724
rect 16672 23672 16724 23724
rect 16948 23672 17000 23724
rect 19984 23715 20036 23724
rect 14188 23604 14240 23656
rect 19524 23604 19576 23656
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 16028 23468 16080 23520
rect 19984 23681 19993 23715
rect 19993 23681 20027 23715
rect 20027 23681 20036 23715
rect 19984 23672 20036 23681
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 20628 23672 20680 23724
rect 20904 23672 20956 23724
rect 21180 23715 21232 23724
rect 21180 23681 21189 23715
rect 21189 23681 21223 23715
rect 21223 23681 21232 23715
rect 21364 23715 21416 23724
rect 21180 23672 21232 23681
rect 21364 23681 21392 23715
rect 21392 23681 21416 23715
rect 21364 23672 21416 23681
rect 21456 23715 21508 23724
rect 21456 23681 21465 23715
rect 21465 23681 21499 23715
rect 21499 23681 21508 23715
rect 23848 23740 23900 23792
rect 21456 23672 21508 23681
rect 19892 23604 19944 23656
rect 21548 23604 21600 23656
rect 17776 23468 17828 23520
rect 17960 23468 18012 23520
rect 18604 23468 18656 23520
rect 19892 23468 19944 23520
rect 21916 23672 21968 23724
rect 22560 23672 22612 23724
rect 21732 23604 21784 23656
rect 22008 23647 22060 23656
rect 22008 23613 22017 23647
rect 22017 23613 22051 23647
rect 22051 23613 22060 23647
rect 22008 23604 22060 23613
rect 23480 23604 23532 23656
rect 25504 23808 25556 23860
rect 27528 23808 27580 23860
rect 24860 23740 24912 23792
rect 27436 23740 27488 23792
rect 24584 23672 24636 23724
rect 26240 23672 26292 23724
rect 26976 23672 27028 23724
rect 27620 23672 27672 23724
rect 28172 23740 28224 23792
rect 28356 23715 28408 23724
rect 28356 23681 28365 23715
rect 28365 23681 28399 23715
rect 28399 23681 28408 23715
rect 28356 23672 28408 23681
rect 28172 23604 28224 23656
rect 23848 23511 23900 23520
rect 23848 23477 23857 23511
rect 23857 23477 23891 23511
rect 23891 23477 23900 23511
rect 27068 23536 27120 23588
rect 23848 23468 23900 23477
rect 26608 23468 26660 23520
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 16304 23264 16356 23316
rect 16764 23307 16816 23316
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 16764 23264 16816 23273
rect 17960 23264 18012 23316
rect 19340 23264 19392 23316
rect 20260 23264 20312 23316
rect 20536 23307 20588 23316
rect 20536 23273 20570 23307
rect 20570 23273 20588 23307
rect 20536 23264 20588 23273
rect 21824 23264 21876 23316
rect 19800 23196 19852 23248
rect 20168 23196 20220 23248
rect 20444 23196 20496 23248
rect 23756 23264 23808 23316
rect 24124 23264 24176 23316
rect 25044 23264 25096 23316
rect 25228 23264 25280 23316
rect 27160 23264 27212 23316
rect 27712 23307 27764 23316
rect 27712 23273 27721 23307
rect 27721 23273 27755 23307
rect 27755 23273 27764 23307
rect 27712 23264 27764 23273
rect 25688 23196 25740 23248
rect 25872 23196 25924 23248
rect 26792 23196 26844 23248
rect 17592 23128 17644 23180
rect 21272 23128 21324 23180
rect 18052 23060 18104 23112
rect 18144 22992 18196 23044
rect 20904 23060 20956 23112
rect 21916 23128 21968 23180
rect 20720 22992 20772 23044
rect 17316 22967 17368 22976
rect 17316 22933 17325 22967
rect 17325 22933 17359 22967
rect 17359 22933 17368 22967
rect 17316 22924 17368 22933
rect 19524 22967 19576 22976
rect 19524 22933 19533 22967
rect 19533 22933 19567 22967
rect 19567 22933 19576 22967
rect 19524 22924 19576 22933
rect 19984 22924 20036 22976
rect 20168 22924 20220 22976
rect 20444 22924 20496 22976
rect 20812 22924 20864 22976
rect 21180 22992 21232 23044
rect 22192 23060 22244 23112
rect 23848 23060 23900 23112
rect 26240 23103 26292 23112
rect 21824 22992 21876 23044
rect 24492 22992 24544 23044
rect 24676 22992 24728 23044
rect 23112 22924 23164 22976
rect 23204 22924 23256 22976
rect 25412 23035 25464 23044
rect 25412 23001 25421 23035
rect 25421 23001 25455 23035
rect 25455 23001 25464 23035
rect 25412 22992 25464 23001
rect 25504 22992 25556 23044
rect 24952 22967 25004 22976
rect 24952 22933 24961 22967
rect 24961 22933 24995 22967
rect 24995 22933 25004 22967
rect 26240 23069 26249 23103
rect 26249 23069 26283 23103
rect 26283 23069 26292 23103
rect 26240 23060 26292 23069
rect 26608 23060 26660 23112
rect 27068 23103 27120 23112
rect 27068 23069 27077 23103
rect 27077 23069 27111 23103
rect 27111 23069 27120 23103
rect 27068 23060 27120 23069
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 24952 22924 25004 22933
rect 26424 22924 26476 22976
rect 26884 22967 26936 22976
rect 26884 22933 26893 22967
rect 26893 22933 26927 22967
rect 26927 22933 26936 22967
rect 26884 22924 26936 22933
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 16396 22720 16448 22772
rect 17224 22720 17276 22772
rect 18972 22720 19024 22772
rect 19800 22763 19852 22772
rect 19800 22729 19809 22763
rect 19809 22729 19843 22763
rect 19843 22729 19852 22763
rect 19800 22720 19852 22729
rect 20260 22720 20312 22772
rect 20904 22720 20956 22772
rect 22100 22720 22152 22772
rect 19892 22652 19944 22704
rect 20444 22695 20496 22704
rect 20444 22661 20471 22695
rect 20471 22661 20496 22695
rect 20444 22652 20496 22661
rect 20720 22652 20772 22704
rect 21088 22695 21140 22704
rect 21088 22661 21097 22695
rect 21097 22661 21131 22695
rect 21131 22661 21140 22695
rect 21088 22652 21140 22661
rect 21824 22584 21876 22636
rect 17500 22516 17552 22568
rect 22468 22720 22520 22772
rect 24216 22763 24268 22772
rect 24216 22729 24243 22763
rect 24243 22729 24268 22763
rect 24216 22720 24268 22729
rect 25780 22763 25832 22772
rect 22284 22627 22336 22670
rect 23112 22652 23164 22704
rect 24308 22652 24360 22704
rect 25780 22729 25789 22763
rect 25789 22729 25823 22763
rect 25823 22729 25832 22763
rect 25780 22720 25832 22729
rect 26240 22720 26292 22772
rect 26792 22720 26844 22772
rect 28172 22763 28224 22772
rect 28172 22729 28181 22763
rect 28181 22729 28215 22763
rect 28215 22729 28224 22763
rect 28172 22720 28224 22729
rect 22284 22618 22301 22627
rect 22301 22618 22335 22627
rect 22335 22618 22336 22627
rect 22836 22584 22888 22636
rect 23020 22627 23072 22636
rect 23020 22593 23029 22627
rect 23029 22593 23063 22627
rect 23063 22593 23072 22627
rect 23020 22584 23072 22593
rect 23572 22627 23624 22636
rect 15476 22448 15528 22500
rect 22928 22516 22980 22568
rect 23572 22593 23581 22627
rect 23581 22593 23615 22627
rect 23615 22593 23624 22627
rect 23572 22584 23624 22593
rect 23940 22584 23992 22636
rect 25504 22652 25556 22704
rect 26700 22652 26752 22704
rect 26884 22584 26936 22636
rect 27896 22584 27948 22636
rect 28264 22584 28316 22636
rect 23848 22516 23900 22568
rect 24952 22516 25004 22568
rect 25596 22516 25648 22568
rect 28632 22516 28684 22568
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 16672 22380 16724 22432
rect 20076 22380 20128 22432
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 21364 22380 21416 22432
rect 22284 22380 22336 22432
rect 25780 22380 25832 22432
rect 27160 22380 27212 22432
rect 27252 22380 27304 22432
rect 29368 22380 29420 22432
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 20444 22176 20496 22228
rect 22284 22176 22336 22228
rect 19892 22108 19944 22160
rect 19984 22108 20036 22160
rect 20168 22151 20220 22160
rect 20168 22117 20177 22151
rect 20177 22117 20211 22151
rect 20211 22117 20220 22151
rect 20168 22108 20220 22117
rect 20260 22108 20312 22160
rect 23020 22219 23072 22228
rect 23020 22185 23029 22219
rect 23029 22185 23063 22219
rect 23063 22185 23072 22219
rect 23020 22176 23072 22185
rect 24400 22176 24452 22228
rect 25872 22176 25924 22228
rect 26148 22176 26200 22228
rect 27344 22176 27396 22228
rect 19800 22040 19852 22092
rect 21364 22040 21416 22092
rect 23388 22108 23440 22160
rect 28540 22108 28592 22160
rect 24124 22040 24176 22092
rect 15936 21972 15988 22024
rect 20260 21972 20312 22024
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 17408 21904 17460 21956
rect 20812 21904 20864 21956
rect 22468 21904 22520 21956
rect 22652 21947 22704 21956
rect 22652 21913 22661 21947
rect 22661 21913 22695 21947
rect 22695 21913 22704 21947
rect 22652 21904 22704 21913
rect 27344 21972 27396 22024
rect 27528 21972 27580 22024
rect 27712 22015 27764 22024
rect 27712 21981 27721 22015
rect 27721 21981 27755 22015
rect 27755 21981 27764 22015
rect 27712 21972 27764 21981
rect 28356 22015 28408 22024
rect 28356 21981 28365 22015
rect 28365 21981 28399 22015
rect 28399 21981 28408 22015
rect 28356 21972 28408 21981
rect 22376 21836 22428 21888
rect 22744 21836 22796 21888
rect 23020 21904 23072 21956
rect 23388 21836 23440 21888
rect 24492 21836 24544 21888
rect 24676 21879 24728 21888
rect 24676 21845 24685 21879
rect 24685 21845 24719 21879
rect 24719 21845 24728 21879
rect 24676 21836 24728 21845
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 19432 21632 19484 21684
rect 21456 21632 21508 21684
rect 24400 21632 24452 21684
rect 25964 21632 26016 21684
rect 18696 21564 18748 21616
rect 21180 21564 21232 21616
rect 21272 21564 21324 21616
rect 22468 21607 22520 21616
rect 22468 21573 22477 21607
rect 22477 21573 22511 21607
rect 22511 21573 22520 21607
rect 22468 21564 22520 21573
rect 23296 21607 23348 21616
rect 23296 21573 23305 21607
rect 23305 21573 23339 21607
rect 23339 21573 23348 21607
rect 23296 21564 23348 21573
rect 23756 21539 23808 21548
rect 23756 21505 23765 21539
rect 23765 21505 23799 21539
rect 23799 21505 23808 21539
rect 23756 21496 23808 21505
rect 1584 21471 1636 21480
rect 1584 21437 1593 21471
rect 1593 21437 1627 21471
rect 1627 21437 1636 21471
rect 1584 21428 1636 21437
rect 12348 21428 12400 21480
rect 24492 21564 24544 21616
rect 25136 21607 25188 21616
rect 25136 21573 25145 21607
rect 25145 21573 25179 21607
rect 25179 21573 25188 21607
rect 25136 21564 25188 21573
rect 26148 21564 26200 21616
rect 26332 21564 26384 21616
rect 24032 21496 24084 21548
rect 27252 21564 27304 21616
rect 28080 21496 28132 21548
rect 19064 21360 19116 21412
rect 18788 21335 18840 21344
rect 18788 21301 18797 21335
rect 18797 21301 18831 21335
rect 18831 21301 18840 21335
rect 18788 21292 18840 21301
rect 20444 21360 20496 21412
rect 24216 21428 24268 21480
rect 20904 21292 20956 21344
rect 21364 21335 21416 21344
rect 21364 21301 21373 21335
rect 21373 21301 21407 21335
rect 21407 21301 21416 21335
rect 21364 21292 21416 21301
rect 21456 21292 21508 21344
rect 22376 21292 22428 21344
rect 22652 21292 22704 21344
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 20352 21088 20404 21140
rect 20444 21131 20496 21140
rect 20444 21097 20453 21131
rect 20453 21097 20487 21131
rect 20487 21097 20496 21131
rect 20444 21088 20496 21097
rect 20812 21088 20864 21140
rect 21364 21088 21416 21140
rect 24860 21088 24912 21140
rect 25136 21131 25188 21140
rect 25136 21097 25145 21131
rect 25145 21097 25179 21131
rect 25179 21097 25188 21131
rect 25136 21088 25188 21097
rect 25780 21131 25832 21140
rect 25780 21097 25789 21131
rect 25789 21097 25823 21131
rect 25823 21097 25832 21131
rect 25780 21088 25832 21097
rect 26332 21088 26384 21140
rect 29184 21088 29236 21140
rect 18788 21020 18840 21072
rect 19524 21020 19576 21072
rect 21088 21020 21140 21072
rect 22376 21020 22428 21072
rect 23756 21063 23808 21072
rect 23756 21029 23765 21063
rect 23765 21029 23799 21063
rect 23799 21029 23808 21063
rect 23756 21020 23808 21029
rect 24216 21020 24268 21072
rect 24768 21020 24820 21072
rect 20536 20884 20588 20936
rect 24676 20952 24728 21004
rect 24860 20952 24912 21004
rect 28448 21020 28500 21072
rect 29276 20952 29328 21004
rect 22652 20884 22704 20936
rect 23020 20884 23072 20936
rect 24584 20884 24636 20936
rect 22560 20859 22612 20868
rect 22560 20825 22569 20859
rect 22569 20825 22603 20859
rect 22603 20825 22612 20859
rect 22560 20816 22612 20825
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 19984 20587 20036 20596
rect 19984 20553 19993 20587
rect 19993 20553 20027 20587
rect 20027 20553 20036 20587
rect 19984 20544 20036 20553
rect 20996 20587 21048 20596
rect 20996 20553 21005 20587
rect 21005 20553 21039 20587
rect 21039 20553 21048 20587
rect 20996 20544 21048 20553
rect 22468 20544 22520 20596
rect 22652 20587 22704 20596
rect 22652 20553 22661 20587
rect 22661 20553 22695 20587
rect 22695 20553 22704 20587
rect 22652 20544 22704 20553
rect 22928 20544 22980 20596
rect 24768 20544 24820 20596
rect 20260 20476 20312 20528
rect 22376 20476 22428 20528
rect 23112 20476 23164 20528
rect 24860 20476 24912 20528
rect 20076 20408 20128 20460
rect 22836 20408 22888 20460
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 26424 20544 26476 20596
rect 27252 20587 27304 20596
rect 27252 20553 27261 20587
rect 27261 20553 27295 20587
rect 27295 20553 27304 20587
rect 27252 20544 27304 20553
rect 29460 20544 29512 20596
rect 28356 20451 28408 20460
rect 28356 20417 28365 20451
rect 28365 20417 28399 20451
rect 28399 20417 28408 20451
rect 28356 20408 28408 20417
rect 25964 20204 26016 20256
rect 26332 20204 26384 20256
rect 26976 20204 27028 20256
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 20628 20043 20680 20052
rect 20628 20009 20637 20043
rect 20637 20009 20671 20043
rect 20671 20009 20680 20043
rect 20628 20000 20680 20009
rect 21640 20043 21692 20052
rect 21640 20009 21649 20043
rect 21649 20009 21683 20043
rect 21683 20009 21692 20043
rect 21640 20000 21692 20009
rect 22284 20043 22336 20052
rect 22284 20009 22293 20043
rect 22293 20009 22327 20043
rect 22327 20009 22336 20043
rect 22284 20000 22336 20009
rect 23756 20000 23808 20052
rect 24124 20000 24176 20052
rect 27528 20000 27580 20052
rect 28356 20000 28408 20052
rect 25780 19932 25832 19984
rect 22652 19864 22704 19916
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 28356 19839 28408 19848
rect 28356 19805 28365 19839
rect 28365 19805 28399 19839
rect 28399 19805 28408 19839
rect 28356 19796 28408 19805
rect 25964 19660 26016 19712
rect 26240 19660 26292 19712
rect 27160 19660 27212 19712
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 21640 19456 21692 19508
rect 22652 19456 22704 19508
rect 23664 19456 23716 19508
rect 26148 19499 26200 19508
rect 26148 19465 26157 19499
rect 26157 19465 26191 19499
rect 26191 19465 26200 19499
rect 26148 19456 26200 19465
rect 28264 19456 28316 19508
rect 26056 19388 26108 19440
rect 24860 19184 24912 19236
rect 28356 19159 28408 19168
rect 28356 19125 28365 19159
rect 28365 19125 28399 19159
rect 28399 19125 28408 19159
rect 28356 19116 28408 19125
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 23572 18955 23624 18964
rect 23572 18921 23581 18955
rect 23581 18921 23615 18955
rect 23615 18921 23624 18955
rect 23572 18912 23624 18921
rect 24952 18912 25004 18964
rect 23756 18844 23808 18896
rect 23572 18776 23624 18828
rect 28356 18751 28408 18760
rect 28356 18717 28365 18751
rect 28365 18717 28399 18751
rect 28399 18717 28408 18751
rect 28356 18708 28408 18717
rect 22376 18615 22428 18624
rect 22376 18581 22385 18615
rect 22385 18581 22419 18615
rect 22419 18581 22428 18615
rect 22376 18572 22428 18581
rect 22468 18572 22520 18624
rect 25688 18572 25740 18624
rect 26884 18615 26936 18624
rect 26884 18581 26893 18615
rect 26893 18581 26927 18615
rect 26927 18581 26936 18615
rect 26884 18572 26936 18581
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 23664 18368 23716 18420
rect 25044 18368 25096 18420
rect 26516 18411 26568 18420
rect 26516 18377 26525 18411
rect 26525 18377 26559 18411
rect 26559 18377 26568 18411
rect 26516 18368 26568 18377
rect 27620 18368 27672 18420
rect 21088 18300 21140 18352
rect 25964 18300 26016 18352
rect 28356 18343 28408 18352
rect 28356 18309 28365 18343
rect 28365 18309 28399 18343
rect 28399 18309 28408 18343
rect 28356 18300 28408 18309
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 24860 18071 24912 18080
rect 24860 18037 24869 18071
rect 24869 18037 24903 18071
rect 24903 18037 24912 18071
rect 24860 18028 24912 18037
rect 25688 18028 25740 18080
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 22744 17824 22796 17876
rect 25596 17867 25648 17876
rect 25596 17833 25605 17867
rect 25605 17833 25639 17867
rect 25639 17833 25648 17867
rect 25596 17824 25648 17833
rect 25780 17824 25832 17876
rect 26976 17867 27028 17876
rect 26976 17833 26985 17867
rect 26985 17833 27019 17867
rect 27019 17833 27028 17867
rect 26976 17824 27028 17833
rect 27804 17824 27856 17876
rect 25504 17756 25556 17808
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 25044 17323 25096 17332
rect 25044 17289 25053 17323
rect 25053 17289 25087 17323
rect 25087 17289 25096 17323
rect 25044 17280 25096 17289
rect 25504 17323 25556 17332
rect 25504 17289 25513 17323
rect 25513 17289 25547 17323
rect 25547 17289 25556 17323
rect 25504 17280 25556 17289
rect 27160 17323 27212 17332
rect 27160 17289 27169 17323
rect 27169 17289 27203 17323
rect 27203 17289 27212 17323
rect 27160 17280 27212 17289
rect 23572 17212 23624 17264
rect 28356 16983 28408 16992
rect 28356 16949 28365 16983
rect 28365 16949 28399 16983
rect 28399 16949 28408 16983
rect 28356 16940 28408 16949
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 24860 16736 24912 16788
rect 26884 16736 26936 16788
rect 25688 16668 25740 16720
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 22376 16192 22428 16244
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 28356 14875 28408 14884
rect 28356 14841 28365 14875
rect 28365 14841 28399 14875
rect 28399 14841 28408 14875
rect 28356 14832 28408 14841
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 28356 13719 28408 13728
rect 28356 13685 28365 13719
rect 28365 13685 28399 13719
rect 28399 13685 28408 13719
rect 28356 13676 28408 13685
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 28356 11543 28408 11552
rect 28356 11509 28365 11543
rect 28365 11509 28399 11543
rect 28399 11509 28408 11543
rect 28356 11500 28408 11509
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 28356 11135 28408 11144
rect 28356 11101 28365 11135
rect 28365 11101 28399 11135
rect 28399 11101 28408 11135
rect 28356 11092 28408 11101
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 28356 9435 28408 9444
rect 28356 9401 28365 9435
rect 28365 9401 28399 9435
rect 28399 9401 28408 9435
rect 28356 9392 28408 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 28356 9095 28408 9104
rect 28356 9061 28365 9095
rect 28365 9061 28399 9095
rect 28399 9061 28408 9095
rect 28356 9052 28408 9061
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 28356 6783 28408 6792
rect 28356 6749 28365 6783
rect 28365 6749 28399 6783
rect 28399 6749 28408 6783
rect 28356 6740 28408 6749
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 28356 5695 28408 5704
rect 28356 5661 28365 5695
rect 28365 5661 28399 5695
rect 28399 5661 28408 5695
rect 28356 5652 28408 5661
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 28356 5015 28408 5024
rect 28356 4981 28365 5015
rect 28365 4981 28399 5015
rect 28399 4981 28408 5015
rect 28356 4972 28408 4981
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 28356 3655 28408 3664
rect 28356 3621 28365 3655
rect 28365 3621 28399 3655
rect 28399 3621 28408 3655
rect 28356 3612 28408 3621
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
<< metal2 >>
rect 570 33200 626 34000
rect 1674 33200 1730 34000
rect 2778 33200 2834 34000
rect 3882 33200 3938 34000
rect 4986 33200 5042 34000
rect 6090 33200 6146 34000
rect 7194 33200 7250 34000
rect 8298 33200 8354 34000
rect 9402 33200 9458 34000
rect 10506 33200 10562 34000
rect 11610 33200 11666 34000
rect 12714 33200 12770 34000
rect 13818 33200 13874 34000
rect 14922 33200 14978 34000
rect 16026 33200 16082 34000
rect 17130 33200 17186 34000
rect 18234 33200 18290 34000
rect 19338 33200 19394 34000
rect 20442 33200 20498 34000
rect 21546 33200 21602 34000
rect 22650 33200 22706 34000
rect 23754 33200 23810 34000
rect 23860 33238 24072 33266
rect 584 31278 612 33200
rect 1688 31482 1716 33200
rect 1676 31476 1728 31482
rect 1676 31418 1728 31424
rect 3896 31346 3924 33200
rect 5000 31482 5028 33200
rect 4988 31476 5040 31482
rect 4988 31418 5040 31424
rect 7208 31346 7236 33200
rect 7896 31580 8204 31589
rect 7896 31578 7902 31580
rect 7958 31578 7982 31580
rect 8038 31578 8062 31580
rect 8118 31578 8142 31580
rect 8198 31578 8204 31580
rect 7958 31526 7960 31578
rect 8140 31526 8142 31578
rect 7896 31524 7902 31526
rect 7958 31524 7982 31526
rect 8038 31524 8062 31526
rect 8118 31524 8142 31526
rect 8198 31524 8204 31526
rect 7896 31515 8204 31524
rect 8312 31482 8340 33200
rect 8392 31952 8444 31958
rect 8392 31894 8444 31900
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 3884 31340 3936 31346
rect 3884 31282 3936 31288
rect 5356 31340 5408 31346
rect 5356 31282 5408 31288
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 572 31272 624 31278
rect 572 31214 624 31220
rect 4423 31036 4731 31045
rect 4423 31034 4429 31036
rect 4485 31034 4509 31036
rect 4565 31034 4589 31036
rect 4645 31034 4669 31036
rect 4725 31034 4731 31036
rect 4485 30982 4487 31034
rect 4667 30982 4669 31034
rect 4423 30980 4429 30982
rect 4485 30980 4509 30982
rect 4565 30980 4589 30982
rect 4645 30980 4669 30982
rect 4725 30980 4731 30982
rect 4423 30971 4731 30980
rect 1584 30728 1636 30734
rect 5368 30705 5396 31282
rect 5816 31136 5868 31142
rect 5816 31078 5868 31084
rect 6184 31136 6236 31142
rect 6184 31078 6236 31084
rect 7656 31136 7708 31142
rect 7656 31078 7708 31084
rect 1584 30670 1636 30676
rect 5354 30696 5410 30705
rect 1596 30297 1624 30670
rect 5354 30631 5410 30640
rect 3424 30592 3476 30598
rect 3424 30534 3476 30540
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 5724 30592 5776 30598
rect 5724 30534 5776 30540
rect 3436 30394 3464 30534
rect 3424 30388 3476 30394
rect 3424 30330 3476 30336
rect 1582 30288 1638 30297
rect 1582 30223 1638 30232
rect 4423 29948 4731 29957
rect 4423 29946 4429 29948
rect 4485 29946 4509 29948
rect 4565 29946 4589 29948
rect 4645 29946 4669 29948
rect 4725 29946 4731 29948
rect 4485 29894 4487 29946
rect 4667 29894 4669 29946
rect 4423 29892 4429 29894
rect 4485 29892 4509 29894
rect 4565 29892 4589 29894
rect 4645 29892 4669 29894
rect 4725 29892 4731 29894
rect 4423 29883 4731 29892
rect 4816 29714 4844 30534
rect 5736 30326 5764 30534
rect 5724 30320 5776 30326
rect 5724 30262 5776 30268
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 5552 29850 5580 30126
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 4804 29708 4856 29714
rect 4804 29650 4856 29656
rect 5736 29646 5764 30262
rect 5828 29850 5856 31078
rect 6196 30938 6224 31078
rect 6184 30932 6236 30938
rect 6184 30874 6236 30880
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 6552 30388 6604 30394
rect 6552 30330 6604 30336
rect 6564 30297 6592 30330
rect 7116 30326 7144 30738
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 7104 30320 7156 30326
rect 6550 30288 6606 30297
rect 7104 30262 7156 30268
rect 6550 30223 6606 30232
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 5816 29844 5868 29850
rect 5816 29786 5868 29792
rect 1584 29640 1636 29646
rect 1582 29608 1584 29617
rect 5724 29640 5776 29646
rect 1636 29608 1638 29617
rect 5724 29582 5776 29588
rect 1582 29543 1638 29552
rect 5264 29504 5316 29510
rect 5264 29446 5316 29452
rect 5276 29306 5304 29446
rect 5264 29300 5316 29306
rect 5264 29242 5316 29248
rect 4423 28860 4731 28869
rect 4423 28858 4429 28860
rect 4485 28858 4509 28860
rect 4565 28858 4589 28860
rect 4645 28858 4669 28860
rect 4725 28858 4731 28860
rect 4485 28806 4487 28858
rect 4667 28806 4669 28858
rect 4423 28804 4429 28806
rect 4485 28804 4509 28806
rect 4565 28804 4589 28806
rect 4645 28804 4669 28806
rect 4725 28804 4731 28806
rect 4423 28795 4731 28804
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1596 28257 1624 28494
rect 1582 28248 1638 28257
rect 1582 28183 1638 28192
rect 6840 28014 6868 29990
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6932 29306 6960 29446
rect 6920 29300 6972 29306
rect 6920 29242 6972 29248
rect 7116 28694 7144 30262
rect 7104 28688 7156 28694
rect 7104 28630 7156 28636
rect 7392 28150 7420 30534
rect 7668 30326 7696 31078
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7656 30320 7708 30326
rect 7656 30262 7708 30268
rect 7760 28694 7788 30874
rect 8404 30734 8432 31894
rect 8576 31748 8628 31754
rect 8576 31690 8628 31696
rect 8484 31408 8536 31414
rect 8484 31350 8536 31356
rect 8496 30938 8524 31350
rect 8588 31346 8616 31690
rect 9864 31408 9916 31414
rect 9864 31350 9916 31356
rect 8576 31340 8628 31346
rect 8576 31282 8628 31288
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 8668 30864 8720 30870
rect 8668 30806 8720 30812
rect 9310 30832 9366 30841
rect 8392 30728 8444 30734
rect 8392 30670 8444 30676
rect 7896 30492 8204 30501
rect 7896 30490 7902 30492
rect 7958 30490 7982 30492
rect 8038 30490 8062 30492
rect 8118 30490 8142 30492
rect 8198 30490 8204 30492
rect 7958 30438 7960 30490
rect 8140 30438 8142 30490
rect 7896 30436 7902 30438
rect 7958 30436 7982 30438
rect 8038 30436 8062 30438
rect 8118 30436 8142 30438
rect 8198 30436 8204 30438
rect 7896 30427 8204 30436
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8312 29850 8340 29990
rect 8300 29844 8352 29850
rect 8300 29786 8352 29792
rect 7896 29404 8204 29413
rect 7896 29402 7902 29404
rect 7958 29402 7982 29404
rect 8038 29402 8062 29404
rect 8118 29402 8142 29404
rect 8198 29402 8204 29404
rect 7958 29350 7960 29402
rect 8140 29350 8142 29402
rect 7896 29348 7902 29350
rect 7958 29348 7982 29350
rect 8038 29348 8062 29350
rect 8118 29348 8142 29350
rect 8198 29348 8204 29350
rect 7896 29339 8204 29348
rect 8404 28762 8432 30670
rect 8484 30660 8536 30666
rect 8484 30602 8536 30608
rect 8496 29850 8524 30602
rect 8680 30598 8708 30806
rect 9310 30767 9366 30776
rect 9324 30734 9352 30767
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 8668 30592 8720 30598
rect 8668 30534 8720 30540
rect 8576 30184 8628 30190
rect 8576 30126 8628 30132
rect 8484 29844 8536 29850
rect 8484 29786 8536 29792
rect 8482 29336 8538 29345
rect 8482 29271 8484 29280
rect 8536 29271 8538 29280
rect 8484 29242 8536 29248
rect 8392 28756 8444 28762
rect 8392 28698 8444 28704
rect 7748 28688 7800 28694
rect 7748 28630 7800 28636
rect 7380 28144 7432 28150
rect 7380 28086 7432 28092
rect 6828 28008 6880 28014
rect 6828 27950 6880 27956
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1596 27577 1624 27814
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 7760 27674 7788 28630
rect 7896 28316 8204 28325
rect 7896 28314 7902 28316
rect 7958 28314 7982 28316
rect 8038 28314 8062 28316
rect 8118 28314 8142 28316
rect 8198 28314 8204 28316
rect 7958 28262 7960 28314
rect 8140 28262 8142 28314
rect 7896 28260 7902 28262
rect 7958 28260 7982 28262
rect 8038 28260 8062 28262
rect 8118 28260 8142 28262
rect 8198 28260 8204 28262
rect 7896 28251 8204 28260
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 8496 27674 8524 27814
rect 7748 27668 7800 27674
rect 7748 27610 7800 27616
rect 8484 27668 8536 27674
rect 8484 27610 8536 27616
rect 1582 27568 1638 27577
rect 1582 27503 1638 27512
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 8312 27033 8340 27270
rect 8298 27024 8354 27033
rect 8298 26959 8354 26968
rect 8588 26926 8616 30126
rect 8680 28762 8708 30534
rect 8944 30320 8996 30326
rect 8944 30262 8996 30268
rect 8760 29300 8812 29306
rect 8760 29242 8812 29248
rect 8772 28966 8800 29242
rect 8956 29034 8984 30262
rect 8944 29028 8996 29034
rect 8944 28970 8996 28976
rect 8760 28960 8812 28966
rect 8760 28902 8812 28908
rect 8668 28756 8720 28762
rect 8668 28698 8720 28704
rect 8956 28558 8984 28970
rect 9220 28960 9272 28966
rect 9220 28902 9272 28908
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 9232 28150 9260 28902
rect 9324 28218 9352 30670
rect 9586 30288 9642 30297
rect 9404 30252 9456 30258
rect 9586 30223 9642 30232
rect 9404 30194 9456 30200
rect 9312 28212 9364 28218
rect 9312 28154 9364 28160
rect 9220 28144 9272 28150
rect 9220 28086 9272 28092
rect 9232 27674 9260 28086
rect 9220 27668 9272 27674
rect 9220 27610 9272 27616
rect 9416 27033 9444 30194
rect 9600 30054 9628 30223
rect 9770 30152 9826 30161
rect 9770 30087 9772 30096
rect 9824 30087 9826 30096
rect 9772 30058 9824 30064
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9634 29844 9686 29850
rect 9634 29786 9686 29792
rect 9646 29696 9674 29786
rect 9770 29744 9826 29753
rect 9646 29688 9770 29696
rect 9646 29679 9826 29688
rect 9646 29668 9812 29679
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9496 29232 9548 29238
rect 9496 29174 9548 29180
rect 9508 28762 9536 29174
rect 9496 28756 9548 28762
rect 9496 28698 9548 28704
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 9508 27130 9536 28562
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9402 27024 9458 27033
rect 9402 26959 9458 26968
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 26217 1624 26318
rect 9600 26234 9628 29514
rect 9876 29492 9904 31350
rect 10140 31136 10192 31142
rect 10140 31078 10192 31084
rect 10048 30660 10100 30666
rect 10048 30602 10100 30608
rect 10060 30433 10088 30602
rect 10046 30424 10102 30433
rect 9956 30388 10008 30394
rect 10152 30394 10180 31078
rect 10046 30359 10102 30368
rect 10140 30388 10192 30394
rect 9956 30330 10008 30336
rect 9968 30122 9996 30330
rect 9956 30116 10008 30122
rect 9956 30058 10008 30064
rect 9956 29504 10008 29510
rect 9876 29464 9956 29492
rect 9956 29446 10008 29452
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 9876 29170 9904 29242
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9678 29064 9734 29073
rect 9678 28999 9734 29008
rect 9692 28490 9720 28999
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9692 27606 9720 28426
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9692 27402 9720 27542
rect 9680 27396 9732 27402
rect 9680 27338 9732 27344
rect 9692 27130 9720 27338
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9772 26784 9824 26790
rect 9876 26772 9904 29106
rect 9824 26744 9904 26772
rect 9772 26726 9824 26732
rect 1582 26208 1638 26217
rect 9600 26206 9720 26234
rect 1582 26143 1638 26152
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 9692 26042 9720 26206
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25537 1624 25638
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 1582 25528 1638 25537
rect 4423 25531 4731 25540
rect 1582 25463 1638 25472
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 1584 24200 1636 24206
rect 1582 24168 1584 24177
rect 1636 24168 1638 24177
rect 1582 24103 1638 24112
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 9784 23730 9812 26726
rect 9864 26376 9916 26382
rect 9862 26344 9864 26353
rect 9968 26364 9996 29446
rect 10060 28218 10088 30359
rect 10140 30330 10192 30336
rect 10520 30190 10548 33200
rect 11624 31482 11652 33200
rect 11796 32224 11848 32230
rect 11796 32166 11848 32172
rect 11704 31816 11756 31822
rect 11704 31758 11756 31764
rect 11612 31476 11664 31482
rect 11612 31418 11664 31424
rect 11150 31376 11206 31385
rect 11150 31311 11152 31320
rect 11204 31311 11206 31320
rect 11152 31282 11204 31288
rect 11369 31036 11677 31045
rect 11369 31034 11375 31036
rect 11431 31034 11455 31036
rect 11511 31034 11535 31036
rect 11591 31034 11615 31036
rect 11671 31034 11677 31036
rect 11431 30982 11433 31034
rect 11613 30982 11615 31034
rect 11369 30980 11375 30982
rect 11431 30980 11455 30982
rect 11511 30980 11535 30982
rect 11591 30980 11615 30982
rect 11671 30980 11677 30982
rect 11369 30971 11677 30980
rect 11244 30932 11296 30938
rect 11244 30874 11296 30880
rect 11152 30660 11204 30666
rect 11152 30602 11204 30608
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10600 30320 10652 30326
rect 10876 30320 10928 30326
rect 10600 30262 10652 30268
rect 10704 30268 10876 30274
rect 10704 30262 10928 30268
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 10324 30116 10376 30122
rect 10324 30058 10376 30064
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10152 29646 10180 29990
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10336 29510 10364 30058
rect 10612 30054 10640 30262
rect 10704 30246 10916 30262
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10324 29504 10376 29510
rect 10324 29446 10376 29452
rect 10140 28552 10192 28558
rect 10140 28494 10192 28500
rect 10152 28218 10180 28494
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 10140 28212 10192 28218
rect 10140 28154 10192 28160
rect 10336 28150 10364 29446
rect 10428 28558 10456 29582
rect 10520 29170 10548 29650
rect 10600 29504 10652 29510
rect 10600 29446 10652 29452
rect 10508 29164 10560 29170
rect 10508 29106 10560 29112
rect 10612 29073 10640 29446
rect 10704 29238 10732 30246
rect 10784 30184 10836 30190
rect 10784 30126 10836 30132
rect 10796 29714 10824 30126
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10784 29708 10836 29714
rect 10784 29650 10836 29656
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10784 29572 10836 29578
rect 10784 29514 10836 29520
rect 10692 29232 10744 29238
rect 10692 29174 10744 29180
rect 10598 29064 10654 29073
rect 10598 28999 10654 29008
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10416 28552 10468 28558
rect 10416 28494 10468 28500
rect 10324 28144 10376 28150
rect 10324 28086 10376 28092
rect 10336 27606 10364 28086
rect 10428 27878 10456 28494
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10416 27872 10468 27878
rect 10416 27814 10468 27820
rect 10520 27606 10548 28154
rect 10612 27878 10640 28902
rect 10600 27872 10652 27878
rect 10600 27814 10652 27820
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 10508 27600 10560 27606
rect 10508 27542 10560 27548
rect 10612 27130 10640 27814
rect 10704 27334 10732 29174
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10600 27124 10652 27130
rect 10600 27066 10652 27072
rect 10612 26586 10640 27066
rect 10704 26586 10732 27270
rect 10600 26580 10652 26586
rect 10600 26522 10652 26528
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 10414 26480 10470 26489
rect 10414 26415 10470 26424
rect 9916 26344 9996 26364
rect 9918 26336 9996 26344
rect 9862 26279 9918 26288
rect 10428 26042 10456 26415
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10612 25906 10640 26522
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10796 25294 10824 29514
rect 10888 28665 10916 29582
rect 10980 28966 11008 29990
rect 11072 29782 11100 30534
rect 11164 30326 11192 30602
rect 11152 30320 11204 30326
rect 11152 30262 11204 30268
rect 11150 30152 11206 30161
rect 11150 30087 11152 30096
rect 11204 30087 11206 30096
rect 11152 30058 11204 30064
rect 11060 29776 11112 29782
rect 11060 29718 11112 29724
rect 11256 29696 11284 30874
rect 11716 30802 11744 31758
rect 11808 31482 11836 32166
rect 13542 31784 13598 31793
rect 13832 31754 13860 33200
rect 14936 32230 14964 33200
rect 14924 32224 14976 32230
rect 14924 32166 14976 32172
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13542 31719 13598 31728
rect 13820 31748 13872 31754
rect 13556 31482 13584 31719
rect 13820 31690 13872 31696
rect 13728 31680 13780 31686
rect 13728 31622 13780 31628
rect 11796 31476 11848 31482
rect 11796 31418 11848 31424
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 13268 31340 13320 31346
rect 13268 31282 13320 31288
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 11992 31249 12020 31282
rect 11978 31240 12034 31249
rect 11978 31175 12034 31184
rect 12164 31136 12216 31142
rect 11978 31104 12034 31113
rect 12164 31078 12216 31084
rect 12716 31136 12768 31142
rect 12716 31078 12768 31084
rect 11978 31039 12034 31048
rect 11796 30932 11848 30938
rect 11796 30874 11848 30880
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 11808 30433 11836 30874
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 11794 30424 11850 30433
rect 11794 30359 11850 30368
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 11369 29948 11677 29957
rect 11369 29946 11375 29948
rect 11431 29946 11455 29948
rect 11511 29946 11535 29948
rect 11591 29946 11615 29948
rect 11671 29946 11677 29948
rect 11431 29894 11433 29946
rect 11613 29894 11615 29946
rect 11369 29892 11375 29894
rect 11431 29892 11455 29894
rect 11511 29892 11535 29894
rect 11591 29892 11615 29894
rect 11671 29892 11677 29894
rect 11369 29883 11677 29892
rect 11612 29776 11664 29782
rect 11164 29668 11284 29696
rect 11334 29744 11390 29753
rect 11612 29718 11664 29724
rect 11334 29679 11336 29688
rect 11060 29640 11112 29646
rect 11060 29582 11112 29588
rect 11072 29034 11100 29582
rect 11060 29028 11112 29034
rect 11060 28970 11112 28976
rect 10968 28960 11020 28966
rect 10968 28902 11020 28908
rect 11164 28762 11192 29668
rect 11388 29679 11390 29688
rect 11336 29650 11388 29656
rect 11244 28960 11296 28966
rect 11624 28948 11652 29718
rect 11716 29209 11744 30194
rect 11900 29730 11928 30738
rect 11992 30598 12020 31039
rect 12070 30968 12126 30977
rect 12070 30903 12126 30912
rect 12084 30666 12112 30903
rect 12072 30660 12124 30666
rect 12072 30602 12124 30608
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 11808 29702 11928 29730
rect 11702 29200 11758 29209
rect 11702 29135 11758 29144
rect 11624 28920 11744 28948
rect 11244 28902 11296 28908
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 10874 28656 10930 28665
rect 10874 28591 10930 28600
rect 11072 28218 11100 28698
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 11164 27130 11192 28698
rect 11256 28626 11284 28902
rect 11369 28860 11677 28869
rect 11369 28858 11375 28860
rect 11431 28858 11455 28860
rect 11511 28858 11535 28860
rect 11591 28858 11615 28860
rect 11671 28858 11677 28860
rect 11431 28806 11433 28858
rect 11613 28806 11615 28858
rect 11369 28804 11375 28806
rect 11431 28804 11455 28806
rect 11511 28804 11535 28806
rect 11591 28804 11615 28806
rect 11671 28804 11677 28806
rect 11369 28795 11677 28804
rect 11612 28756 11664 28762
rect 11612 28698 11664 28704
rect 11244 28620 11296 28626
rect 11244 28562 11296 28568
rect 11428 28484 11480 28490
rect 11428 28426 11480 28432
rect 11440 28121 11468 28426
rect 11426 28112 11482 28121
rect 11426 28047 11482 28056
rect 11624 27946 11652 28698
rect 11716 28393 11744 28920
rect 11808 28490 11836 29702
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11900 29073 11928 29582
rect 11886 29064 11942 29073
rect 11886 28999 11942 29008
rect 11992 28914 12020 30534
rect 12176 30054 12204 31078
rect 12440 30932 12492 30938
rect 12440 30874 12492 30880
rect 12452 30802 12480 30874
rect 12440 30796 12492 30802
rect 12440 30738 12492 30744
rect 12348 30728 12400 30734
rect 12268 30688 12348 30716
rect 12268 30258 12296 30688
rect 12348 30670 12400 30676
rect 12452 30580 12480 30738
rect 12360 30552 12480 30580
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12072 30048 12124 30054
rect 12072 29990 12124 29996
rect 12164 30048 12216 30054
rect 12164 29990 12216 29996
rect 11900 28886 12020 28914
rect 11796 28484 11848 28490
rect 11796 28426 11848 28432
rect 11702 28384 11758 28393
rect 11702 28319 11758 28328
rect 11612 27940 11664 27946
rect 11612 27882 11664 27888
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 11716 27606 11744 28319
rect 11808 28218 11836 28426
rect 11900 28422 11928 28886
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11796 28212 11848 28218
rect 11796 28154 11848 28160
rect 11808 28014 11836 28154
rect 11900 28150 11928 28358
rect 11888 28144 11940 28150
rect 11888 28086 11940 28092
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11704 27600 11756 27606
rect 11704 27542 11756 27548
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 11348 27334 11376 27474
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 11900 27130 11928 28086
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 11888 27124 11940 27130
rect 11888 27066 11940 27072
rect 11164 26518 11192 27066
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 11152 26512 11204 26518
rect 11152 26454 11204 26460
rect 11900 26314 11928 27066
rect 11888 26308 11940 26314
rect 11888 26250 11940 26256
rect 11992 25702 12020 27950
rect 12084 27577 12112 29990
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 12176 29238 12204 29582
rect 12164 29232 12216 29238
rect 12164 29174 12216 29180
rect 12176 28694 12204 29174
rect 12268 29170 12296 30194
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12164 28688 12216 28694
rect 12164 28630 12216 28636
rect 12176 27674 12204 28630
rect 12268 28014 12296 29106
rect 12360 28558 12388 30552
rect 12624 30252 12676 30258
rect 12624 30194 12676 30200
rect 12636 29850 12664 30194
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12544 29730 12572 29786
rect 12728 29730 12756 31078
rect 13280 30938 13308 31282
rect 13372 31113 13400 31282
rect 13740 31278 13768 31622
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13912 31136 13964 31142
rect 13358 31104 13414 31113
rect 13912 31078 13964 31084
rect 13358 31039 13414 31048
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 12808 30116 12860 30122
rect 12808 30058 12860 30064
rect 12544 29702 12756 29730
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 12452 29170 12480 29514
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12624 29164 12676 29170
rect 12624 29106 12676 29112
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12360 28257 12388 28494
rect 12346 28248 12402 28257
rect 12346 28183 12402 28192
rect 12348 28144 12400 28150
rect 12348 28086 12400 28092
rect 12256 28008 12308 28014
rect 12256 27950 12308 27956
rect 12256 27872 12308 27878
rect 12256 27814 12308 27820
rect 12268 27674 12296 27814
rect 12164 27668 12216 27674
rect 12164 27610 12216 27616
rect 12256 27668 12308 27674
rect 12256 27610 12308 27616
rect 12070 27568 12126 27577
rect 12070 27503 12126 27512
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 11992 25430 12020 25638
rect 12084 25498 12112 26522
rect 12176 26042 12204 27610
rect 12360 27062 12388 28086
rect 12452 27441 12480 29106
rect 12532 28552 12584 28558
rect 12530 28520 12532 28529
rect 12584 28520 12586 28529
rect 12530 28455 12586 28464
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12544 27713 12572 28018
rect 12530 27704 12586 27713
rect 12530 27639 12586 27648
rect 12438 27432 12494 27441
rect 12438 27367 12494 27376
rect 12636 27130 12664 29106
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12348 27056 12400 27062
rect 12348 26998 12400 27004
rect 12360 26586 12388 26998
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12348 26444 12400 26450
rect 12624 26444 12676 26450
rect 12400 26404 12624 26432
rect 12348 26386 12400 26392
rect 12624 26386 12676 26392
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 12360 25770 12388 26386
rect 12348 25764 12400 25770
rect 12348 25706 12400 25712
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 11980 25424 12032 25430
rect 11980 25366 12032 25372
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22137 1624 22374
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 12360 21486 12388 25706
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12544 25158 12572 25638
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12728 23798 12756 29702
rect 12820 28994 12848 30058
rect 12912 29481 12940 30262
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 12898 29472 12954 29481
rect 12898 29407 12954 29416
rect 13004 29034 13032 29514
rect 12992 29028 13044 29034
rect 12820 28966 12940 28994
rect 12992 28970 13044 28976
rect 13084 29028 13136 29034
rect 13084 28970 13136 28976
rect 12808 27600 12860 27606
rect 12808 27542 12860 27548
rect 12820 25498 12848 27542
rect 12912 27402 12940 28966
rect 13096 28642 13124 28970
rect 13188 28762 13216 30670
rect 13280 30025 13308 30670
rect 13360 30252 13412 30258
rect 13360 30194 13412 30200
rect 13266 30016 13322 30025
rect 13266 29951 13322 29960
rect 13280 29617 13308 29951
rect 13266 29608 13322 29617
rect 13266 29543 13322 29552
rect 13372 29345 13400 30194
rect 13464 29782 13492 30670
rect 13636 30592 13688 30598
rect 13636 30534 13688 30540
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13358 29336 13414 29345
rect 13358 29271 13414 29280
rect 13176 28756 13228 28762
rect 13176 28698 13228 28704
rect 13266 28656 13322 28665
rect 13096 28614 13216 28642
rect 13084 28416 13136 28422
rect 13084 28358 13136 28364
rect 12990 28248 13046 28257
rect 13096 28218 13124 28358
rect 12990 28183 13046 28192
rect 13084 28212 13136 28218
rect 13004 28082 13032 28183
rect 13084 28154 13136 28160
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12912 25945 12940 27338
rect 13004 26994 13032 28018
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 13004 26761 13032 26930
rect 12990 26752 13046 26761
rect 12990 26687 13046 26696
rect 12898 25936 12954 25945
rect 12898 25871 12954 25880
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 13096 24313 13124 27814
rect 13188 25158 13216 28614
rect 13266 28591 13322 28600
rect 13280 28422 13308 28591
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 13268 28008 13320 28014
rect 13266 27976 13268 27985
rect 13320 27976 13322 27985
rect 13266 27911 13322 27920
rect 13372 27520 13400 29271
rect 13544 29232 13596 29238
rect 13544 29174 13596 29180
rect 13556 28014 13584 29174
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13544 27532 13596 27538
rect 13372 27492 13492 27520
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 13372 27305 13400 27338
rect 13358 27296 13414 27305
rect 13358 27231 13414 27240
rect 13360 26784 13412 26790
rect 13360 26726 13412 26732
rect 13372 26450 13400 26726
rect 13360 26444 13412 26450
rect 13360 26386 13412 26392
rect 13266 26344 13322 26353
rect 13266 26279 13322 26288
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13280 24342 13308 26279
rect 13372 24818 13400 26386
rect 13464 25362 13492 27492
rect 13544 27474 13596 27480
rect 13556 27334 13584 27474
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13556 25974 13584 27270
rect 13648 26994 13676 30534
rect 13728 29776 13780 29782
rect 13728 29718 13780 29724
rect 13740 29617 13768 29718
rect 13726 29608 13782 29617
rect 13726 29543 13782 29552
rect 13820 28620 13872 28626
rect 13820 28562 13872 28568
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13636 26988 13688 26994
rect 13636 26930 13688 26936
rect 13544 25968 13596 25974
rect 13544 25910 13596 25916
rect 13740 25498 13768 28494
rect 13832 28393 13860 28562
rect 13818 28384 13874 28393
rect 13818 28319 13874 28328
rect 13832 27538 13860 28319
rect 13924 27946 13952 31078
rect 14016 30734 14044 31826
rect 16580 31748 16632 31754
rect 16580 31690 16632 31696
rect 14842 31580 15150 31589
rect 14842 31578 14848 31580
rect 14904 31578 14928 31580
rect 14984 31578 15008 31580
rect 15064 31578 15088 31580
rect 15144 31578 15150 31580
rect 14904 31526 14906 31578
rect 15086 31526 15088 31578
rect 14842 31524 14848 31526
rect 14904 31524 14928 31526
rect 14984 31524 15008 31526
rect 15064 31524 15088 31526
rect 15144 31524 15150 31526
rect 14842 31515 15150 31524
rect 15658 31512 15714 31521
rect 15658 31447 15714 31456
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 14004 30728 14056 30734
rect 14004 30670 14056 30676
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 15108 30728 15160 30734
rect 15292 30728 15344 30734
rect 15160 30688 15240 30716
rect 15108 30670 15160 30676
rect 14372 30320 14424 30326
rect 14186 30288 14242 30297
rect 14372 30262 14424 30268
rect 14186 30223 14242 30232
rect 14200 29889 14228 30223
rect 14186 29880 14242 29889
rect 14186 29815 14242 29824
rect 14280 29844 14332 29850
rect 14280 29786 14332 29792
rect 14004 29572 14056 29578
rect 14004 29514 14056 29520
rect 14016 28490 14044 29514
rect 14094 29472 14150 29481
rect 14094 29407 14150 29416
rect 14004 28484 14056 28490
rect 14004 28426 14056 28432
rect 13912 27940 13964 27946
rect 13912 27882 13964 27888
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13832 26994 13860 27338
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 13924 26314 13952 26862
rect 13912 26308 13964 26314
rect 13912 26250 13964 26256
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 13556 24854 13584 25434
rect 13820 24880 13872 24886
rect 13556 24828 13820 24854
rect 13556 24826 13872 24828
rect 13820 24822 13872 24826
rect 13924 24818 13952 26250
rect 14016 25265 14044 28426
rect 14108 27946 14136 29407
rect 14096 27940 14148 27946
rect 14096 27882 14148 27888
rect 14002 25256 14058 25265
rect 14002 25191 14058 25200
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13268 24336 13320 24342
rect 13082 24304 13138 24313
rect 13268 24278 13320 24284
rect 14016 24274 14044 25094
rect 14108 24857 14136 27882
rect 14186 27704 14242 27713
rect 14186 27639 14242 27648
rect 14200 27334 14228 27639
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14200 26586 14228 26726
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 14188 25764 14240 25770
rect 14188 25706 14240 25712
rect 14094 24848 14150 24857
rect 14094 24783 14150 24792
rect 13082 24239 13138 24248
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 14200 23662 14228 25706
rect 14292 24138 14320 29786
rect 14384 27606 14412 30262
rect 14464 30116 14516 30122
rect 14464 30058 14516 30064
rect 14476 29170 14504 30058
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 14462 29064 14518 29073
rect 14462 28999 14518 29008
rect 14476 28966 14504 28999
rect 14464 28960 14516 28966
rect 14464 28902 14516 28908
rect 14568 28694 14596 30670
rect 14648 30592 14700 30598
rect 14648 30534 14700 30540
rect 14660 30326 14688 30534
rect 14842 30492 15150 30501
rect 14842 30490 14848 30492
rect 14904 30490 14928 30492
rect 14984 30490 15008 30492
rect 15064 30490 15088 30492
rect 15144 30490 15150 30492
rect 14904 30438 14906 30490
rect 15086 30438 15088 30490
rect 14842 30436 14848 30438
rect 14904 30436 14928 30438
rect 14984 30436 15008 30438
rect 15064 30436 15088 30438
rect 15144 30436 15150 30438
rect 14842 30427 15150 30436
rect 14648 30320 14700 30326
rect 14648 30262 14700 30268
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 15014 30016 15070 30025
rect 14844 29578 14872 29990
rect 15014 29951 15070 29960
rect 15028 29646 15056 29951
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14832 29572 14884 29578
rect 14832 29514 14884 29520
rect 14648 29504 14700 29510
rect 14648 29446 14700 29452
rect 14556 28688 14608 28694
rect 14556 28630 14608 28636
rect 14568 28558 14596 28630
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14476 27849 14504 27950
rect 14568 27946 14596 28494
rect 14660 28150 14688 29446
rect 14842 29404 15150 29413
rect 14842 29402 14848 29404
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 15144 29402 15150 29404
rect 14904 29350 14906 29402
rect 15086 29350 15088 29402
rect 14842 29348 14848 29350
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 15144 29348 15150 29350
rect 14842 29339 15150 29348
rect 15212 29288 15240 30688
rect 15292 30670 15344 30676
rect 15304 30297 15332 30670
rect 15290 30288 15346 30297
rect 15290 30223 15346 30232
rect 15292 29776 15344 29782
rect 15292 29718 15344 29724
rect 15120 29260 15240 29288
rect 15016 29232 15068 29238
rect 15016 29174 15068 29180
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14752 28082 14780 29038
rect 15028 28694 15056 29174
rect 15016 28688 15068 28694
rect 15016 28630 15068 28636
rect 15120 28558 15148 29260
rect 15304 28937 15332 29718
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15396 29238 15424 29582
rect 15488 29238 15516 31282
rect 15580 29850 15608 31350
rect 15672 30598 15700 31447
rect 16488 31272 16540 31278
rect 16488 31214 16540 31220
rect 16304 30660 16356 30666
rect 16304 30602 16356 30608
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15752 30252 15804 30258
rect 16028 30252 16080 30258
rect 15804 30212 15976 30240
rect 15752 30194 15804 30200
rect 15948 30054 15976 30212
rect 16028 30194 16080 30200
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15568 29844 15620 29850
rect 15568 29786 15620 29792
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15476 29232 15528 29238
rect 15476 29174 15528 29180
rect 15290 28928 15346 28937
rect 15290 28863 15346 28872
rect 15476 28688 15528 28694
rect 15476 28630 15528 28636
rect 15292 28620 15344 28626
rect 15292 28562 15344 28568
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 14842 28316 15150 28325
rect 14842 28314 14848 28316
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 15144 28314 15150 28316
rect 14904 28262 14906 28314
rect 15086 28262 15088 28314
rect 14842 28260 14848 28262
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 15144 28260 15150 28262
rect 14842 28251 15150 28260
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14648 28008 14700 28014
rect 14648 27950 14700 27956
rect 14556 27940 14608 27946
rect 14556 27882 14608 27888
rect 14462 27840 14518 27849
rect 14462 27775 14518 27784
rect 14372 27600 14424 27606
rect 14372 27542 14424 27548
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14462 27296 14518 27305
rect 14462 27231 14518 27240
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14384 26897 14412 26998
rect 14370 26888 14426 26897
rect 14370 26823 14426 26832
rect 14372 26512 14424 26518
rect 14372 26454 14424 26460
rect 14384 25430 14412 26454
rect 14372 25424 14424 25430
rect 14372 25366 14424 25372
rect 14476 24177 14504 27231
rect 14568 26790 14596 27474
rect 14556 26784 14608 26790
rect 14556 26726 14608 26732
rect 14568 25770 14596 26726
rect 14660 26518 14688 27950
rect 14752 27674 14780 28018
rect 14832 27940 14884 27946
rect 14832 27882 14884 27888
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 14844 27538 14872 27882
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14832 27532 14884 27538
rect 14832 27474 14884 27480
rect 14936 27470 14964 27814
rect 15198 27704 15254 27713
rect 15304 27690 15332 28562
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15396 28257 15424 28494
rect 15488 28393 15516 28630
rect 15474 28384 15530 28393
rect 15474 28319 15530 28328
rect 15382 28248 15438 28257
rect 15382 28183 15438 28192
rect 15474 27704 15530 27713
rect 15304 27662 15474 27690
rect 15198 27639 15254 27648
rect 15474 27639 15530 27648
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14648 26512 14700 26518
rect 14648 26454 14700 26460
rect 14646 26344 14702 26353
rect 14646 26279 14648 26288
rect 14700 26279 14702 26288
rect 14648 26250 14700 26256
rect 14752 26042 14780 27066
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14844 26761 14872 26930
rect 14830 26752 14886 26761
rect 14830 26687 14886 26696
rect 15106 26616 15162 26625
rect 15106 26551 15162 26560
rect 15120 26382 15148 26551
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 15212 26042 15240 27639
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15304 26994 15332 27406
rect 15382 27296 15438 27305
rect 15382 27231 15438 27240
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 15290 26752 15346 26761
rect 15290 26687 15346 26696
rect 14740 26036 14792 26042
rect 14740 25978 14792 25984
rect 15200 26036 15252 26042
rect 15200 25978 15252 25984
rect 14738 25936 14794 25945
rect 14648 25900 14700 25906
rect 15304 25922 15332 26687
rect 14738 25871 14740 25880
rect 14648 25842 14700 25848
rect 14792 25871 14794 25880
rect 15212 25894 15332 25922
rect 14740 25842 14792 25848
rect 14660 25770 14688 25842
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14648 25764 14700 25770
rect 14648 25706 14700 25712
rect 14740 25424 14792 25430
rect 14740 25366 14792 25372
rect 14752 25158 14780 25366
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14752 24410 14780 25094
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 15212 24818 15240 25894
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15212 24682 15240 24754
rect 15396 24682 15424 27231
rect 15488 27130 15516 27639
rect 15476 27124 15528 27130
rect 15476 27066 15528 27072
rect 15580 27062 15608 29650
rect 15568 27056 15620 27062
rect 15568 26998 15620 27004
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15474 26616 15530 26625
rect 15474 26551 15530 26560
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 14740 24404 14792 24410
rect 14740 24346 14792 24352
rect 14462 24168 14518 24177
rect 14280 24132 14332 24138
rect 14462 24103 14518 24112
rect 14280 24074 14332 24080
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 14188 23656 14240 23662
rect 14188 23598 14240 23604
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 15488 22506 15516 26551
rect 15580 26382 15608 26726
rect 15672 26518 15700 29990
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 15752 29572 15804 29578
rect 15752 29514 15804 29520
rect 15764 29481 15792 29514
rect 15750 29472 15806 29481
rect 15750 29407 15806 29416
rect 15750 29336 15806 29345
rect 15750 29271 15806 29280
rect 15764 29170 15792 29271
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15750 28928 15806 28937
rect 15750 28863 15806 28872
rect 15764 26858 15792 28863
rect 15752 26852 15804 26858
rect 15752 26794 15804 26800
rect 15660 26512 15712 26518
rect 15660 26454 15712 26460
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15672 24614 15700 25774
rect 15764 25430 15792 26794
rect 15856 25974 15884 29786
rect 16040 28200 16068 30194
rect 16210 29880 16266 29889
rect 16210 29815 16266 29824
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 15948 28172 16068 28200
rect 15948 27878 15976 28172
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 16040 27674 16068 28018
rect 16132 28014 16160 28358
rect 16120 28008 16172 28014
rect 16120 27950 16172 27956
rect 15936 27668 15988 27674
rect 15936 27610 15988 27616
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 15948 26761 15976 27610
rect 16028 27532 16080 27538
rect 16028 27474 16080 27480
rect 16040 27305 16068 27474
rect 16120 27396 16172 27402
rect 16120 27338 16172 27344
rect 16026 27296 16082 27305
rect 16026 27231 16082 27240
rect 16132 26994 16160 27338
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16120 26784 16172 26790
rect 15934 26752 15990 26761
rect 16120 26726 16172 26732
rect 15934 26687 15990 26696
rect 16132 26625 16160 26726
rect 15934 26616 15990 26625
rect 15934 26551 15990 26560
rect 16118 26616 16174 26625
rect 16118 26551 16174 26560
rect 15844 25968 15896 25974
rect 15844 25910 15896 25916
rect 15752 25424 15804 25430
rect 15752 25366 15804 25372
rect 15948 25344 15976 26551
rect 16120 26512 16172 26518
rect 16116 26466 16120 26500
rect 16040 26460 16120 26466
rect 16040 26454 16172 26460
rect 16040 26438 16144 26454
rect 16040 25838 16068 26438
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16132 26217 16160 26318
rect 16118 26208 16174 26217
rect 16118 26143 16174 26152
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 16028 25696 16080 25702
rect 16132 25684 16160 26143
rect 16224 26058 16252 29815
rect 16316 28422 16344 30602
rect 16396 30388 16448 30394
rect 16396 30330 16448 30336
rect 16408 29850 16436 30330
rect 16500 30122 16528 31214
rect 16488 30116 16540 30122
rect 16488 30058 16540 30064
rect 16396 29844 16448 29850
rect 16396 29786 16448 29792
rect 16500 29646 16528 30058
rect 16488 29640 16540 29646
rect 16488 29582 16540 29588
rect 16592 29306 16620 31690
rect 17144 31657 17172 33200
rect 18248 31754 18276 33200
rect 20260 32088 20312 32094
rect 20260 32030 20312 32036
rect 18696 31884 18748 31890
rect 18696 31826 18748 31832
rect 18064 31726 18276 31754
rect 17130 31648 17186 31657
rect 17130 31583 17186 31592
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 16776 29345 16804 31282
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16960 30258 16988 31078
rect 17052 30394 17080 31282
rect 17958 30968 18014 30977
rect 17958 30903 18014 30912
rect 17500 30864 17552 30870
rect 17500 30806 17552 30812
rect 17316 30796 17368 30802
rect 17316 30738 17368 30744
rect 17328 30394 17356 30738
rect 17512 30705 17540 30806
rect 17684 30728 17736 30734
rect 17498 30696 17554 30705
rect 17498 30631 17554 30640
rect 17682 30696 17684 30705
rect 17736 30696 17738 30705
rect 17972 30666 18000 30903
rect 17682 30631 17738 30640
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 17868 30592 17920 30598
rect 17868 30534 17920 30540
rect 17590 30424 17646 30433
rect 17040 30388 17092 30394
rect 17040 30330 17092 30336
rect 17316 30388 17368 30394
rect 17368 30348 17448 30376
rect 17646 30368 17658 30410
rect 17590 30359 17658 30368
rect 17316 30330 17368 30336
rect 17130 30288 17186 30297
rect 16948 30252 17000 30258
rect 17130 30223 17186 30232
rect 16948 30194 17000 30200
rect 16856 30184 16908 30190
rect 16856 30126 16908 30132
rect 16762 29336 16818 29345
rect 16580 29300 16632 29306
rect 16762 29271 16818 29280
rect 16580 29242 16632 29248
rect 16764 29232 16816 29238
rect 16764 29174 16816 29180
rect 16776 29034 16804 29174
rect 16764 29028 16816 29034
rect 16764 28970 16816 28976
rect 16396 28960 16448 28966
rect 16396 28902 16448 28908
rect 16488 28960 16540 28966
rect 16488 28902 16540 28908
rect 16304 28416 16356 28422
rect 16304 28358 16356 28364
rect 16304 28144 16356 28150
rect 16304 28086 16356 28092
rect 16316 27674 16344 28086
rect 16304 27668 16356 27674
rect 16304 27610 16356 27616
rect 16302 27160 16358 27169
rect 16302 27095 16358 27104
rect 16316 26858 16344 27095
rect 16304 26852 16356 26858
rect 16304 26794 16356 26800
rect 16316 26246 16344 26794
rect 16408 26296 16436 28902
rect 16500 28393 16528 28902
rect 16764 28688 16816 28694
rect 16764 28630 16816 28636
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 16486 28384 16542 28393
rect 16486 28319 16542 28328
rect 16578 28248 16634 28257
rect 16578 28183 16634 28192
rect 16592 27962 16620 28183
rect 16500 27934 16620 27962
rect 16500 27130 16528 27934
rect 16684 27860 16712 28562
rect 16592 27832 16712 27860
rect 16488 27124 16540 27130
rect 16488 27066 16540 27072
rect 16592 27010 16620 27832
rect 16672 27328 16724 27334
rect 16672 27270 16724 27276
rect 16500 26982 16620 27010
rect 16500 26518 16528 26982
rect 16684 26625 16712 27270
rect 16776 27169 16804 28630
rect 16762 27160 16818 27169
rect 16762 27095 16818 27104
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16776 26790 16804 26862
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16670 26616 16726 26625
rect 16670 26551 16726 26560
rect 16488 26512 16540 26518
rect 16488 26454 16540 26460
rect 16580 26512 16632 26518
rect 16580 26454 16632 26460
rect 16408 26268 16528 26296
rect 16304 26240 16356 26246
rect 16356 26206 16436 26234
rect 16500 26217 16528 26268
rect 16304 26182 16356 26188
rect 16224 26030 16344 26058
rect 16212 25968 16264 25974
rect 16212 25910 16264 25916
rect 16080 25656 16160 25684
rect 16028 25638 16080 25644
rect 15948 25316 16068 25344
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 23633 15700 24550
rect 15658 23624 15714 23633
rect 15658 23559 15714 23568
rect 15476 22500 15528 22506
rect 15476 22442 15528 22448
rect 15948 22030 15976 25162
rect 16040 23526 16068 25316
rect 16132 24041 16160 25656
rect 16224 25226 16252 25910
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 16224 24886 16252 25162
rect 16316 25158 16344 26030
rect 16408 25673 16436 26206
rect 16486 26208 16542 26217
rect 16486 26143 16542 26152
rect 16488 25764 16540 25770
rect 16488 25706 16540 25712
rect 16394 25664 16450 25673
rect 16394 25599 16450 25608
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 16224 24206 16252 24822
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16118 24032 16174 24041
rect 16118 23967 16174 23976
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 16316 23322 16344 24754
rect 16408 23866 16436 25599
rect 16500 24585 16528 25706
rect 16592 24721 16620 26454
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16684 26042 16712 26318
rect 16762 26072 16818 26081
rect 16672 26036 16724 26042
rect 16762 26007 16818 26016
rect 16672 25978 16724 25984
rect 16684 25786 16712 25978
rect 16776 25974 16804 26007
rect 16764 25968 16816 25974
rect 16868 25945 16896 30126
rect 17144 29889 17172 30223
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17130 29880 17186 29889
rect 17130 29815 17186 29824
rect 17040 29776 17092 29782
rect 17040 29718 17092 29724
rect 16948 29504 17000 29510
rect 16948 29446 17000 29452
rect 16960 29102 16988 29446
rect 16948 29096 17000 29102
rect 17052 29073 17080 29718
rect 16948 29038 17000 29044
rect 17038 29064 17094 29073
rect 17038 28999 17094 29008
rect 17040 28008 17092 28014
rect 17092 27956 17172 27962
rect 17040 27950 17172 27956
rect 17052 27934 17172 27950
rect 17040 27872 17092 27878
rect 17040 27814 17092 27820
rect 16948 27396 17000 27402
rect 16948 27338 17000 27344
rect 16764 25910 16816 25916
rect 16854 25936 16910 25945
rect 16854 25871 16910 25880
rect 16684 25758 16804 25786
rect 16672 25696 16724 25702
rect 16672 25638 16724 25644
rect 16684 25498 16712 25638
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16578 24712 16634 24721
rect 16578 24647 16634 24656
rect 16486 24576 16542 24585
rect 16486 24511 16542 24520
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16408 22778 16436 23802
rect 16592 23712 16620 24647
rect 16684 24614 16712 25434
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16776 24426 16804 25758
rect 16684 24398 16804 24426
rect 16684 24274 16712 24398
rect 16764 24336 16816 24342
rect 16764 24278 16816 24284
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 16776 24070 16804 24278
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 16672 23724 16724 23730
rect 16592 23684 16672 23712
rect 16672 23666 16724 23672
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16684 22438 16712 23666
rect 16776 23322 16804 24006
rect 16960 23730 16988 27338
rect 17052 23769 17080 27814
rect 17144 27606 17172 27934
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 17132 27396 17184 27402
rect 17132 27338 17184 27344
rect 17144 26518 17172 27338
rect 17132 26512 17184 26518
rect 17132 26454 17184 26460
rect 17236 26081 17264 30126
rect 17314 29880 17370 29889
rect 17314 29815 17370 29824
rect 17328 29714 17356 29815
rect 17316 29708 17368 29714
rect 17316 29650 17368 29656
rect 17420 29646 17448 30348
rect 17630 30308 17658 30359
rect 17630 30280 17724 30308
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17512 29170 17540 30194
rect 17316 29164 17368 29170
rect 17316 29106 17368 29112
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17222 26072 17278 26081
rect 17222 26007 17278 26016
rect 17328 25922 17356 29106
rect 17406 29064 17462 29073
rect 17406 28999 17462 29008
rect 17420 27305 17448 28999
rect 17512 28014 17540 29106
rect 17592 28484 17644 28490
rect 17592 28426 17644 28432
rect 17500 28008 17552 28014
rect 17500 27950 17552 27956
rect 17604 27946 17632 28426
rect 17696 28218 17724 30280
rect 17880 29481 17908 30534
rect 18064 30054 18092 31726
rect 18512 31680 18564 31686
rect 18234 31648 18290 31657
rect 18512 31622 18564 31628
rect 18234 31583 18290 31592
rect 18144 31408 18196 31414
rect 18144 31350 18196 31356
rect 18156 30705 18184 31350
rect 18248 30818 18276 31583
rect 18524 31278 18552 31622
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18315 31036 18623 31045
rect 18315 31034 18321 31036
rect 18377 31034 18401 31036
rect 18457 31034 18481 31036
rect 18537 31034 18561 31036
rect 18617 31034 18623 31036
rect 18377 30982 18379 31034
rect 18559 30982 18561 31034
rect 18315 30980 18321 30982
rect 18377 30980 18401 30982
rect 18457 30980 18481 30982
rect 18537 30980 18561 30982
rect 18617 30980 18623 30982
rect 18315 30971 18623 30980
rect 18708 30977 18736 31826
rect 18788 31748 18840 31754
rect 18788 31690 18840 31696
rect 19984 31748 20036 31754
rect 19984 31690 20036 31696
rect 18694 30968 18750 30977
rect 18694 30903 18750 30912
rect 18248 30790 18368 30818
rect 18236 30728 18288 30734
rect 18142 30696 18198 30705
rect 18236 30670 18288 30676
rect 18142 30631 18198 30640
rect 18052 30048 18104 30054
rect 17958 30016 18014 30025
rect 18052 29990 18104 29996
rect 18144 30048 18196 30054
rect 18144 29990 18196 29996
rect 17958 29951 18014 29960
rect 17972 29510 18000 29951
rect 18050 29880 18106 29889
rect 18050 29815 18106 29824
rect 18064 29646 18092 29815
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 18156 29578 18184 29990
rect 18144 29572 18196 29578
rect 18144 29514 18196 29520
rect 17960 29504 18012 29510
rect 17866 29472 17922 29481
rect 17960 29446 18012 29452
rect 17866 29407 17922 29416
rect 17958 29336 18014 29345
rect 17958 29271 18014 29280
rect 17866 29200 17922 29209
rect 17972 29170 18000 29271
rect 17866 29135 17922 29144
rect 17960 29164 18012 29170
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17788 28490 17816 28562
rect 17776 28484 17828 28490
rect 17776 28426 17828 28432
rect 17684 28212 17736 28218
rect 17684 28154 17736 28160
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17592 27940 17644 27946
rect 17592 27882 17644 27888
rect 17498 27704 17554 27713
rect 17696 27690 17724 28018
rect 17788 27713 17816 28018
rect 17498 27639 17554 27648
rect 17604 27662 17724 27690
rect 17774 27704 17830 27713
rect 17512 27470 17540 27639
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17406 27296 17462 27305
rect 17406 27231 17462 27240
rect 17408 26920 17460 26926
rect 17408 26862 17460 26868
rect 17144 25894 17356 25922
rect 17144 25412 17172 25894
rect 17224 25832 17276 25838
rect 17276 25792 17356 25820
rect 17224 25774 17276 25780
rect 17224 25424 17276 25430
rect 17144 25384 17224 25412
rect 17224 25366 17276 25372
rect 17328 25294 17356 25792
rect 17224 25288 17276 25294
rect 17222 25256 17224 25265
rect 17316 25288 17368 25294
rect 17276 25256 17278 25265
rect 17316 25230 17368 25236
rect 17222 25191 17278 25200
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17236 24721 17264 24890
rect 17222 24712 17278 24721
rect 17222 24647 17278 24656
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17132 24404 17184 24410
rect 17132 24346 17184 24352
rect 17144 23798 17172 24346
rect 17236 24342 17264 24550
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17328 24274 17356 25230
rect 17316 24268 17368 24274
rect 17316 24210 17368 24216
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17132 23792 17184 23798
rect 17038 23760 17094 23769
rect 16948 23724 17000 23730
rect 17132 23734 17184 23740
rect 17038 23695 17094 23704
rect 16948 23666 17000 23672
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 17236 22778 17264 24142
rect 17328 23866 17356 24210
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17316 22976 17368 22982
rect 17314 22944 17316 22953
rect 17368 22944 17370 22953
rect 17314 22879 17370 22888
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 17420 21962 17448 26862
rect 17512 26450 17540 27406
rect 17500 26444 17552 26450
rect 17500 26386 17552 26392
rect 17512 26353 17540 26386
rect 17498 26344 17554 26353
rect 17498 26279 17554 26288
rect 17498 26208 17554 26217
rect 17498 26143 17554 26152
rect 17512 25906 17540 26143
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17512 25702 17540 25842
rect 17604 25770 17632 27662
rect 17774 27639 17830 27648
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 17696 27305 17724 27542
rect 17682 27296 17738 27305
rect 17682 27231 17738 27240
rect 17880 27130 17908 29135
rect 17960 29106 18012 29112
rect 17972 28937 18000 29106
rect 18052 29096 18104 29102
rect 18052 29038 18104 29044
rect 17958 28928 18014 28937
rect 17958 28863 18014 28872
rect 17958 28792 18014 28801
rect 17958 28727 18014 28736
rect 17972 28393 18000 28727
rect 17958 28384 18014 28393
rect 17958 28319 18014 28328
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17868 27124 17920 27130
rect 17868 27066 17920 27072
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17696 26024 17724 26930
rect 17774 26752 17830 26761
rect 17774 26687 17830 26696
rect 17788 26314 17816 26687
rect 17866 26616 17922 26625
rect 17866 26551 17922 26560
rect 17880 26353 17908 26551
rect 17866 26344 17922 26353
rect 17776 26308 17828 26314
rect 17866 26279 17922 26288
rect 17776 26250 17828 26256
rect 17776 26036 17828 26042
rect 17696 25996 17776 26024
rect 17592 25764 17644 25770
rect 17592 25706 17644 25712
rect 17500 25696 17552 25702
rect 17696 25673 17724 25996
rect 17776 25978 17828 25984
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17500 25638 17552 25644
rect 17682 25664 17738 25673
rect 17682 25599 17738 25608
rect 17788 25537 17816 25842
rect 17498 25528 17554 25537
rect 17498 25463 17554 25472
rect 17774 25528 17830 25537
rect 17774 25463 17830 25472
rect 17512 22574 17540 25463
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 17696 24857 17724 25162
rect 17682 24848 17738 24857
rect 17682 24783 17738 24792
rect 17590 24576 17646 24585
rect 17590 24511 17646 24520
rect 17604 23186 17632 24511
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 17696 22953 17724 24783
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 23526 17816 24550
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17682 22944 17738 22953
rect 17682 22879 17738 22888
rect 17500 22568 17552 22574
rect 17880 22545 17908 25230
rect 17972 23798 18000 27950
rect 18064 24886 18092 29038
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 18050 24712 18106 24721
rect 18050 24647 18106 24656
rect 18064 24138 18092 24647
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 17960 23520 18012 23526
rect 17960 23462 18012 23468
rect 18050 23488 18106 23497
rect 17972 23322 18000 23462
rect 18050 23423 18106 23432
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 18064 23118 18092 23423
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18156 23050 18184 29514
rect 18248 28218 18276 30670
rect 18340 30054 18368 30790
rect 18800 30580 18828 31690
rect 19156 31476 19208 31482
rect 19156 31418 19208 31424
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18892 30802 18920 31282
rect 18972 30932 19024 30938
rect 18972 30874 19024 30880
rect 18880 30796 18932 30802
rect 18880 30738 18932 30744
rect 18800 30552 18920 30580
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18328 30048 18380 30054
rect 18616 30036 18644 30126
rect 18616 30008 18736 30036
rect 18328 29990 18380 29996
rect 18315 29948 18623 29957
rect 18315 29946 18321 29948
rect 18377 29946 18401 29948
rect 18457 29946 18481 29948
rect 18537 29946 18561 29948
rect 18617 29946 18623 29948
rect 18377 29894 18379 29946
rect 18559 29894 18561 29946
rect 18315 29892 18321 29894
rect 18377 29892 18401 29894
rect 18457 29892 18481 29894
rect 18537 29892 18561 29894
rect 18617 29892 18623 29894
rect 18315 29883 18623 29892
rect 18708 29714 18736 30008
rect 18788 29776 18840 29782
rect 18788 29718 18840 29724
rect 18696 29708 18748 29714
rect 18696 29650 18748 29656
rect 18328 29572 18380 29578
rect 18328 29514 18380 29520
rect 18340 29345 18368 29514
rect 18512 29504 18564 29510
rect 18696 29504 18748 29510
rect 18512 29446 18564 29452
rect 18694 29472 18696 29481
rect 18748 29472 18750 29481
rect 18524 29345 18552 29446
rect 18694 29407 18750 29416
rect 18326 29336 18382 29345
rect 18326 29271 18382 29280
rect 18510 29336 18566 29345
rect 18510 29271 18566 29280
rect 18800 29170 18828 29718
rect 18892 29306 18920 30552
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18984 29220 19012 30874
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 19076 30433 19104 30670
rect 19062 30424 19118 30433
rect 19062 30359 19118 30368
rect 19168 30161 19196 31418
rect 19524 31340 19576 31346
rect 19524 31282 19576 31288
rect 19248 31136 19300 31142
rect 19248 31078 19300 31084
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19154 30152 19210 30161
rect 19154 30087 19210 30096
rect 18984 29192 19104 29220
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 18880 29164 18932 29170
rect 18880 29106 18932 29112
rect 18786 28928 18842 28937
rect 18315 28860 18623 28869
rect 18786 28863 18842 28872
rect 18315 28858 18321 28860
rect 18377 28858 18401 28860
rect 18457 28858 18481 28860
rect 18537 28858 18561 28860
rect 18617 28858 18623 28860
rect 18377 28806 18379 28858
rect 18559 28806 18561 28858
rect 18315 28804 18321 28806
rect 18377 28804 18401 28806
rect 18457 28804 18481 28806
rect 18537 28804 18561 28806
rect 18617 28804 18623 28806
rect 18315 28795 18623 28804
rect 18800 28744 18828 28863
rect 18524 28716 18828 28744
rect 18524 28490 18552 28716
rect 18512 28484 18564 28490
rect 18512 28426 18564 28432
rect 18788 28416 18840 28422
rect 18788 28358 18840 28364
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 18604 27872 18656 27878
rect 18656 27849 18736 27860
rect 18656 27840 18750 27849
rect 18656 27832 18694 27840
rect 18604 27814 18656 27820
rect 18315 27772 18623 27781
rect 18694 27775 18750 27784
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 18328 27056 18380 27062
rect 18696 27056 18748 27062
rect 18380 27016 18696 27044
rect 18328 26998 18380 27004
rect 18696 26998 18748 27004
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 18696 26512 18748 26518
rect 18696 26454 18748 26460
rect 18512 26444 18564 26450
rect 18512 26386 18564 26392
rect 18524 25922 18552 26386
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18340 25906 18552 25922
rect 18328 25900 18552 25906
rect 18380 25894 18552 25900
rect 18328 25842 18380 25848
rect 18616 25684 18644 26182
rect 18708 26081 18736 26454
rect 18694 26072 18750 26081
rect 18694 26007 18750 26016
rect 18248 25656 18644 25684
rect 18248 25480 18276 25656
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18708 25537 18736 26007
rect 18694 25528 18750 25537
rect 18328 25492 18380 25498
rect 18248 25452 18328 25480
rect 18694 25463 18750 25472
rect 18328 25434 18380 25440
rect 18696 25424 18748 25430
rect 18696 25366 18748 25372
rect 18708 25294 18736 25366
rect 18236 25288 18288 25294
rect 18696 25288 18748 25294
rect 18236 25230 18288 25236
rect 18604 25266 18656 25272
rect 18248 24818 18276 25230
rect 18696 25230 18748 25236
rect 18604 25208 18656 25214
rect 18328 24948 18380 24954
rect 18616 24936 18644 25208
rect 18616 24908 18736 24936
rect 18328 24890 18380 24896
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18236 24676 18288 24682
rect 18236 24618 18288 24624
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 18248 22817 18276 24618
rect 18340 24614 18368 24890
rect 18708 24857 18736 24908
rect 18694 24848 18750 24857
rect 18694 24783 18750 24792
rect 18512 24744 18564 24750
rect 18510 24712 18512 24721
rect 18564 24712 18566 24721
rect 18510 24647 18566 24656
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18616 23526 18644 24346
rect 18708 23866 18736 24618
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18800 23798 18828 28358
rect 18892 24818 18920 29106
rect 19076 28994 19104 29192
rect 18984 28966 19104 28994
rect 18984 26246 19012 28966
rect 19062 28792 19118 28801
rect 19062 28727 19118 28736
rect 19076 28218 19104 28727
rect 19260 28490 19288 31078
rect 19444 30569 19472 31078
rect 19430 30560 19486 30569
rect 19430 30495 19486 30504
rect 19536 30433 19564 31282
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 19904 30802 19932 31078
rect 19892 30796 19944 30802
rect 19892 30738 19944 30744
rect 19616 30660 19668 30666
rect 19616 30602 19668 30608
rect 19628 30569 19656 30602
rect 19614 30560 19670 30569
rect 19614 30495 19670 30504
rect 19522 30424 19578 30433
rect 19522 30359 19578 30368
rect 19708 30252 19760 30258
rect 19536 30212 19708 30240
rect 19430 30152 19486 30161
rect 19430 30087 19486 30096
rect 19338 29880 19394 29889
rect 19338 29815 19394 29824
rect 19352 28626 19380 29815
rect 19444 29714 19472 30087
rect 19432 29708 19484 29714
rect 19432 29650 19484 29656
rect 19432 28960 19484 28966
rect 19430 28928 19432 28937
rect 19484 28928 19486 28937
rect 19430 28863 19486 28872
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 19248 28144 19300 28150
rect 19246 28112 19248 28121
rect 19300 28112 19302 28121
rect 19064 28076 19116 28082
rect 19246 28047 19302 28056
rect 19064 28018 19116 28024
rect 19076 27606 19104 28018
rect 19352 27962 19380 28562
rect 19260 27934 19380 27962
rect 19064 27600 19116 27606
rect 19064 27542 19116 27548
rect 19064 27396 19116 27402
rect 19116 27356 19196 27384
rect 19064 27338 19116 27344
rect 19062 26344 19118 26353
rect 19062 26279 19118 26288
rect 18972 26240 19024 26246
rect 18972 26182 19024 26188
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18984 25430 19012 25842
rect 19076 25809 19104 26279
rect 19168 26058 19196 27356
rect 19260 27062 19288 27934
rect 19338 27840 19394 27849
rect 19338 27775 19394 27784
rect 19352 27538 19380 27775
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19248 27056 19300 27062
rect 19248 26998 19300 27004
rect 19248 26920 19300 26926
rect 19248 26862 19300 26868
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19260 26761 19288 26862
rect 19246 26752 19302 26761
rect 19246 26687 19302 26696
rect 19352 26314 19380 26862
rect 19340 26308 19392 26314
rect 19340 26250 19392 26256
rect 19168 26030 19288 26058
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 19062 25800 19118 25809
rect 19062 25735 19118 25744
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 19064 25424 19116 25430
rect 19064 25366 19116 25372
rect 18972 25288 19024 25294
rect 18972 25230 19024 25236
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18788 23792 18840 23798
rect 18984 23746 19012 25230
rect 19076 25158 19104 25366
rect 19064 25152 19116 25158
rect 19064 25094 19116 25100
rect 19062 24848 19118 24857
rect 19062 24783 19064 24792
rect 19116 24783 19118 24792
rect 19064 24754 19116 24760
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 19076 24070 19104 24278
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 19076 23798 19104 24006
rect 19168 23866 19196 25910
rect 19260 25498 19288 26030
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19352 25809 19380 25910
rect 19338 25800 19394 25809
rect 19338 25735 19394 25744
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19260 24800 19288 25434
rect 19444 25158 19472 28630
rect 19536 28150 19564 30212
rect 19708 30194 19760 30200
rect 19800 30184 19852 30190
rect 19800 30126 19852 30132
rect 19812 29889 19840 30126
rect 19798 29880 19854 29889
rect 19798 29815 19854 29824
rect 19616 29708 19668 29714
rect 19616 29650 19668 29656
rect 19628 28966 19656 29650
rect 19708 29640 19760 29646
rect 19708 29582 19760 29588
rect 19892 29640 19944 29646
rect 19892 29582 19944 29588
rect 19616 28960 19668 28966
rect 19720 28937 19748 29582
rect 19904 29050 19932 29582
rect 19812 29022 19932 29050
rect 19616 28902 19668 28908
rect 19706 28928 19762 28937
rect 19706 28863 19762 28872
rect 19524 28144 19576 28150
rect 19524 28086 19576 28092
rect 19720 28014 19748 28863
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 19614 27704 19670 27713
rect 19614 27639 19670 27648
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19536 26450 19564 27406
rect 19628 27062 19656 27639
rect 19720 27470 19748 27950
rect 19708 27464 19760 27470
rect 19708 27406 19760 27412
rect 19708 27328 19760 27334
rect 19708 27270 19760 27276
rect 19616 27056 19668 27062
rect 19616 26998 19668 27004
rect 19720 26625 19748 27270
rect 19812 26874 19840 29022
rect 19892 28960 19944 28966
rect 19892 28902 19944 28908
rect 19904 27606 19932 28902
rect 19996 28370 20024 31690
rect 20272 30870 20300 32030
rect 20352 30932 20404 30938
rect 20352 30874 20404 30880
rect 20260 30864 20312 30870
rect 20260 30806 20312 30812
rect 20168 30796 20220 30802
rect 20168 30738 20220 30744
rect 20076 30660 20128 30666
rect 20076 30602 20128 30608
rect 20088 28762 20116 30602
rect 20180 29578 20208 30738
rect 20364 30734 20392 30874
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20260 30660 20312 30666
rect 20260 30602 20312 30608
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 20180 28506 20208 29514
rect 20272 28966 20300 30602
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20364 29034 20392 30194
rect 20456 29850 20484 33200
rect 21560 32094 21588 33200
rect 23768 33130 23796 33200
rect 23860 33130 23888 33238
rect 23768 33102 23888 33130
rect 21548 32088 21600 32094
rect 21548 32030 21600 32036
rect 21640 31748 21692 31754
rect 21640 31690 21692 31696
rect 21100 31470 21404 31498
rect 21100 31414 21128 31470
rect 21376 31414 21404 31470
rect 20628 31408 20680 31414
rect 20628 31350 20680 31356
rect 21088 31408 21140 31414
rect 21088 31350 21140 31356
rect 21180 31408 21232 31414
rect 21364 31408 21416 31414
rect 21232 31368 21312 31396
rect 21180 31350 21232 31356
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20548 30802 20576 31078
rect 20640 30938 20668 31350
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20904 31340 20956 31346
rect 20956 31300 21036 31328
rect 20904 31282 20956 31288
rect 20720 31136 20772 31142
rect 20720 31078 20772 31084
rect 20628 30932 20680 30938
rect 20628 30874 20680 30880
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 20444 29844 20496 29850
rect 20444 29786 20496 29792
rect 20444 29572 20496 29578
rect 20444 29514 20496 29520
rect 20456 29306 20484 29514
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20352 29028 20404 29034
rect 20352 28970 20404 28976
rect 20260 28960 20312 28966
rect 20260 28902 20312 28908
rect 20444 28960 20496 28966
rect 20444 28902 20496 28908
rect 20272 28762 20300 28902
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20456 28626 20484 28902
rect 20444 28620 20496 28626
rect 20444 28562 20496 28568
rect 20180 28478 20300 28506
rect 20168 28416 20220 28422
rect 20074 28384 20130 28393
rect 19996 28342 20074 28370
rect 20168 28358 20220 28364
rect 20074 28319 20130 28328
rect 19984 28144 20036 28150
rect 19984 28086 20036 28092
rect 19996 28014 20024 28086
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19892 27600 19944 27606
rect 19892 27542 19944 27548
rect 19996 26926 20024 27950
rect 20088 27878 20116 28319
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 20180 27713 20208 28358
rect 20272 28257 20300 28478
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 20258 28248 20314 28257
rect 20258 28183 20314 28192
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20166 27704 20222 27713
rect 20166 27639 20222 27648
rect 20166 27568 20222 27577
rect 20166 27503 20222 27512
rect 20180 27470 20208 27503
rect 20168 27464 20220 27470
rect 20168 27406 20220 27412
rect 20166 27296 20222 27305
rect 20166 27231 20222 27240
rect 19984 26920 20036 26926
rect 19812 26846 19932 26874
rect 19984 26862 20036 26868
rect 19800 26784 19852 26790
rect 19800 26726 19852 26732
rect 19706 26616 19762 26625
rect 19706 26551 19762 26560
rect 19524 26444 19576 26450
rect 19524 26386 19576 26392
rect 19720 26234 19748 26551
rect 19812 26382 19840 26726
rect 19800 26376 19852 26382
rect 19798 26344 19800 26353
rect 19852 26344 19854 26353
rect 19798 26279 19854 26288
rect 19720 26206 19840 26234
rect 19522 26072 19578 26081
rect 19522 26007 19578 26016
rect 19616 26036 19668 26042
rect 19536 25294 19564 26007
rect 19616 25978 19668 25984
rect 19708 26036 19760 26042
rect 19708 25978 19760 25984
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19340 24812 19392 24818
rect 19260 24772 19340 24800
rect 19340 24754 19392 24760
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 18788 23734 18840 23740
rect 18892 23718 19012 23746
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18234 22808 18290 22817
rect 18234 22743 18290 22752
rect 17500 22510 17552 22516
rect 17866 22536 17922 22545
rect 17866 22471 17922 22480
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18892 22094 18920 23718
rect 18972 22772 19024 22778
rect 19076 22760 19104 23734
rect 19352 23322 19380 24550
rect 19430 24440 19486 24449
rect 19430 24375 19486 24384
rect 19444 23798 19472 24375
rect 19536 24070 19564 24890
rect 19628 24868 19656 25978
rect 19720 25129 19748 25978
rect 19812 25362 19840 26206
rect 19800 25356 19852 25362
rect 19800 25298 19852 25304
rect 19800 25220 19852 25226
rect 19800 25162 19852 25168
rect 19706 25120 19762 25129
rect 19706 25055 19762 25064
rect 19708 24880 19760 24886
rect 19628 24840 19708 24868
rect 19708 24822 19760 24828
rect 19812 24449 19840 25162
rect 19798 24440 19854 24449
rect 19708 24404 19760 24410
rect 19798 24375 19854 24384
rect 19708 24346 19760 24352
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19614 23624 19670 23633
rect 19536 23497 19564 23598
rect 19614 23559 19670 23568
rect 19522 23488 19578 23497
rect 19522 23423 19578 23432
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19522 23080 19578 23089
rect 19522 23015 19578 23024
rect 19536 22982 19564 23015
rect 19524 22976 19576 22982
rect 19524 22918 19576 22924
rect 19024 22732 19104 22760
rect 18972 22714 19024 22720
rect 18708 22066 18920 22094
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 18708 21622 18736 22066
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 1584 21480 1636 21486
rect 1582 21448 1584 21457
rect 12348 21480 12400 21486
rect 1636 21448 1638 21457
rect 12348 21422 12400 21428
rect 19076 21418 19104 22732
rect 19628 21978 19656 23559
rect 19720 23361 19748 24346
rect 19904 24342 19932 26846
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 19996 25838 20024 26726
rect 20180 26246 20208 27231
rect 20168 26240 20220 26246
rect 20168 26182 20220 26188
rect 20074 25936 20130 25945
rect 20074 25871 20130 25880
rect 20168 25900 20220 25906
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 20088 25702 20116 25871
rect 20168 25842 20220 25848
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 20180 25498 20208 25842
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 19984 25220 20036 25226
rect 19984 25162 20036 25168
rect 19996 25129 20024 25162
rect 19982 25120 20038 25129
rect 19982 25055 20038 25064
rect 20166 25120 20222 25129
rect 20166 25055 20222 25064
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19984 24676 20036 24682
rect 19984 24618 20036 24624
rect 19892 24336 19944 24342
rect 19892 24278 19944 24284
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19904 24070 19932 24142
rect 19800 24064 19852 24070
rect 19800 24006 19852 24012
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19706 23352 19762 23361
rect 19706 23287 19762 23296
rect 19812 23254 19840 24006
rect 19996 23848 20024 24618
rect 20088 24585 20116 24754
rect 20074 24576 20130 24585
rect 20074 24511 20130 24520
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19904 23820 20024 23848
rect 19904 23662 19932 23820
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19892 23656 19944 23662
rect 19892 23598 19944 23604
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19800 23248 19852 23254
rect 19800 23190 19852 23196
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19812 22098 19840 22714
rect 19904 22710 19932 23462
rect 19996 22982 20024 23666
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19996 22817 20024 22918
rect 19982 22808 20038 22817
rect 19982 22743 20038 22752
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19904 22166 19932 22646
rect 19996 22166 20024 22743
rect 20088 22438 20116 24142
rect 20180 24138 20208 25055
rect 20272 24342 20300 28018
rect 20350 27568 20406 27577
rect 20350 27503 20406 27512
rect 20364 26994 20392 27503
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 20364 25906 20392 26930
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 20364 24342 20392 25706
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20352 24336 20404 24342
rect 20352 24278 20404 24284
rect 20258 24168 20314 24177
rect 20168 24132 20220 24138
rect 20258 24103 20314 24112
rect 20168 24074 20220 24080
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20180 23610 20208 23734
rect 20272 23730 20300 24103
rect 20350 24032 20406 24041
rect 20350 23967 20406 23976
rect 20364 23798 20392 23967
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20180 23582 20300 23610
rect 20272 23322 20300 23582
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20168 23248 20220 23254
rect 20168 23190 20220 23196
rect 20180 22982 20208 23190
rect 20168 22976 20220 22982
rect 20168 22918 20220 22924
rect 20272 22778 20300 23258
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19892 22160 19944 22166
rect 19892 22102 19944 22108
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19800 22092 19852 22098
rect 19800 22034 19852 22040
rect 19536 21950 19656 21978
rect 19430 21856 19486 21865
rect 19430 21791 19486 21800
rect 19444 21690 19472 21791
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 1582 21383 1638 21392
rect 19064 21412 19116 21418
rect 19064 21354 19116 21360
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18800 21078 18828 21286
rect 19536 21078 19564 21950
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 19982 20632 20038 20641
rect 19982 20567 19984 20576
rect 20036 20567 20038 20576
rect 19984 20538 20036 20544
rect 20088 20466 20116 22374
rect 20166 22264 20222 22273
rect 20166 22199 20222 22208
rect 20180 22166 20208 22199
rect 20272 22166 20300 22714
rect 20168 22160 20220 22166
rect 20168 22102 20220 22108
rect 20260 22160 20312 22166
rect 20260 22102 20312 22108
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20272 20534 20300 21966
rect 20364 21146 20392 23734
rect 20456 23254 20484 28358
rect 20548 27849 20576 30602
rect 20626 30424 20682 30433
rect 20626 30359 20682 30368
rect 20640 30326 20668 30359
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20626 29608 20682 29617
rect 20626 29543 20682 29552
rect 20640 28937 20668 29543
rect 20732 29238 20760 31078
rect 20824 29714 20852 31282
rect 21008 30297 21036 31300
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 20994 30288 21050 30297
rect 20994 30223 21050 30232
rect 21192 30190 21220 30670
rect 21284 30569 21312 31368
rect 21364 31350 21416 31356
rect 21548 31340 21600 31346
rect 21468 31300 21548 31328
rect 21468 30648 21496 31300
rect 21548 31282 21600 31288
rect 21652 30784 21680 31690
rect 22652 31680 22704 31686
rect 22652 31622 22704 31628
rect 22744 31680 22796 31686
rect 22744 31622 22796 31628
rect 21788 31580 22096 31589
rect 21788 31578 21794 31580
rect 21850 31578 21874 31580
rect 21930 31578 21954 31580
rect 22010 31578 22034 31580
rect 22090 31578 22096 31580
rect 21850 31526 21852 31578
rect 22032 31526 22034 31578
rect 21788 31524 21794 31526
rect 21850 31524 21874 31526
rect 21930 31524 21954 31526
rect 22010 31524 22034 31526
rect 22090 31524 22096 31526
rect 21788 31515 22096 31524
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21916 31204 21968 31210
rect 21916 31146 21968 31152
rect 21730 31104 21786 31113
rect 21730 31039 21786 31048
rect 21744 30938 21772 31039
rect 21732 30932 21784 30938
rect 21732 30874 21784 30880
rect 21652 30756 21772 30784
rect 21744 30666 21772 30756
rect 21928 30734 21956 31146
rect 22112 30802 22140 31214
rect 22100 30796 22152 30802
rect 22100 30738 22152 30744
rect 22664 30734 22692 31622
rect 21916 30728 21968 30734
rect 21916 30670 21968 30676
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 21367 30620 21496 30648
rect 21640 30660 21692 30666
rect 21270 30560 21326 30569
rect 21367 30546 21395 30620
rect 21640 30602 21692 30608
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 21548 30592 21600 30598
rect 21454 30560 21510 30569
rect 21367 30518 21404 30546
rect 21270 30495 21326 30504
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 21272 30116 21324 30122
rect 21272 30058 21324 30064
rect 21180 30048 21232 30054
rect 21180 29990 21232 29996
rect 21086 29744 21142 29753
rect 20812 29708 20864 29714
rect 21086 29679 21142 29688
rect 20812 29650 20864 29656
rect 20720 29232 20772 29238
rect 20720 29174 20772 29180
rect 20626 28928 20682 28937
rect 20626 28863 20682 28872
rect 20824 28694 20852 29650
rect 21100 29646 21128 29679
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 21088 29504 21140 29510
rect 20994 29472 21050 29481
rect 21088 29446 21140 29452
rect 20994 29407 21050 29416
rect 21008 29238 21036 29407
rect 21100 29306 21128 29446
rect 21088 29300 21140 29306
rect 21088 29242 21140 29248
rect 20996 29232 21048 29238
rect 20996 29174 21048 29180
rect 20994 29064 21050 29073
rect 20994 28999 21050 29008
rect 20812 28688 20864 28694
rect 20812 28630 20864 28636
rect 20718 28248 20774 28257
rect 20718 28183 20774 28192
rect 20534 27840 20590 27849
rect 20534 27775 20590 27784
rect 20732 27470 20760 28183
rect 20812 28144 20864 28150
rect 20812 28086 20864 28092
rect 20824 27996 20852 28086
rect 20824 27968 20944 27996
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 20536 27056 20588 27062
rect 20536 26998 20588 27004
rect 20548 25140 20576 26998
rect 20640 25242 20668 27406
rect 20718 27160 20774 27169
rect 20718 27095 20774 27104
rect 20732 26761 20760 27095
rect 20718 26752 20774 26761
rect 20718 26687 20774 26696
rect 20824 26518 20852 27814
rect 20812 26512 20864 26518
rect 20718 26480 20774 26489
rect 20812 26454 20864 26460
rect 20718 26415 20774 26424
rect 20732 26314 20760 26415
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20810 25936 20866 25945
rect 20810 25871 20812 25880
rect 20864 25871 20866 25880
rect 20812 25842 20864 25848
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20640 25226 20760 25242
rect 20640 25220 20772 25226
rect 20640 25214 20720 25220
rect 20720 25162 20772 25168
rect 20548 25112 20668 25140
rect 20640 24138 20668 25112
rect 20824 24993 20852 25638
rect 20810 24984 20866 24993
rect 20810 24919 20866 24928
rect 20718 24440 20774 24449
rect 20718 24375 20774 24384
rect 20732 24206 20760 24375
rect 20810 24304 20866 24313
rect 20810 24239 20866 24248
rect 20824 24206 20852 24239
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20626 23896 20682 23905
rect 20626 23831 20682 23840
rect 20640 23730 20668 23831
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20626 23488 20682 23497
rect 20626 23423 20682 23432
rect 20534 23352 20590 23361
rect 20534 23287 20536 23296
rect 20588 23287 20590 23296
rect 20536 23258 20588 23264
rect 20444 23248 20496 23254
rect 20444 23190 20496 23196
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20456 22710 20484 22918
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20444 22432 20496 22438
rect 20548 22420 20576 23258
rect 20496 22392 20576 22420
rect 20444 22374 20496 22380
rect 20456 22234 20484 22374
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20456 21418 20484 22170
rect 20534 21584 20590 21593
rect 20534 21519 20590 21528
rect 20444 21412 20496 21418
rect 20444 21354 20496 21360
rect 20456 21146 20484 21354
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20548 20942 20576 21519
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20097 1624 20198
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 1582 20088 1638 20097
rect 4423 20091 4731 20100
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 20640 20058 20668 23423
rect 20732 23050 20760 24142
rect 20916 23905 20944 27968
rect 21008 27606 21036 28999
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 20996 27600 21048 27606
rect 20996 27542 21048 27548
rect 20996 26512 21048 26518
rect 20996 26454 21048 26460
rect 20902 23896 20958 23905
rect 20812 23860 20864 23866
rect 20902 23831 20958 23840
rect 20812 23802 20864 23808
rect 20824 23361 20852 23802
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 20810 23352 20866 23361
rect 20810 23287 20866 23296
rect 20916 23118 20944 23666
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 20718 22808 20774 22817
rect 20718 22743 20774 22752
rect 20732 22710 20760 22743
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20824 21962 20852 22918
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20812 21956 20864 21962
rect 20812 21898 20864 21904
rect 20824 21865 20852 21898
rect 20810 21856 20866 21865
rect 20810 21791 20866 21800
rect 20824 21146 20852 21791
rect 20916 21350 20944 22714
rect 21008 22001 21036 26454
rect 21100 26382 21128 28358
rect 21192 28150 21220 29990
rect 21284 29782 21312 30058
rect 21272 29776 21324 29782
rect 21272 29718 21324 29724
rect 21272 29300 21324 29306
rect 21272 29242 21324 29248
rect 21180 28144 21232 28150
rect 21180 28086 21232 28092
rect 21284 26790 21312 29242
rect 21376 27305 21404 30518
rect 21548 30534 21600 30540
rect 21454 30495 21510 30504
rect 21468 27860 21496 30495
rect 21560 28082 21588 30534
rect 21652 29034 21680 30602
rect 22652 30592 22704 30598
rect 22652 30534 22704 30540
rect 21788 30492 22096 30501
rect 21788 30490 21794 30492
rect 21850 30490 21874 30492
rect 21930 30490 21954 30492
rect 22010 30490 22034 30492
rect 22090 30490 22096 30492
rect 21850 30438 21852 30490
rect 22032 30438 22034 30490
rect 21788 30436 21794 30438
rect 21850 30436 21874 30438
rect 21930 30436 21954 30438
rect 22010 30436 22034 30438
rect 22090 30436 22096 30438
rect 21788 30427 22096 30436
rect 22558 30424 22614 30433
rect 22558 30359 22614 30368
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 21788 29404 22096 29413
rect 21788 29402 21794 29404
rect 21850 29402 21874 29404
rect 21930 29402 21954 29404
rect 22010 29402 22034 29404
rect 22090 29402 22096 29404
rect 21850 29350 21852 29402
rect 22032 29350 22034 29402
rect 21788 29348 21794 29350
rect 21850 29348 21874 29350
rect 21930 29348 21954 29350
rect 22010 29348 22034 29350
rect 22090 29348 22096 29350
rect 21788 29339 22096 29348
rect 22296 29073 22324 30194
rect 22376 29640 22428 29646
rect 22376 29582 22428 29588
rect 22388 29102 22416 29582
rect 22376 29096 22428 29102
rect 22282 29064 22338 29073
rect 21640 29028 21692 29034
rect 22376 29038 22428 29044
rect 22282 28999 22338 29008
rect 21640 28970 21692 28976
rect 21548 28076 21600 28082
rect 21548 28018 21600 28024
rect 21548 27872 21600 27878
rect 21468 27832 21548 27860
rect 21548 27814 21600 27820
rect 21362 27296 21418 27305
rect 21362 27231 21418 27240
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21178 26616 21234 26625
rect 21178 26551 21234 26560
rect 21192 26382 21220 26551
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21178 26208 21234 26217
rect 21178 26143 21234 26152
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 21100 22710 21128 25434
rect 21192 24596 21220 26143
rect 21284 24954 21312 26726
rect 21376 26042 21404 27066
rect 21454 26888 21510 26897
rect 21454 26823 21510 26832
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 21468 25945 21496 26823
rect 21560 26081 21588 27814
rect 21546 26072 21602 26081
rect 21546 26007 21602 26016
rect 21454 25936 21510 25945
rect 21454 25871 21510 25880
rect 21362 25528 21418 25537
rect 21362 25463 21418 25472
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 21376 24886 21404 25463
rect 21364 24880 21416 24886
rect 21364 24822 21416 24828
rect 21468 24614 21496 25871
rect 21652 25129 21680 28970
rect 22388 28694 22416 29038
rect 22376 28688 22428 28694
rect 22376 28630 22428 28636
rect 22388 28558 22416 28630
rect 22376 28552 22428 28558
rect 22020 28490 22232 28506
rect 22376 28494 22428 28500
rect 22008 28484 22232 28490
rect 22060 28478 22232 28484
rect 22008 28426 22060 28432
rect 21788 28316 22096 28325
rect 21788 28314 21794 28316
rect 21850 28314 21874 28316
rect 21930 28314 21954 28316
rect 22010 28314 22034 28316
rect 22090 28314 22096 28316
rect 21850 28262 21852 28314
rect 22032 28262 22034 28314
rect 21788 28260 21794 28262
rect 21850 28260 21874 28262
rect 21930 28260 21954 28262
rect 22010 28260 22034 28262
rect 22090 28260 22096 28262
rect 21788 28251 22096 28260
rect 21732 28144 21784 28150
rect 21732 28086 21784 28092
rect 21744 27334 21772 28086
rect 21732 27328 21784 27334
rect 21732 27270 21784 27276
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 22006 27024 22062 27033
rect 22006 26959 22062 26968
rect 22020 26926 22048 26959
rect 22008 26920 22060 26926
rect 21730 26888 21786 26897
rect 22008 26862 22060 26868
rect 22204 26874 22232 28478
rect 22284 28484 22336 28490
rect 22284 28426 22336 28432
rect 22296 27849 22324 28426
rect 22388 28014 22416 28494
rect 22376 28008 22428 28014
rect 22428 27968 22508 27996
rect 22376 27950 22428 27956
rect 22376 27872 22428 27878
rect 22282 27840 22338 27849
rect 22376 27814 22428 27820
rect 22282 27775 22338 27784
rect 22388 27470 22416 27814
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 22296 26994 22324 27066
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 22204 26846 22416 26874
rect 21730 26823 21732 26832
rect 21784 26823 21786 26832
rect 21732 26794 21784 26800
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 22098 26616 22154 26625
rect 22098 26551 22154 26560
rect 22112 26314 22140 26551
rect 22100 26308 22152 26314
rect 22100 26250 22152 26256
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 21732 25900 21784 25906
rect 21732 25842 21784 25848
rect 21744 25702 21772 25842
rect 22008 25832 22060 25838
rect 22204 25820 22232 26182
rect 22060 25792 22232 25820
rect 22008 25774 22060 25780
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 21824 25696 21876 25702
rect 21824 25638 21876 25644
rect 21836 25294 21864 25638
rect 22098 25528 22154 25537
rect 22098 25463 22154 25472
rect 22112 25294 22140 25463
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 22100 25288 22152 25294
rect 22152 25248 22232 25276
rect 22100 25230 22152 25236
rect 21638 25120 21694 25129
rect 21638 25055 21694 25064
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 22204 24614 22232 25248
rect 21456 24608 21508 24614
rect 21192 24568 21312 24596
rect 21178 24440 21234 24449
rect 21178 24375 21234 24384
rect 21192 24342 21220 24375
rect 21180 24336 21232 24342
rect 21180 24278 21232 24284
rect 21284 24206 21312 24568
rect 21456 24550 21508 24556
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 21192 23730 21220 24074
rect 21284 24041 21312 24142
rect 21640 24132 21692 24138
rect 21376 24092 21640 24120
rect 21270 24032 21326 24041
rect 21270 23967 21326 23976
rect 21270 23760 21326 23769
rect 21180 23724 21232 23730
rect 21376 23730 21404 24092
rect 21640 24074 21692 24080
rect 21638 24032 21694 24041
rect 21638 23967 21694 23976
rect 21546 23760 21602 23769
rect 21270 23695 21326 23704
rect 21364 23724 21416 23730
rect 21180 23666 21232 23672
rect 21192 23633 21220 23666
rect 21178 23624 21234 23633
rect 21178 23559 21234 23568
rect 21284 23186 21312 23695
rect 21364 23666 21416 23672
rect 21456 23724 21508 23730
rect 21546 23695 21602 23704
rect 21456 23666 21508 23672
rect 21376 23497 21404 23666
rect 21362 23488 21418 23497
rect 21362 23423 21418 23432
rect 21272 23180 21324 23186
rect 21272 23122 21324 23128
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 21192 22012 21220 22986
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21270 22128 21326 22137
rect 21376 22098 21404 22374
rect 21270 22063 21326 22072
rect 21364 22092 21416 22098
rect 21284 22030 21312 22063
rect 21364 22034 21416 22040
rect 20994 21992 21050 22001
rect 20994 21927 21050 21936
rect 21100 21984 21220 22012
rect 21272 22024 21324 22030
rect 21100 21400 21128 21984
rect 21272 21966 21324 21972
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 21376 21570 21404 22034
rect 21468 21690 21496 23666
rect 21560 23662 21588 23695
rect 21548 23656 21600 23662
rect 21548 23598 21600 23604
rect 21652 23644 21680 23967
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 22190 23896 22246 23905
rect 21836 23840 22190 23848
rect 21836 23831 22246 23840
rect 21836 23820 22232 23831
rect 21732 23656 21784 23662
rect 21652 23616 21732 23644
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21008 21372 21128 21400
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 21008 20602 21036 21372
rect 21192 21321 21220 21558
rect 21284 21332 21312 21558
rect 21376 21542 21496 21570
rect 21468 21350 21496 21542
rect 21364 21344 21416 21350
rect 21178 21312 21234 21321
rect 21284 21304 21364 21332
rect 21364 21286 21416 21292
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21178 21247 21234 21256
rect 21376 21146 21404 21286
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 1582 20023 1638 20032
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19417 1624 19790
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 21100 18358 21128 21014
rect 21652 20058 21680 23616
rect 21732 23598 21784 23604
rect 21836 23322 21864 23820
rect 21916 23724 21968 23730
rect 21916 23666 21968 23672
rect 21824 23316 21876 23322
rect 21824 23258 21876 23264
rect 21928 23186 21956 23666
rect 22008 23656 22060 23662
rect 22006 23624 22008 23633
rect 22060 23624 22062 23633
rect 22006 23559 22062 23568
rect 22098 23488 22154 23497
rect 22098 23423 22154 23432
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 21822 23080 21878 23089
rect 21822 23015 21824 23024
rect 21876 23015 21878 23024
rect 21824 22986 21876 22992
rect 22112 22964 22140 23423
rect 22192 23112 22244 23118
rect 22192 23054 22244 23060
rect 22112 22936 22171 22964
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 22143 22778 22171 22936
rect 22100 22772 22171 22778
rect 22152 22732 22171 22772
rect 22100 22714 22152 22720
rect 22204 22681 22232 23054
rect 21822 22672 21878 22681
rect 21822 22607 21824 22616
rect 21876 22607 21878 22616
rect 22190 22672 22246 22681
rect 22296 22676 22324 26726
rect 22388 24818 22416 26846
rect 22480 25537 22508 27968
rect 22572 27713 22600 30359
rect 22558 27704 22614 27713
rect 22558 27639 22614 27648
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 22572 27169 22600 27542
rect 22664 27402 22692 30534
rect 22756 28150 22784 31622
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 22928 29640 22980 29646
rect 22926 29608 22928 29617
rect 22980 29608 22982 29617
rect 22926 29543 22982 29552
rect 22926 29472 22982 29481
rect 22926 29407 22982 29416
rect 22834 28792 22890 28801
rect 22834 28727 22890 28736
rect 22744 28144 22796 28150
rect 22744 28086 22796 28092
rect 22742 27840 22798 27849
rect 22742 27775 22798 27784
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22558 27160 22614 27169
rect 22558 27095 22614 27104
rect 22558 27024 22614 27033
rect 22558 26959 22614 26968
rect 22466 25528 22522 25537
rect 22466 25463 22522 25472
rect 22468 24880 22520 24886
rect 22468 24822 22520 24828
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22190 22607 22246 22616
rect 22284 22670 22336 22676
rect 22284 22612 22336 22618
rect 21824 22578 21876 22584
rect 22284 22432 22336 22438
rect 22282 22400 22284 22409
rect 22336 22400 22338 22409
rect 22282 22335 22338 22344
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 22296 20058 22324 22170
rect 22388 21894 22416 24550
rect 22480 23032 22508 24822
rect 22572 23730 22600 26959
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22480 23004 22600 23032
rect 22466 22808 22522 22817
rect 22466 22743 22468 22752
rect 22520 22743 22522 22752
rect 22468 22714 22520 22720
rect 22466 22128 22522 22137
rect 22466 22063 22522 22072
rect 22480 21962 22508 22063
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22468 21616 22520 21622
rect 22466 21584 22468 21593
rect 22520 21584 22522 21593
rect 22466 21519 22522 21528
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 21078 22416 21286
rect 22376 21072 22428 21078
rect 22428 21032 22508 21060
rect 22376 21014 22428 21020
rect 22480 20602 22508 21032
rect 22572 20874 22600 23004
rect 22664 21962 22692 27338
rect 22756 25498 22784 27775
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22756 24886 22784 25230
rect 22848 25129 22876 28727
rect 22940 28558 22968 29407
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 23124 28937 23152 29106
rect 23110 28928 23166 28937
rect 23110 28863 23166 28872
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 22928 28552 22980 28558
rect 22980 28500 23060 28506
rect 22928 28494 23060 28500
rect 22940 28478 23060 28494
rect 23032 28393 23060 28478
rect 23018 28384 23074 28393
rect 23018 28319 23074 28328
rect 23124 27713 23152 28562
rect 23110 27704 23166 27713
rect 23110 27639 23166 27648
rect 23110 27568 23166 27577
rect 23110 27503 23166 27512
rect 23020 27464 23072 27470
rect 22940 27424 23020 27452
rect 22834 25120 22890 25129
rect 22834 25055 22890 25064
rect 22744 24880 22796 24886
rect 22744 24822 22796 24828
rect 22834 24440 22890 24449
rect 22834 24375 22890 24384
rect 22848 24342 22876 24375
rect 22940 24342 22968 27424
rect 23020 27406 23072 27412
rect 23124 27169 23152 27503
rect 23110 27160 23166 27169
rect 23110 27095 23166 27104
rect 23020 26852 23072 26858
rect 23020 26794 23072 26800
rect 23032 26382 23060 26794
rect 23216 26518 23244 31418
rect 23940 31272 23992 31278
rect 23940 31214 23992 31220
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 23480 30728 23532 30734
rect 23480 30670 23532 30676
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23492 30598 23520 30670
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23388 30048 23440 30054
rect 23388 29990 23440 29996
rect 23400 29782 23428 29990
rect 23388 29776 23440 29782
rect 23388 29718 23440 29724
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23296 28076 23348 28082
rect 23296 28018 23348 28024
rect 23308 27849 23336 28018
rect 23400 28014 23428 29038
rect 23570 28928 23626 28937
rect 23570 28863 23626 28872
rect 23388 28008 23440 28014
rect 23388 27950 23440 27956
rect 23294 27840 23350 27849
rect 23294 27775 23350 27784
rect 23584 27606 23612 28863
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23676 28665 23704 28698
rect 23662 28656 23718 28665
rect 23662 28591 23718 28600
rect 23768 28393 23796 30670
rect 23860 30326 23888 31078
rect 23952 30734 23980 31214
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23848 30320 23900 30326
rect 23848 30262 23900 30268
rect 23848 30184 23900 30190
rect 23848 30126 23900 30132
rect 23860 29578 23888 30126
rect 23848 29572 23900 29578
rect 23848 29514 23900 29520
rect 23860 29102 23888 29514
rect 23848 29096 23900 29102
rect 23848 29038 23900 29044
rect 23848 28960 23900 28966
rect 23848 28902 23900 28908
rect 23860 28762 23888 28902
rect 23848 28756 23900 28762
rect 23848 28698 23900 28704
rect 23754 28384 23810 28393
rect 23754 28319 23810 28328
rect 23756 28076 23808 28082
rect 23676 28036 23756 28064
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23308 26625 23336 27406
rect 23388 27396 23440 27402
rect 23388 27338 23440 27344
rect 23400 26897 23428 27338
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23386 26888 23442 26897
rect 23386 26823 23442 26832
rect 23294 26616 23350 26625
rect 23294 26551 23350 26560
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23204 26512 23256 26518
rect 23204 26454 23256 26460
rect 23400 26382 23428 26522
rect 23020 26376 23072 26382
rect 23388 26376 23440 26382
rect 23072 26336 23244 26364
rect 23020 26318 23072 26324
rect 23112 26240 23164 26246
rect 23110 26208 23112 26217
rect 23164 26208 23166 26217
rect 23110 26143 23166 26152
rect 23112 25764 23164 25770
rect 23032 25724 23112 25752
rect 23032 25226 23060 25724
rect 23112 25706 23164 25712
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 22836 24336 22888 24342
rect 22836 24278 22888 24284
rect 22928 24336 22980 24342
rect 22928 24278 22980 24284
rect 22848 24177 22876 24278
rect 23032 24274 23060 25162
rect 23124 24410 23152 25434
rect 23216 24886 23244 26336
rect 23388 26318 23440 26324
rect 23296 26240 23348 26246
rect 23296 26182 23348 26188
rect 23308 25294 23336 26182
rect 23386 26072 23442 26081
rect 23386 26007 23442 26016
rect 23400 25702 23428 26007
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 23308 24993 23336 25094
rect 23294 24984 23350 24993
rect 23294 24919 23350 24928
rect 23204 24880 23256 24886
rect 23204 24822 23256 24828
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23020 24268 23072 24274
rect 23020 24210 23072 24216
rect 23216 24177 23244 24550
rect 22834 24168 22890 24177
rect 22834 24103 22890 24112
rect 23202 24168 23258 24177
rect 23202 24103 23258 24112
rect 22834 24032 22890 24041
rect 22834 23967 22890 23976
rect 22848 22642 22876 23967
rect 23112 22976 23164 22982
rect 23018 22944 23074 22953
rect 23112 22918 23164 22924
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 23018 22879 23074 22888
rect 23032 22642 23060 22879
rect 23124 22710 23152 22918
rect 23112 22704 23164 22710
rect 23112 22646 23164 22652
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22652 21344 22704 21350
rect 22650 21312 22652 21321
rect 22704 21312 22706 21321
rect 22650 21247 22706 21256
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 21652 19514 21680 19994
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 22388 18630 22416 20470
rect 22572 19334 22600 20810
rect 22664 20602 22692 20878
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22664 19922 22692 20538
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22664 19514 22692 19858
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22480 19306 22600 19334
rect 22480 18630 22508 19306
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 1584 18080 1636 18086
rect 1582 18048 1584 18057
rect 1636 18048 1638 18057
rect 1582 17983 1638 17992
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 17377 1624 17614
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 1582 17368 1638 17377
rect 7896 17371 8204 17380
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 1582 17303 1638 17312
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 22388 16250 22416 18566
rect 22756 17882 22784 21830
rect 22848 20466 22876 22578
rect 22928 22568 22980 22574
rect 22928 22510 22980 22516
rect 22940 20602 22968 22510
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 23032 22137 23060 22170
rect 23018 22128 23074 22137
rect 23018 22063 23074 22072
rect 23018 21992 23074 22001
rect 23018 21927 23020 21936
rect 23072 21927 23074 21936
rect 23020 21898 23072 21904
rect 23124 21434 23152 22646
rect 23216 22273 23244 22918
rect 23308 22817 23336 24754
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 23361 23428 24550
rect 23492 24070 23520 25094
rect 23584 24410 23612 27270
rect 23676 26790 23704 28036
rect 23756 28018 23808 28024
rect 23848 28008 23900 28014
rect 23900 27968 23980 27996
rect 23848 27950 23900 27956
rect 23848 27872 23900 27878
rect 23846 27840 23848 27849
rect 23900 27840 23902 27849
rect 23846 27775 23902 27784
rect 23848 27668 23900 27674
rect 23848 27610 23900 27616
rect 23754 27568 23810 27577
rect 23754 27503 23810 27512
rect 23664 26784 23716 26790
rect 23664 26726 23716 26732
rect 23768 26518 23796 27503
rect 23860 27130 23888 27610
rect 23952 27470 23980 27968
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23848 27124 23900 27130
rect 23848 27066 23900 27072
rect 23952 26858 23980 27406
rect 23940 26852 23992 26858
rect 23940 26794 23992 26800
rect 23756 26512 23808 26518
rect 23662 26480 23718 26489
rect 23756 26454 23808 26460
rect 23662 26415 23718 26424
rect 23676 26314 23704 26415
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 23664 26308 23716 26314
rect 23664 26250 23716 26256
rect 23860 26042 23888 26318
rect 23940 26240 23992 26246
rect 23940 26182 23992 26188
rect 23664 26036 23716 26042
rect 23664 25978 23716 25984
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23676 25906 23704 25978
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 23676 25294 23704 25842
rect 23952 25786 23980 26182
rect 23860 25758 23980 25786
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23572 24404 23624 24410
rect 23572 24346 23624 24352
rect 23572 24200 23624 24206
rect 23768 24188 23796 25434
rect 23624 24160 23796 24188
rect 23572 24142 23624 24148
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23584 23866 23612 24142
rect 23572 23860 23624 23866
rect 23624 23820 23704 23848
rect 23572 23802 23624 23808
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23386 23352 23442 23361
rect 23386 23287 23442 23296
rect 23294 22808 23350 22817
rect 23294 22743 23350 22752
rect 23386 22536 23442 22545
rect 23492 22522 23520 23598
rect 23570 22672 23626 22681
rect 23570 22607 23572 22616
rect 23624 22607 23626 22616
rect 23572 22578 23624 22584
rect 23492 22494 23612 22522
rect 23386 22471 23442 22480
rect 23202 22264 23258 22273
rect 23202 22199 23258 22208
rect 23400 22166 23428 22471
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 23386 21992 23442 22001
rect 23386 21927 23442 21936
rect 23400 21894 23428 21927
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23294 21720 23350 21729
rect 23294 21655 23350 21664
rect 23308 21622 23336 21655
rect 23296 21616 23348 21622
rect 23296 21558 23348 21564
rect 23032 21406 23152 21434
rect 23032 20942 23060 21406
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23124 20534 23152 21286
rect 23112 20528 23164 20534
rect 23112 20470 23164 20476
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 23584 18970 23612 22494
rect 23676 19514 23704 23820
rect 23860 23798 23888 25758
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23848 23792 23900 23798
rect 23848 23734 23900 23740
rect 23848 23520 23900 23526
rect 23952 23497 23980 25638
rect 23848 23462 23900 23468
rect 23938 23488 23994 23497
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23768 21554 23796 23258
rect 23860 23118 23888 23462
rect 23938 23423 23994 23432
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23860 22574 23888 23054
rect 23938 22808 23994 22817
rect 23938 22743 23994 22752
rect 23952 22642 23980 22743
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 24044 21554 24072 33238
rect 24858 33200 24914 34000
rect 24964 33238 25820 33266
rect 24872 33130 24900 33200
rect 24964 33130 24992 33238
rect 24872 33102 24992 33130
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 24492 31272 24544 31278
rect 24492 31214 24544 31220
rect 24308 30592 24360 30598
rect 24308 30534 24360 30540
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24124 29640 24176 29646
rect 24124 29582 24176 29588
rect 24136 27130 24164 29582
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 24136 25838 24164 27066
rect 24124 25832 24176 25838
rect 24124 25774 24176 25780
rect 24228 24664 24256 30262
rect 24136 24636 24256 24664
rect 24136 24449 24164 24636
rect 24320 24562 24348 30534
rect 24398 29336 24454 29345
rect 24398 29271 24454 29280
rect 24412 28626 24440 29271
rect 24400 28620 24452 28626
rect 24400 28562 24452 28568
rect 24504 28234 24532 31214
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24596 30394 24624 30534
rect 24584 30388 24636 30394
rect 24584 30330 24636 30336
rect 24582 30288 24638 30297
rect 24582 30223 24638 30232
rect 24596 28370 24624 30223
rect 24676 29504 24728 29510
rect 24676 29446 24728 29452
rect 24688 28558 24716 29446
rect 24768 29232 24820 29238
rect 24768 29174 24820 29180
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24596 28342 24716 28370
rect 24504 28206 24624 28234
rect 24492 28144 24544 28150
rect 24492 28086 24544 28092
rect 24398 27024 24454 27033
rect 24398 26959 24454 26968
rect 24412 26382 24440 26959
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24228 24534 24348 24562
rect 24122 24440 24178 24449
rect 24122 24375 24178 24384
rect 24124 23316 24176 23322
rect 24124 23258 24176 23264
rect 24136 22098 24164 23258
rect 24228 22778 24256 24534
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24320 23474 24348 24142
rect 24412 23633 24440 25230
rect 24398 23624 24454 23633
rect 24398 23559 24454 23568
rect 24320 23446 24440 23474
rect 24306 23352 24362 23361
rect 24306 23287 24362 23296
rect 24216 22772 24268 22778
rect 24216 22714 24268 22720
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 23754 21312 23810 21321
rect 23754 21247 23810 21256
rect 23768 21078 23796 21247
rect 23756 21072 23808 21078
rect 23756 21014 23808 21020
rect 24136 20058 24164 22034
rect 24228 21486 24256 22714
rect 24320 22710 24348 23287
rect 24308 22704 24360 22710
rect 24308 22646 24360 22652
rect 24412 22234 24440 23446
rect 24504 23050 24532 28086
rect 24596 27470 24624 28206
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24596 26518 24624 26930
rect 24584 26512 24636 26518
rect 24584 26454 24636 26460
rect 24582 26072 24638 26081
rect 24582 26007 24638 26016
rect 24596 24614 24624 26007
rect 24584 24608 24636 24614
rect 24582 24576 24584 24585
rect 24636 24576 24638 24585
rect 24582 24511 24638 24520
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24492 23044 24544 23050
rect 24492 22986 24544 22992
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24504 22094 24532 22986
rect 24412 22066 24532 22094
rect 24412 21690 24440 22066
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24504 21622 24532 21830
rect 24492 21616 24544 21622
rect 24492 21558 24544 21564
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 24228 21078 24256 21422
rect 24216 21072 24268 21078
rect 24216 21014 24268 21020
rect 24596 20942 24624 23666
rect 24688 23050 24716 28342
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24780 22794 24808 29174
rect 24872 28506 24900 31282
rect 25261 31036 25569 31045
rect 25261 31034 25267 31036
rect 25323 31034 25347 31036
rect 25403 31034 25427 31036
rect 25483 31034 25507 31036
rect 25563 31034 25569 31036
rect 25323 30982 25325 31034
rect 25505 30982 25507 31034
rect 25261 30980 25267 30982
rect 25323 30980 25347 30982
rect 25403 30980 25427 30982
rect 25483 30980 25507 30982
rect 25563 30980 25569 30982
rect 25261 30971 25569 30980
rect 25044 30592 25096 30598
rect 25044 30534 25096 30540
rect 25056 30394 25084 30534
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 25228 30388 25280 30394
rect 25228 30330 25280 30336
rect 25240 30297 25268 30330
rect 25226 30288 25282 30297
rect 25226 30223 25282 30232
rect 25134 30152 25190 30161
rect 25134 30087 25190 30096
rect 25688 30116 25740 30122
rect 25044 30048 25096 30054
rect 25042 30016 25044 30025
rect 25096 30016 25098 30025
rect 25042 29951 25098 29960
rect 25148 29730 25176 30087
rect 25688 30058 25740 30064
rect 25261 29948 25569 29957
rect 25261 29946 25267 29948
rect 25323 29946 25347 29948
rect 25403 29946 25427 29948
rect 25483 29946 25507 29948
rect 25563 29946 25569 29948
rect 25323 29894 25325 29946
rect 25505 29894 25507 29946
rect 25261 29892 25267 29894
rect 25323 29892 25347 29894
rect 25403 29892 25427 29894
rect 25483 29892 25507 29894
rect 25563 29892 25569 29894
rect 25261 29883 25569 29892
rect 25148 29702 25268 29730
rect 25136 29572 25188 29578
rect 25136 29514 25188 29520
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 24952 29028 25004 29034
rect 24952 28970 25004 28976
rect 24964 28937 24992 28970
rect 24950 28928 25006 28937
rect 24950 28863 25006 28872
rect 24872 28478 24992 28506
rect 24964 28422 24992 28478
rect 24952 28416 25004 28422
rect 24952 28358 25004 28364
rect 24952 28008 25004 28014
rect 24952 27950 25004 27956
rect 24860 27668 24912 27674
rect 24860 27610 24912 27616
rect 24872 26246 24900 27610
rect 24964 26761 24992 27950
rect 25056 27878 25084 29446
rect 25148 29306 25176 29514
rect 25136 29300 25188 29306
rect 25136 29242 25188 29248
rect 25240 29050 25268 29702
rect 25148 29022 25268 29050
rect 25044 27872 25096 27878
rect 25044 27814 25096 27820
rect 25042 27704 25098 27713
rect 25042 27639 25098 27648
rect 25056 27402 25084 27639
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 25148 27130 25176 29022
rect 25261 28860 25569 28869
rect 25261 28858 25267 28860
rect 25323 28858 25347 28860
rect 25403 28858 25427 28860
rect 25483 28858 25507 28860
rect 25563 28858 25569 28860
rect 25323 28806 25325 28858
rect 25505 28806 25507 28858
rect 25261 28804 25267 28806
rect 25323 28804 25347 28806
rect 25403 28804 25427 28806
rect 25483 28804 25507 28806
rect 25563 28804 25569 28806
rect 25261 28795 25569 28804
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 25412 28552 25464 28558
rect 25410 28520 25412 28529
rect 25464 28520 25466 28529
rect 25410 28455 25466 28464
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 25240 27946 25268 28358
rect 25516 28014 25544 28698
rect 25596 28416 25648 28422
rect 25596 28358 25648 28364
rect 25504 28008 25556 28014
rect 25318 27976 25374 27985
rect 25228 27940 25280 27946
rect 25318 27911 25374 27920
rect 25502 27976 25504 27985
rect 25556 27976 25558 27985
rect 25502 27911 25558 27920
rect 25228 27882 25280 27888
rect 25332 27878 25360 27911
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 25502 27160 25558 27169
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 25136 27124 25188 27130
rect 25502 27095 25558 27104
rect 25136 27066 25188 27072
rect 25056 26790 25084 27066
rect 25228 26920 25280 26926
rect 25226 26888 25228 26897
rect 25280 26888 25282 26897
rect 25516 26858 25544 27095
rect 25608 26994 25636 28358
rect 25700 27674 25728 30058
rect 25688 27668 25740 27674
rect 25688 27610 25740 27616
rect 25686 27568 25742 27577
rect 25686 27503 25742 27512
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25700 26926 25728 27503
rect 25688 26920 25740 26926
rect 25792 26897 25820 33238
rect 25962 33200 26018 34000
rect 27066 33200 27122 34000
rect 28170 33200 28226 34000
rect 28276 33238 28488 33266
rect 26884 31952 26936 31958
rect 26884 31894 26936 31900
rect 26700 31340 26752 31346
rect 26700 31282 26752 31288
rect 26148 31272 26200 31278
rect 26148 31214 26200 31220
rect 26422 31240 26478 31249
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25976 30938 26004 31078
rect 25964 30932 26016 30938
rect 25964 30874 26016 30880
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 25976 29646 26004 30670
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25976 29345 26004 29582
rect 25962 29336 26018 29345
rect 25962 29271 26018 29280
rect 25964 29096 26016 29102
rect 25964 29038 26016 29044
rect 25872 27668 25924 27674
rect 25872 27610 25924 27616
rect 25884 27441 25912 27610
rect 25870 27432 25926 27441
rect 25870 27367 25926 27376
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25884 26994 25912 27066
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 25688 26862 25740 26868
rect 25778 26888 25834 26897
rect 25226 26823 25282 26832
rect 25504 26852 25556 26858
rect 25778 26823 25834 26832
rect 25504 26794 25556 26800
rect 25044 26784 25096 26790
rect 24950 26752 25006 26761
rect 25044 26726 25096 26732
rect 24950 26687 25006 26696
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25686 26616 25742 26625
rect 25608 26574 25686 26602
rect 25608 26466 25636 26574
rect 25686 26551 25742 26560
rect 25148 26438 25636 26466
rect 24860 26240 24912 26246
rect 24860 26182 24912 26188
rect 25044 26240 25096 26246
rect 25148 26217 25176 26438
rect 25884 26330 25912 26930
rect 25976 26625 26004 29038
rect 26160 28422 26188 31214
rect 26422 31175 26478 31184
rect 26436 31142 26464 31175
rect 26424 31136 26476 31142
rect 26424 31078 26476 31084
rect 26424 30592 26476 30598
rect 26424 30534 26476 30540
rect 26436 30433 26464 30534
rect 26422 30424 26478 30433
rect 26712 30376 26740 31282
rect 26422 30359 26478 30368
rect 26528 30348 26740 30376
rect 26528 29322 26556 30348
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 26344 29294 26556 29322
rect 26344 28994 26372 29294
rect 26252 28966 26372 28994
rect 26148 28416 26200 28422
rect 26148 28358 26200 28364
rect 26148 28008 26200 28014
rect 26148 27950 26200 27956
rect 26056 27872 26108 27878
rect 26056 27814 26108 27820
rect 26068 27674 26096 27814
rect 26056 27668 26108 27674
rect 26056 27610 26108 27616
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 25962 26616 26018 26625
rect 25962 26551 26018 26560
rect 26068 26466 26096 27406
rect 26160 26489 26188 27950
rect 25608 26314 25912 26330
rect 25596 26308 25912 26314
rect 25648 26302 25912 26308
rect 25596 26250 25648 26256
rect 25044 26182 25096 26188
rect 25134 26208 25190 26217
rect 24858 25528 24914 25537
rect 24858 25463 24860 25472
rect 24912 25463 24914 25472
rect 24860 25434 24912 25440
rect 24950 25392 25006 25401
rect 24860 25356 24912 25362
rect 24950 25327 25006 25336
rect 24860 25298 24912 25304
rect 24872 24410 24900 25298
rect 24964 25158 24992 25327
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 24964 24818 24992 25094
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24950 24712 25006 24721
rect 24950 24647 25006 24656
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 24872 23798 24900 24346
rect 24964 24274 24992 24647
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 25056 23322 25084 26182
rect 25134 26143 25190 26152
rect 25318 26208 25374 26217
rect 25318 26143 25374 26152
rect 25226 26072 25282 26081
rect 25226 26007 25282 26016
rect 25240 25906 25268 26007
rect 25228 25900 25280 25906
rect 25228 25842 25280 25848
rect 25332 25786 25360 26143
rect 25884 25906 25912 26302
rect 25976 26450 26096 26466
rect 26146 26480 26202 26489
rect 25976 26444 26108 26450
rect 25976 26438 26056 26444
rect 25872 25900 25924 25906
rect 25872 25842 25924 25848
rect 25148 25758 25360 25786
rect 25780 25764 25832 25770
rect 25148 25537 25176 25758
rect 25780 25706 25832 25712
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25134 25528 25190 25537
rect 25261 25531 25569 25540
rect 25134 25463 25190 25472
rect 25226 25392 25282 25401
rect 25226 25327 25282 25336
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25148 24313 25176 25162
rect 25240 24818 25268 25327
rect 25596 24880 25648 24886
rect 25596 24822 25648 24828
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25608 24392 25636 24822
rect 25792 24721 25820 25706
rect 25870 25528 25926 25537
rect 25870 25463 25926 25472
rect 25884 24993 25912 25463
rect 25976 25294 26004 26438
rect 26146 26415 26202 26424
rect 26056 26386 26108 26392
rect 26056 26308 26108 26314
rect 26056 26250 26108 26256
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26068 26042 26096 26250
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 25964 25288 26016 25294
rect 25964 25230 26016 25236
rect 26160 25106 26188 26250
rect 26252 26246 26280 28966
rect 26516 28484 26568 28490
rect 26516 28426 26568 28432
rect 26332 28144 26384 28150
rect 26332 28086 26384 28092
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 25976 25078 26188 25106
rect 25870 24984 25926 24993
rect 25976 24954 26004 25078
rect 25870 24919 25926 24928
rect 25964 24948 26016 24954
rect 25964 24890 26016 24896
rect 26148 24880 26200 24886
rect 26148 24822 26200 24828
rect 25778 24712 25834 24721
rect 25778 24647 25834 24656
rect 25964 24676 26016 24682
rect 25792 24449 25820 24647
rect 25964 24618 26016 24624
rect 25516 24364 25636 24392
rect 25778 24440 25834 24449
rect 25778 24375 25834 24384
rect 25134 24304 25190 24313
rect 25134 24239 25190 24248
rect 25410 24304 25466 24313
rect 25410 24239 25466 24248
rect 25148 24041 25176 24239
rect 25134 24032 25190 24041
rect 25134 23967 25190 23976
rect 25424 23746 25452 24239
rect 25516 23866 25544 24364
rect 25976 24290 26004 24618
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 25700 24262 26004 24290
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 25608 23905 25636 24074
rect 25594 23896 25650 23905
rect 25504 23860 25556 23866
rect 25594 23831 25650 23840
rect 25504 23802 25556 23808
rect 25424 23718 25636 23746
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 24952 22976 25004 22982
rect 25240 22930 25268 23258
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25004 22924 25268 22930
rect 24952 22918 25268 22924
rect 24964 22902 25268 22918
rect 25424 22817 25452 22986
rect 24688 22766 24808 22794
rect 25410 22808 25466 22817
rect 24688 22409 24716 22766
rect 25410 22743 25466 22752
rect 25516 22710 25544 22986
rect 25504 22704 25556 22710
rect 25504 22646 25556 22652
rect 25608 22574 25636 23718
rect 25700 23254 25728 24262
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 25872 23248 25924 23254
rect 25872 23190 25924 23196
rect 25778 22808 25834 22817
rect 25778 22743 25780 22752
rect 25832 22743 25834 22752
rect 25780 22714 25832 22720
rect 25884 22681 25912 23190
rect 25870 22672 25926 22681
rect 25870 22607 25926 22616
rect 24952 22568 25004 22574
rect 24952 22510 25004 22516
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 24674 22400 24730 22409
rect 24674 22335 24730 22344
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24688 21010 24716 21830
rect 24858 21448 24914 21457
rect 24858 21383 24914 21392
rect 24872 21146 24900 21383
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24780 20602 24808 21014
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24872 20534 24900 20946
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23584 18834 23612 18906
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 23584 17270 23612 18770
rect 23676 18426 23704 19450
rect 23768 18902 23796 19994
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 24872 18086 24900 19178
rect 24964 18970 24992 22510
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25136 21616 25188 21622
rect 25136 21558 25188 21564
rect 25148 21146 25176 21558
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25792 21146 25820 22374
rect 25870 22264 25926 22273
rect 25870 22199 25872 22208
rect 25924 22199 25926 22208
rect 25872 22170 25924 22176
rect 25976 21690 26004 24142
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 25594 20360 25650 20369
rect 25594 20295 25650 20304
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 23572 17264 23624 17270
rect 23572 17206 23624 17212
rect 24872 16794 24900 18022
rect 25056 17338 25084 18362
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25608 17882 25636 20295
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25700 18086 25728 18566
rect 25688 18080 25740 18086
rect 25688 18022 25740 18028
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25504 17808 25556 17814
rect 25504 17750 25556 17756
rect 25516 17338 25544 17750
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 25700 16726 25728 18022
rect 25792 17882 25820 19926
rect 25976 19718 26004 20198
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25976 18358 26004 19654
rect 26068 19446 26096 24550
rect 26160 22234 26188 24822
rect 26252 24070 26280 25298
rect 26344 24993 26372 28086
rect 26424 27872 26476 27878
rect 26424 27814 26476 27820
rect 26436 26926 26464 27814
rect 26424 26920 26476 26926
rect 26424 26862 26476 26868
rect 26422 26344 26478 26353
rect 26422 26279 26478 26288
rect 26330 24984 26386 24993
rect 26330 24919 26386 24928
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 26344 24206 26372 24618
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 26436 24138 26464 26279
rect 26528 25945 26556 28426
rect 26620 26994 26648 30194
rect 26700 30184 26752 30190
rect 26700 30126 26752 30132
rect 26712 29034 26740 30126
rect 26896 29306 26924 31894
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 26884 29300 26936 29306
rect 26884 29242 26936 29248
rect 26700 29028 26752 29034
rect 26700 28970 26752 28976
rect 26884 29028 26936 29034
rect 26884 28970 26936 28976
rect 26896 28150 26924 28970
rect 26884 28144 26936 28150
rect 26884 28086 26936 28092
rect 26792 27940 26844 27946
rect 26792 27882 26844 27888
rect 26698 27840 26754 27849
rect 26698 27775 26754 27784
rect 26608 26988 26660 26994
rect 26608 26930 26660 26936
rect 26606 26888 26662 26897
rect 26606 26823 26608 26832
rect 26660 26823 26662 26832
rect 26608 26794 26660 26800
rect 26620 25974 26648 26794
rect 26608 25968 26660 25974
rect 26514 25936 26570 25945
rect 26608 25910 26660 25916
rect 26514 25871 26570 25880
rect 26712 25378 26740 27775
rect 26804 27402 26832 27882
rect 26792 27396 26844 27402
rect 26792 27338 26844 27344
rect 26884 25900 26936 25906
rect 26884 25842 26936 25848
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26528 25350 26740 25378
rect 26528 24886 26556 25350
rect 26606 25256 26662 25265
rect 26606 25191 26608 25200
rect 26660 25191 26662 25200
rect 26608 25162 26660 25168
rect 26516 24880 26568 24886
rect 26516 24822 26568 24828
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 26516 24132 26568 24138
rect 26516 24074 26568 24080
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26332 24064 26384 24070
rect 26332 24006 26384 24012
rect 26238 23896 26294 23905
rect 26238 23831 26294 23840
rect 26252 23730 26280 23831
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 26252 23118 26280 23666
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26252 22953 26280 23054
rect 26238 22944 26294 22953
rect 26238 22879 26294 22888
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 26160 19514 26188 21558
rect 26252 19718 26280 22714
rect 26344 21622 26372 24006
rect 26528 23712 26556 24074
rect 26436 23684 26556 23712
rect 26436 22982 26464 23684
rect 26620 23610 26648 25162
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 26528 23582 26648 23610
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26332 21616 26384 21622
rect 26332 21558 26384 21564
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 26344 20262 26372 21082
rect 26436 20602 26464 22918
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26056 19440 26108 19446
rect 26056 19382 26108 19388
rect 26528 18426 26556 23582
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26620 23118 26648 23462
rect 26608 23112 26660 23118
rect 26608 23054 26660 23060
rect 26712 22710 26740 24822
rect 26804 24410 26832 25774
rect 26896 24818 26924 25842
rect 26988 25498 27016 30194
rect 27080 27402 27108 33200
rect 28184 33130 28212 33200
rect 28276 33130 28304 33238
rect 28184 33102 28304 33130
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 28172 31476 28224 31482
rect 28172 31418 28224 31424
rect 28184 31385 28212 31418
rect 28170 31376 28226 31385
rect 27252 31340 27304 31346
rect 27252 31282 27304 31288
rect 27896 31340 27948 31346
rect 28368 31346 28396 31622
rect 28170 31311 28226 31320
rect 28356 31340 28408 31346
rect 27896 31282 27948 31288
rect 28356 31282 28408 31288
rect 27158 30832 27214 30841
rect 27158 30767 27214 30776
rect 27172 30394 27200 30767
rect 27160 30388 27212 30394
rect 27160 30330 27212 30336
rect 27160 29164 27212 29170
rect 27160 29106 27212 29112
rect 27068 27396 27120 27402
rect 27068 27338 27120 27344
rect 27172 27146 27200 29106
rect 27080 27118 27200 27146
rect 27264 27146 27292 31282
rect 27344 30388 27396 30394
rect 27528 30388 27580 30394
rect 27344 30330 27396 30336
rect 27448 30348 27528 30376
rect 27356 28257 27384 30330
rect 27342 28248 27398 28257
rect 27342 28183 27398 28192
rect 27448 28121 27476 30348
rect 27908 30374 27936 31282
rect 28080 30728 28132 30734
rect 28080 30670 28132 30676
rect 27528 30330 27580 30336
rect 27724 30346 27936 30374
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27540 29170 27568 30194
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27620 29164 27672 29170
rect 27620 29106 27672 29112
rect 27540 28665 27568 29106
rect 27632 29073 27660 29106
rect 27618 29064 27674 29073
rect 27618 28999 27674 29008
rect 27526 28656 27582 28665
rect 27526 28591 27582 28600
rect 27434 28112 27490 28121
rect 27344 28076 27396 28082
rect 27434 28047 27490 28056
rect 27620 28076 27672 28082
rect 27344 28018 27396 28024
rect 27620 28018 27672 28024
rect 27356 27334 27384 28018
rect 27436 27940 27488 27946
rect 27436 27882 27488 27888
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 27264 27118 27384 27146
rect 26976 25492 27028 25498
rect 26976 25434 27028 25440
rect 27080 24954 27108 27118
rect 27158 27024 27214 27033
rect 27158 26959 27214 26968
rect 27252 26988 27304 26994
rect 27172 26926 27200 26959
rect 27252 26930 27304 26936
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27160 26308 27212 26314
rect 27160 26250 27212 26256
rect 27172 25974 27200 26250
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 27158 25800 27214 25809
rect 27158 25735 27160 25744
rect 27212 25735 27214 25744
rect 27160 25706 27212 25712
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 27068 24948 27120 24954
rect 27068 24890 27120 24896
rect 27172 24854 27200 25094
rect 26988 24826 27200 24854
rect 26884 24812 26936 24818
rect 26884 24754 26936 24760
rect 26792 24404 26844 24410
rect 26792 24346 26844 24352
rect 26792 24064 26844 24070
rect 26792 24006 26844 24012
rect 26804 23254 26832 24006
rect 26896 23633 26924 24754
rect 26988 24750 27016 24826
rect 26976 24744 27028 24750
rect 26976 24686 27028 24692
rect 26988 23730 27016 24686
rect 27264 24614 27292 26930
rect 27356 25362 27384 27118
rect 27344 25356 27396 25362
rect 27344 25298 27396 25304
rect 27342 24984 27398 24993
rect 27342 24919 27398 24928
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27252 24608 27304 24614
rect 27252 24550 27304 24556
rect 27068 24404 27120 24410
rect 27068 24346 27120 24352
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26882 23624 26938 23633
rect 26882 23559 26938 23568
rect 26792 23248 26844 23254
rect 26792 23190 26844 23196
rect 26896 23066 26924 23559
rect 26988 23089 27016 23666
rect 27080 23594 27108 24346
rect 27172 24177 27200 24550
rect 27264 24313 27292 24550
rect 27250 24304 27306 24313
rect 27250 24239 27306 24248
rect 27158 24168 27214 24177
rect 27158 24103 27214 24112
rect 27158 24032 27214 24041
rect 27158 23967 27214 23976
rect 27068 23588 27120 23594
rect 27068 23530 27120 23536
rect 27172 23322 27200 23967
rect 27160 23316 27212 23322
rect 27160 23258 27212 23264
rect 27066 23216 27122 23225
rect 27066 23151 27122 23160
rect 27080 23118 27108 23151
rect 27068 23112 27120 23118
rect 26804 23038 26924 23066
rect 26974 23080 27030 23089
rect 26804 22778 26832 23038
rect 27068 23054 27120 23060
rect 26974 23015 27030 23024
rect 26884 22976 26936 22982
rect 26884 22918 26936 22924
rect 26792 22772 26844 22778
rect 26792 22714 26844 22720
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 26896 22642 26924 22918
rect 26884 22636 26936 22642
rect 26884 22578 26936 22584
rect 26988 20714 27016 23015
rect 27172 22438 27200 23258
rect 27160 22432 27212 22438
rect 27160 22374 27212 22380
rect 27252 22432 27304 22438
rect 27252 22374 27304 22380
rect 27264 21622 27292 22374
rect 27356 22234 27384 24919
rect 27448 24750 27476 27882
rect 27528 27328 27580 27334
rect 27528 27270 27580 27276
rect 27540 26994 27568 27270
rect 27632 26994 27660 28018
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27632 26897 27660 26930
rect 27618 26888 27674 26897
rect 27528 26852 27580 26858
rect 27618 26823 27674 26832
rect 27528 26794 27580 26800
rect 27540 26081 27568 26794
rect 27724 26217 27752 30346
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 27802 29200 27858 29209
rect 27802 29135 27804 29144
rect 27856 29135 27858 29144
rect 27804 29106 27856 29112
rect 28000 28994 28028 29446
rect 27908 28966 28028 28994
rect 27804 28416 27856 28422
rect 27804 28358 27856 28364
rect 27816 28218 27844 28358
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 27804 28076 27856 28082
rect 27804 28018 27856 28024
rect 27816 27985 27844 28018
rect 27802 27976 27858 27985
rect 27802 27911 27858 27920
rect 27908 27674 27936 28966
rect 27988 28144 28040 28150
rect 27988 28086 28040 28092
rect 27896 27668 27948 27674
rect 27896 27610 27948 27616
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27710 26208 27766 26217
rect 27710 26143 27766 26152
rect 27526 26072 27582 26081
rect 27526 26007 27582 26016
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27540 25226 27568 25842
rect 27724 25362 27752 26143
rect 27908 25922 27936 27338
rect 28000 26042 28028 28086
rect 28092 26994 28120 30670
rect 28264 30592 28316 30598
rect 28264 30534 28316 30540
rect 28276 29646 28304 30534
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 28356 28960 28408 28966
rect 28356 28902 28408 28908
rect 28170 28520 28226 28529
rect 28170 28455 28226 28464
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 28184 26738 28212 28455
rect 28368 28422 28396 28902
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28264 27872 28316 27878
rect 28264 27814 28316 27820
rect 28276 27305 28304 27814
rect 28368 27334 28396 28358
rect 28356 27328 28408 27334
rect 28262 27296 28318 27305
rect 28356 27270 28408 27276
rect 28262 27231 28318 27240
rect 28184 26710 28304 26738
rect 27988 26036 28040 26042
rect 27988 25978 28040 25984
rect 27804 25900 27856 25906
rect 27908 25894 28120 25922
rect 27804 25842 27856 25848
rect 27816 25401 27844 25842
rect 27894 25800 27950 25809
rect 27894 25735 27950 25744
rect 27802 25392 27858 25401
rect 27712 25356 27764 25362
rect 27802 25327 27858 25336
rect 27712 25298 27764 25304
rect 27816 25294 27844 25327
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27528 25220 27580 25226
rect 27528 25162 27580 25168
rect 27526 25120 27582 25129
rect 27526 25055 27582 25064
rect 27540 24886 27568 25055
rect 27528 24880 27580 24886
rect 27528 24822 27580 24828
rect 27436 24744 27488 24750
rect 27436 24686 27488 24692
rect 27436 24608 27488 24614
rect 27436 24550 27488 24556
rect 27448 23798 27476 24550
rect 27526 24304 27582 24313
rect 27526 24239 27582 24248
rect 27540 24206 27568 24239
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 27540 23866 27568 24142
rect 27632 24070 27660 25230
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 27710 24848 27766 24857
rect 27816 24818 27844 25094
rect 27710 24783 27766 24792
rect 27804 24812 27856 24818
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27356 22030 27384 22170
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27252 21616 27304 21622
rect 27252 21558 27304 21564
rect 26896 20686 27016 20714
rect 26896 18630 26924 20686
rect 27264 20602 27292 21558
rect 27252 20596 27304 20602
rect 27252 20538 27304 20544
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26884 18624 26936 18630
rect 26884 18566 26936 18572
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 26896 16794 26924 18566
rect 26988 17882 27016 20198
rect 27540 20058 27568 21966
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 26976 17876 27028 17882
rect 26976 17818 27028 17824
rect 27172 17338 27200 19654
rect 27632 18426 27660 23666
rect 27724 23322 27752 24783
rect 27804 24754 27856 24760
rect 27816 24410 27844 24754
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27710 22128 27766 22137
rect 27710 22063 27766 22072
rect 27724 22030 27752 22063
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 27816 17882 27844 24074
rect 27908 22642 27936 25735
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 28000 24342 28028 25230
rect 27988 24336 28040 24342
rect 27988 24278 28040 24284
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 28092 21554 28120 25894
rect 28170 24440 28226 24449
rect 28170 24375 28226 24384
rect 28184 23798 28212 24375
rect 28276 24138 28304 26710
rect 28368 26586 28396 27270
rect 28356 26580 28408 26586
rect 28356 26522 28408 26528
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 28368 25430 28396 25842
rect 28356 25424 28408 25430
rect 28356 25366 28408 25372
rect 28264 24132 28316 24138
rect 28264 24074 28316 24080
rect 28172 23792 28224 23798
rect 28172 23734 28224 23740
rect 28354 23760 28410 23769
rect 28354 23695 28356 23704
rect 28408 23695 28410 23704
rect 28356 23666 28408 23672
rect 28172 23656 28224 23662
rect 28172 23598 28224 23604
rect 28184 22778 28212 23598
rect 28356 23112 28408 23118
rect 28354 23080 28356 23089
rect 28408 23080 28410 23089
rect 28354 23015 28410 23024
rect 28172 22772 28224 22778
rect 28172 22714 28224 22720
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28276 22409 28304 22578
rect 28262 22400 28318 22409
rect 28262 22335 28318 22344
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 28276 19514 28304 22335
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28368 21593 28396 21966
rect 28354 21584 28410 21593
rect 28354 21519 28410 21528
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28368 21049 28396 21286
rect 28460 21078 28488 33238
rect 29274 33200 29330 34000
rect 29288 31770 29316 33200
rect 29288 31742 29408 31770
rect 28734 31580 29042 31589
rect 28734 31578 28740 31580
rect 28796 31578 28820 31580
rect 28876 31578 28900 31580
rect 28956 31578 28980 31580
rect 29036 31578 29042 31580
rect 28796 31526 28798 31578
rect 28978 31526 28980 31578
rect 28734 31524 28740 31526
rect 28796 31524 28820 31526
rect 28876 31524 28900 31526
rect 28956 31524 28980 31526
rect 29036 31524 29042 31526
rect 28734 31515 29042 31524
rect 28998 31240 29054 31249
rect 29054 31198 29316 31226
rect 28998 31175 29054 31184
rect 28734 30492 29042 30501
rect 28734 30490 28740 30492
rect 28796 30490 28820 30492
rect 28876 30490 28900 30492
rect 28956 30490 28980 30492
rect 29036 30490 29042 30492
rect 28796 30438 28798 30490
rect 28978 30438 28980 30490
rect 28734 30436 28740 30438
rect 28796 30436 28820 30438
rect 28876 30436 28900 30438
rect 28956 30436 28980 30438
rect 29036 30436 29042 30438
rect 28734 30427 29042 30436
rect 28538 29880 28594 29889
rect 28538 29815 28594 29824
rect 28552 22166 28580 29815
rect 28632 29640 28684 29646
rect 28632 29582 28684 29588
rect 28644 28966 28672 29582
rect 28734 29404 29042 29413
rect 28734 29402 28740 29404
rect 28796 29402 28820 29404
rect 28876 29402 28900 29404
rect 28956 29402 28980 29404
rect 29036 29402 29042 29404
rect 28796 29350 28798 29402
rect 28978 29350 28980 29402
rect 28734 29348 28740 29350
rect 28796 29348 28820 29350
rect 28876 29348 28900 29350
rect 28956 29348 28980 29350
rect 29036 29348 29042 29350
rect 28734 29339 29042 29348
rect 28998 29200 29054 29209
rect 29054 29158 29224 29186
rect 28998 29135 29054 29144
rect 28632 28960 28684 28966
rect 28632 28902 28684 28908
rect 28734 28316 29042 28325
rect 28734 28314 28740 28316
rect 28796 28314 28820 28316
rect 28876 28314 28900 28316
rect 28956 28314 28980 28316
rect 29036 28314 29042 28316
rect 28796 28262 28798 28314
rect 28978 28262 28980 28314
rect 28734 28260 28740 28262
rect 28796 28260 28820 28262
rect 28876 28260 28900 28262
rect 28956 28260 28980 28262
rect 29036 28260 29042 28262
rect 28734 28251 29042 28260
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28630 27024 28686 27033
rect 28630 26959 28686 26968
rect 28644 22574 28672 26959
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 28632 22568 28684 22574
rect 28632 22510 28684 22516
rect 28540 22160 28592 22166
rect 28540 22102 28592 22108
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 29196 21146 29224 29158
rect 29184 21140 29236 21146
rect 29184 21082 29236 21088
rect 28448 21072 28500 21078
rect 28354 21040 28410 21049
rect 28448 21014 28500 21020
rect 29288 21010 29316 31198
rect 29380 22438 29408 31742
rect 29460 25968 29512 25974
rect 29460 25910 29512 25916
rect 29368 22432 29420 22438
rect 29368 22374 29420 22380
rect 28354 20975 28410 20984
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 29472 20602 29500 25910
rect 29460 20596 29512 20602
rect 29460 20538 29512 20544
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 28368 20369 28396 20402
rect 28354 20360 28410 20369
rect 28354 20295 28410 20304
rect 28368 20058 28396 20295
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28356 19848 28408 19854
rect 28354 19816 28356 19825
rect 28408 19816 28410 19825
rect 28354 19751 28410 19760
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28368 19009 28396 19110
rect 28354 19000 28410 19009
rect 28354 18935 28410 18944
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28368 18358 28396 18702
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28356 18352 28408 18358
rect 28354 18320 28356 18329
rect 28408 18320 28410 18329
rect 28354 18255 28410 18264
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 28356 17672 28408 17678
rect 28354 17640 28356 17649
rect 28408 17640 28410 17649
rect 28354 17575 28410 17584
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 28356 16992 28408 16998
rect 28354 16960 28356 16969
rect 28408 16960 28410 16969
rect 28354 16895 28410 16904
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 25688 16720 25740 16726
rect 25688 16662 25740 16668
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 1584 16040 1636 16046
rect 1582 16008 1584 16017
rect 1636 16008 1638 16017
rect 1582 15943 1638 15952
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 28368 15609 28396 15846
rect 28354 15600 28410 15609
rect 28354 15535 28410 15544
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 15337 1624 15438
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28354 14920 28410 14929
rect 28354 14855 28356 14864
rect 28408 14855 28410 14864
rect 28356 14826 28408 14832
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13977 1624 14350
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 28356 13728 28408 13734
rect 28356 13670 28408 13676
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 28368 13569 28396 13670
rect 28354 13560 28410 13569
rect 28354 13495 28410 13504
rect 1584 13320 1636 13326
rect 1582 13288 1584 13297
rect 28356 13320 28408 13326
rect 1636 13288 1638 13297
rect 28356 13262 28408 13268
rect 1582 13223 1638 13232
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 28368 12889 28396 13262
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28354 12880 28410 12889
rect 28354 12815 28410 12824
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11937 1624 12174
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 1582 11928 1638 11937
rect 7896 11931 8204 11940
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 1582 11863 1638 11872
rect 1584 11552 1636 11558
rect 28356 11552 28408 11558
rect 1584 11494 1636 11500
rect 28354 11520 28356 11529
rect 28408 11520 28410 11529
rect 1596 11257 1624 11494
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 25261 11452 25569 11461
rect 28354 11455 28410 11464
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 1582 11248 1638 11257
rect 1582 11183 1638 11192
rect 28356 11144 28408 11150
rect 28354 11112 28356 11121
rect 28408 11112 28410 11121
rect 28354 11047 28410 11056
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9897 1624 9998
rect 1582 9888 1638 9897
rect 1582 9823 1638 9832
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28354 9480 28410 9489
rect 28354 9415 28356 9424
rect 28408 9415 28410 9424
rect 28356 9386 28408 9392
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9217 1624 9318
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 1582 9208 1638 9217
rect 4423 9211 4731 9220
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 1582 9143 1638 9152
rect 28356 9104 28408 9110
rect 28354 9072 28356 9081
rect 28408 9072 28410 9081
rect 28354 9007 28410 9016
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 1584 7880 1636 7886
rect 1582 7848 1584 7857
rect 28356 7880 28408 7886
rect 1636 7848 1638 7857
rect 28356 7822 28408 7828
rect 1582 7783 1638 7792
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 28368 7449 28396 7822
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 28354 7440 28410 7449
rect 28354 7375 28410 7384
rect 1584 7200 1636 7206
rect 1582 7168 1584 7177
rect 1636 7168 1638 7177
rect 1582 7103 1638 7112
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 28356 6792 28408 6798
rect 28354 6760 28356 6769
rect 28408 6760 28410 6769
rect 28354 6695 28410 6704
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5817 1624 6054
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 1582 5808 1638 5817
rect 1582 5743 1638 5752
rect 28356 5704 28408 5710
rect 28354 5672 28356 5681
rect 28408 5672 28410 5681
rect 28354 5607 28410 5616
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 1584 5160 1636 5166
rect 1582 5128 1584 5137
rect 1636 5128 1638 5137
rect 1582 5063 1638 5072
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 28368 4729 28396 4966
rect 28354 4720 28410 4729
rect 28354 4655 28410 4664
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3777 1624 3878
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 1582 3768 1638 3777
rect 4423 3771 4731 3780
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 1582 3703 1638 3712
rect 28356 3664 28408 3670
rect 28354 3632 28356 3641
rect 28408 3632 28410 3641
rect 28354 3567 28410 3576
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 3097 1624 3470
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 28368 2689 28396 2790
rect 28354 2680 28410 2689
rect 28354 2615 28410 2624
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
<< via2 >>
rect 7902 31578 7958 31580
rect 7982 31578 8038 31580
rect 8062 31578 8118 31580
rect 8142 31578 8198 31580
rect 7902 31526 7948 31578
rect 7948 31526 7958 31578
rect 7982 31526 8012 31578
rect 8012 31526 8024 31578
rect 8024 31526 8038 31578
rect 8062 31526 8076 31578
rect 8076 31526 8088 31578
rect 8088 31526 8118 31578
rect 8142 31526 8152 31578
rect 8152 31526 8198 31578
rect 7902 31524 7958 31526
rect 7982 31524 8038 31526
rect 8062 31524 8118 31526
rect 8142 31524 8198 31526
rect 4429 31034 4485 31036
rect 4509 31034 4565 31036
rect 4589 31034 4645 31036
rect 4669 31034 4725 31036
rect 4429 30982 4475 31034
rect 4475 30982 4485 31034
rect 4509 30982 4539 31034
rect 4539 30982 4551 31034
rect 4551 30982 4565 31034
rect 4589 30982 4603 31034
rect 4603 30982 4615 31034
rect 4615 30982 4645 31034
rect 4669 30982 4679 31034
rect 4679 30982 4725 31034
rect 4429 30980 4485 30982
rect 4509 30980 4565 30982
rect 4589 30980 4645 30982
rect 4669 30980 4725 30982
rect 5354 30640 5410 30696
rect 1582 30232 1638 30288
rect 4429 29946 4485 29948
rect 4509 29946 4565 29948
rect 4589 29946 4645 29948
rect 4669 29946 4725 29948
rect 4429 29894 4475 29946
rect 4475 29894 4485 29946
rect 4509 29894 4539 29946
rect 4539 29894 4551 29946
rect 4551 29894 4565 29946
rect 4589 29894 4603 29946
rect 4603 29894 4615 29946
rect 4615 29894 4645 29946
rect 4669 29894 4679 29946
rect 4679 29894 4725 29946
rect 4429 29892 4485 29894
rect 4509 29892 4565 29894
rect 4589 29892 4645 29894
rect 4669 29892 4725 29894
rect 6550 30232 6606 30288
rect 1582 29588 1584 29608
rect 1584 29588 1636 29608
rect 1636 29588 1638 29608
rect 1582 29552 1638 29588
rect 4429 28858 4485 28860
rect 4509 28858 4565 28860
rect 4589 28858 4645 28860
rect 4669 28858 4725 28860
rect 4429 28806 4475 28858
rect 4475 28806 4485 28858
rect 4509 28806 4539 28858
rect 4539 28806 4551 28858
rect 4551 28806 4565 28858
rect 4589 28806 4603 28858
rect 4603 28806 4615 28858
rect 4615 28806 4645 28858
rect 4669 28806 4679 28858
rect 4679 28806 4725 28858
rect 4429 28804 4485 28806
rect 4509 28804 4565 28806
rect 4589 28804 4645 28806
rect 4669 28804 4725 28806
rect 1582 28192 1638 28248
rect 7902 30490 7958 30492
rect 7982 30490 8038 30492
rect 8062 30490 8118 30492
rect 8142 30490 8198 30492
rect 7902 30438 7948 30490
rect 7948 30438 7958 30490
rect 7982 30438 8012 30490
rect 8012 30438 8024 30490
rect 8024 30438 8038 30490
rect 8062 30438 8076 30490
rect 8076 30438 8088 30490
rect 8088 30438 8118 30490
rect 8142 30438 8152 30490
rect 8152 30438 8198 30490
rect 7902 30436 7958 30438
rect 7982 30436 8038 30438
rect 8062 30436 8118 30438
rect 8142 30436 8198 30438
rect 7902 29402 7958 29404
rect 7982 29402 8038 29404
rect 8062 29402 8118 29404
rect 8142 29402 8198 29404
rect 7902 29350 7948 29402
rect 7948 29350 7958 29402
rect 7982 29350 8012 29402
rect 8012 29350 8024 29402
rect 8024 29350 8038 29402
rect 8062 29350 8076 29402
rect 8076 29350 8088 29402
rect 8088 29350 8118 29402
rect 8142 29350 8152 29402
rect 8152 29350 8198 29402
rect 7902 29348 7958 29350
rect 7982 29348 8038 29350
rect 8062 29348 8118 29350
rect 8142 29348 8198 29350
rect 9310 30776 9366 30832
rect 8482 29300 8538 29336
rect 8482 29280 8484 29300
rect 8484 29280 8536 29300
rect 8536 29280 8538 29300
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 7902 28314 7958 28316
rect 7982 28314 8038 28316
rect 8062 28314 8118 28316
rect 8142 28314 8198 28316
rect 7902 28262 7948 28314
rect 7948 28262 7958 28314
rect 7982 28262 8012 28314
rect 8012 28262 8024 28314
rect 8024 28262 8038 28314
rect 8062 28262 8076 28314
rect 8076 28262 8088 28314
rect 8088 28262 8118 28314
rect 8142 28262 8152 28314
rect 8152 28262 8198 28314
rect 7902 28260 7958 28262
rect 7982 28260 8038 28262
rect 8062 28260 8118 28262
rect 8142 28260 8198 28262
rect 1582 27512 1638 27568
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 8298 26968 8354 27024
rect 9586 30232 9642 30288
rect 9770 30116 9826 30152
rect 9770 30096 9772 30116
rect 9772 30096 9824 30116
rect 9824 30096 9826 30116
rect 9770 29688 9826 29744
rect 9402 26968 9458 27024
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 10046 30368 10102 30424
rect 9678 29008 9734 29064
rect 1582 26152 1638 26208
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 1582 25472 1638 25528
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 1582 24148 1584 24168
rect 1584 24148 1636 24168
rect 1636 24148 1638 24168
rect 1582 24112 1638 24148
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 11150 31340 11206 31376
rect 11150 31320 11152 31340
rect 11152 31320 11204 31340
rect 11204 31320 11206 31340
rect 11375 31034 11431 31036
rect 11455 31034 11511 31036
rect 11535 31034 11591 31036
rect 11615 31034 11671 31036
rect 11375 30982 11421 31034
rect 11421 30982 11431 31034
rect 11455 30982 11485 31034
rect 11485 30982 11497 31034
rect 11497 30982 11511 31034
rect 11535 30982 11549 31034
rect 11549 30982 11561 31034
rect 11561 30982 11591 31034
rect 11615 30982 11625 31034
rect 11625 30982 11671 31034
rect 11375 30980 11431 30982
rect 11455 30980 11511 30982
rect 11535 30980 11591 30982
rect 11615 30980 11671 30982
rect 10598 29008 10654 29064
rect 10414 26424 10470 26480
rect 9862 26324 9864 26344
rect 9864 26324 9916 26344
rect 9916 26324 9918 26344
rect 9862 26288 9918 26324
rect 11150 30116 11206 30152
rect 11150 30096 11152 30116
rect 11152 30096 11204 30116
rect 11204 30096 11206 30116
rect 13542 31728 13598 31784
rect 11978 31184 12034 31240
rect 11978 31048 12034 31104
rect 11794 30368 11850 30424
rect 11375 29946 11431 29948
rect 11455 29946 11511 29948
rect 11535 29946 11591 29948
rect 11615 29946 11671 29948
rect 11375 29894 11421 29946
rect 11421 29894 11431 29946
rect 11455 29894 11485 29946
rect 11485 29894 11497 29946
rect 11497 29894 11511 29946
rect 11535 29894 11549 29946
rect 11549 29894 11561 29946
rect 11561 29894 11591 29946
rect 11615 29894 11625 29946
rect 11625 29894 11671 29946
rect 11375 29892 11431 29894
rect 11455 29892 11511 29894
rect 11535 29892 11591 29894
rect 11615 29892 11671 29894
rect 11334 29708 11390 29744
rect 11334 29688 11336 29708
rect 11336 29688 11388 29708
rect 11388 29688 11390 29708
rect 12070 30912 12126 30968
rect 11702 29144 11758 29200
rect 10874 28600 10930 28656
rect 11375 28858 11431 28860
rect 11455 28858 11511 28860
rect 11535 28858 11591 28860
rect 11615 28858 11671 28860
rect 11375 28806 11421 28858
rect 11421 28806 11431 28858
rect 11455 28806 11485 28858
rect 11485 28806 11497 28858
rect 11497 28806 11511 28858
rect 11535 28806 11549 28858
rect 11549 28806 11561 28858
rect 11561 28806 11591 28858
rect 11615 28806 11625 28858
rect 11625 28806 11671 28858
rect 11375 28804 11431 28806
rect 11455 28804 11511 28806
rect 11535 28804 11591 28806
rect 11615 28804 11671 28806
rect 11426 28056 11482 28112
rect 11886 29008 11942 29064
rect 11702 28328 11758 28384
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 13358 31048 13414 31104
rect 12346 28192 12402 28248
rect 12070 27512 12126 27568
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 12530 28500 12532 28520
rect 12532 28500 12584 28520
rect 12584 28500 12586 28520
rect 12530 28464 12586 28500
rect 12530 27648 12586 27704
rect 12438 27376 12494 27432
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 1582 22072 1638 22128
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 12898 29416 12954 29472
rect 13266 29960 13322 30016
rect 13266 29552 13322 29608
rect 13358 29280 13414 29336
rect 12990 28192 13046 28248
rect 12990 26696 13046 26752
rect 12898 25880 12954 25936
rect 13266 28600 13322 28656
rect 13266 27956 13268 27976
rect 13268 27956 13320 27976
rect 13320 27956 13322 27976
rect 13266 27920 13322 27956
rect 13358 27240 13414 27296
rect 13266 26288 13322 26344
rect 13726 29552 13782 29608
rect 13818 28328 13874 28384
rect 14848 31578 14904 31580
rect 14928 31578 14984 31580
rect 15008 31578 15064 31580
rect 15088 31578 15144 31580
rect 14848 31526 14894 31578
rect 14894 31526 14904 31578
rect 14928 31526 14958 31578
rect 14958 31526 14970 31578
rect 14970 31526 14984 31578
rect 15008 31526 15022 31578
rect 15022 31526 15034 31578
rect 15034 31526 15064 31578
rect 15088 31526 15098 31578
rect 15098 31526 15144 31578
rect 14848 31524 14904 31526
rect 14928 31524 14984 31526
rect 15008 31524 15064 31526
rect 15088 31524 15144 31526
rect 15658 31456 15714 31512
rect 14186 30232 14242 30288
rect 14186 29824 14242 29880
rect 14094 29416 14150 29472
rect 14002 25200 14058 25256
rect 13082 24248 13138 24304
rect 14186 27648 14242 27704
rect 14094 24792 14150 24848
rect 14462 29008 14518 29064
rect 14848 30490 14904 30492
rect 14928 30490 14984 30492
rect 15008 30490 15064 30492
rect 15088 30490 15144 30492
rect 14848 30438 14894 30490
rect 14894 30438 14904 30490
rect 14928 30438 14958 30490
rect 14958 30438 14970 30490
rect 14970 30438 14984 30490
rect 15008 30438 15022 30490
rect 15022 30438 15034 30490
rect 15034 30438 15064 30490
rect 15088 30438 15098 30490
rect 15098 30438 15144 30490
rect 14848 30436 14904 30438
rect 14928 30436 14984 30438
rect 15008 30436 15064 30438
rect 15088 30436 15144 30438
rect 15014 29960 15070 30016
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14894 29402
rect 14894 29350 14904 29402
rect 14928 29350 14958 29402
rect 14958 29350 14970 29402
rect 14970 29350 14984 29402
rect 15008 29350 15022 29402
rect 15022 29350 15034 29402
rect 15034 29350 15064 29402
rect 15088 29350 15098 29402
rect 15098 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 15290 30232 15346 30288
rect 15290 28872 15346 28928
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14894 28314
rect 14894 28262 14904 28314
rect 14928 28262 14958 28314
rect 14958 28262 14970 28314
rect 14970 28262 14984 28314
rect 15008 28262 15022 28314
rect 15022 28262 15034 28314
rect 15034 28262 15064 28314
rect 15088 28262 15098 28314
rect 15098 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 14462 27784 14518 27840
rect 14462 27240 14518 27296
rect 14370 26832 14426 26888
rect 15198 27648 15254 27704
rect 15474 28328 15530 28384
rect 15382 28192 15438 28248
rect 15474 27648 15530 27704
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 14646 26308 14702 26344
rect 14646 26288 14648 26308
rect 14648 26288 14700 26308
rect 14700 26288 14702 26308
rect 14830 26696 14886 26752
rect 15106 26560 15162 26616
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 15382 27240 15438 27296
rect 15290 26696 15346 26752
rect 14738 25900 14794 25936
rect 14738 25880 14740 25900
rect 14740 25880 14792 25900
rect 14792 25880 14794 25900
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 15474 26560 15530 26616
rect 14462 24112 14518 24168
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 15750 29416 15806 29472
rect 15750 29280 15806 29336
rect 15750 28872 15806 28928
rect 16210 29824 16266 29880
rect 16026 27240 16082 27296
rect 15934 26696 15990 26752
rect 15934 26560 15990 26616
rect 16118 26560 16174 26616
rect 16118 26152 16174 26208
rect 17130 31592 17186 31648
rect 17958 30912 18014 30968
rect 17498 30640 17554 30696
rect 17682 30676 17684 30696
rect 17684 30676 17736 30696
rect 17736 30676 17738 30696
rect 17682 30640 17738 30676
rect 17590 30368 17646 30424
rect 17130 30232 17186 30288
rect 16762 29280 16818 29336
rect 16302 27104 16358 27160
rect 16486 28328 16542 28384
rect 16578 28192 16634 28248
rect 16762 27104 16818 27160
rect 16670 26560 16726 26616
rect 15658 23568 15714 23624
rect 16486 26152 16542 26208
rect 16394 25608 16450 25664
rect 16118 23976 16174 24032
rect 16762 26016 16818 26072
rect 17130 29824 17186 29880
rect 17038 29008 17094 29064
rect 16854 25880 16910 25936
rect 16578 24656 16634 24712
rect 16486 24520 16542 24576
rect 17314 29824 17370 29880
rect 17222 26016 17278 26072
rect 17406 29008 17462 29064
rect 18234 31592 18290 31648
rect 18321 31034 18377 31036
rect 18401 31034 18457 31036
rect 18481 31034 18537 31036
rect 18561 31034 18617 31036
rect 18321 30982 18367 31034
rect 18367 30982 18377 31034
rect 18401 30982 18431 31034
rect 18431 30982 18443 31034
rect 18443 30982 18457 31034
rect 18481 30982 18495 31034
rect 18495 30982 18507 31034
rect 18507 30982 18537 31034
rect 18561 30982 18571 31034
rect 18571 30982 18617 31034
rect 18321 30980 18377 30982
rect 18401 30980 18457 30982
rect 18481 30980 18537 30982
rect 18561 30980 18617 30982
rect 18694 30912 18750 30968
rect 18142 30640 18198 30696
rect 17958 29960 18014 30016
rect 18050 29824 18106 29880
rect 17866 29416 17922 29472
rect 17958 29280 18014 29336
rect 17866 29144 17922 29200
rect 17498 27648 17554 27704
rect 17406 27240 17462 27296
rect 17222 25236 17224 25256
rect 17224 25236 17276 25256
rect 17276 25236 17278 25256
rect 17222 25200 17278 25236
rect 17222 24656 17278 24712
rect 17038 23704 17094 23760
rect 17314 22924 17316 22944
rect 17316 22924 17368 22944
rect 17368 22924 17370 22944
rect 17314 22888 17370 22924
rect 17498 26288 17554 26344
rect 17498 26152 17554 26208
rect 17774 27648 17830 27704
rect 17682 27240 17738 27296
rect 17958 28872 18014 28928
rect 17958 28736 18014 28792
rect 17958 28328 18014 28384
rect 17774 26696 17830 26752
rect 17866 26560 17922 26616
rect 17866 26288 17922 26344
rect 17682 25608 17738 25664
rect 17498 25472 17554 25528
rect 17774 25472 17830 25528
rect 17682 24792 17738 24848
rect 17590 24520 17646 24576
rect 17682 22888 17738 22944
rect 18050 24656 18106 24712
rect 18050 23432 18106 23488
rect 18321 29946 18377 29948
rect 18401 29946 18457 29948
rect 18481 29946 18537 29948
rect 18561 29946 18617 29948
rect 18321 29894 18367 29946
rect 18367 29894 18377 29946
rect 18401 29894 18431 29946
rect 18431 29894 18443 29946
rect 18443 29894 18457 29946
rect 18481 29894 18495 29946
rect 18495 29894 18507 29946
rect 18507 29894 18537 29946
rect 18561 29894 18571 29946
rect 18571 29894 18617 29946
rect 18321 29892 18377 29894
rect 18401 29892 18457 29894
rect 18481 29892 18537 29894
rect 18561 29892 18617 29894
rect 18694 29452 18696 29472
rect 18696 29452 18748 29472
rect 18748 29452 18750 29472
rect 18694 29416 18750 29452
rect 18326 29280 18382 29336
rect 18510 29280 18566 29336
rect 19062 30368 19118 30424
rect 19154 30096 19210 30152
rect 18786 28872 18842 28928
rect 18321 28858 18377 28860
rect 18401 28858 18457 28860
rect 18481 28858 18537 28860
rect 18561 28858 18617 28860
rect 18321 28806 18367 28858
rect 18367 28806 18377 28858
rect 18401 28806 18431 28858
rect 18431 28806 18443 28858
rect 18443 28806 18457 28858
rect 18481 28806 18495 28858
rect 18495 28806 18507 28858
rect 18507 28806 18537 28858
rect 18561 28806 18571 28858
rect 18571 28806 18617 28858
rect 18321 28804 18377 28806
rect 18401 28804 18457 28806
rect 18481 28804 18537 28806
rect 18561 28804 18617 28806
rect 18694 27784 18750 27840
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 18694 26016 18750 26072
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18694 25472 18750 25528
rect 18694 24792 18750 24848
rect 18510 24692 18512 24712
rect 18512 24692 18564 24712
rect 18564 24692 18566 24712
rect 18510 24656 18566 24692
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 19062 28736 19118 28792
rect 19430 30504 19486 30560
rect 19614 30504 19670 30560
rect 19522 30368 19578 30424
rect 19430 30096 19486 30152
rect 19338 29824 19394 29880
rect 19430 28908 19432 28928
rect 19432 28908 19484 28928
rect 19484 28908 19486 28928
rect 19430 28872 19486 28908
rect 19246 28092 19248 28112
rect 19248 28092 19300 28112
rect 19300 28092 19302 28112
rect 19246 28056 19302 28092
rect 19062 26288 19118 26344
rect 19338 27784 19394 27840
rect 19246 26696 19302 26752
rect 19062 25744 19118 25800
rect 19062 24812 19118 24848
rect 19062 24792 19064 24812
rect 19064 24792 19116 24812
rect 19116 24792 19118 24812
rect 19338 25744 19394 25800
rect 19798 29824 19854 29880
rect 19706 28872 19762 28928
rect 19614 27648 19670 27704
rect 20074 28328 20130 28384
rect 20258 28192 20314 28248
rect 20166 27648 20222 27704
rect 20166 27512 20222 27568
rect 20166 27240 20222 27296
rect 19706 26560 19762 26616
rect 19798 26324 19800 26344
rect 19800 26324 19852 26344
rect 19852 26324 19854 26344
rect 19798 26288 19854 26324
rect 19522 26016 19578 26072
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 18234 22752 18290 22808
rect 17866 22480 17922 22536
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 19430 24384 19486 24440
rect 19706 25064 19762 25120
rect 19798 24384 19854 24440
rect 19614 23568 19670 23624
rect 19522 23432 19578 23488
rect 19522 23024 19578 23080
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 1582 21428 1584 21448
rect 1584 21428 1636 21448
rect 1636 21428 1638 21448
rect 1582 21392 1638 21428
rect 20074 25880 20130 25936
rect 19982 25064 20038 25120
rect 20166 25064 20222 25120
rect 19706 23296 19762 23352
rect 20074 24520 20130 24576
rect 19982 22752 20038 22808
rect 20350 27512 20406 27568
rect 20258 24112 20314 24168
rect 20350 23976 20406 24032
rect 19430 21800 19486 21856
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 19982 20596 20038 20632
rect 19982 20576 19984 20596
rect 19984 20576 20036 20596
rect 20036 20576 20038 20596
rect 20166 22208 20222 22264
rect 20626 30368 20682 30424
rect 20626 29552 20682 29608
rect 20994 30232 21050 30288
rect 21794 31578 21850 31580
rect 21874 31578 21930 31580
rect 21954 31578 22010 31580
rect 22034 31578 22090 31580
rect 21794 31526 21840 31578
rect 21840 31526 21850 31578
rect 21874 31526 21904 31578
rect 21904 31526 21916 31578
rect 21916 31526 21930 31578
rect 21954 31526 21968 31578
rect 21968 31526 21980 31578
rect 21980 31526 22010 31578
rect 22034 31526 22044 31578
rect 22044 31526 22090 31578
rect 21794 31524 21850 31526
rect 21874 31524 21930 31526
rect 21954 31524 22010 31526
rect 22034 31524 22090 31526
rect 21730 31048 21786 31104
rect 21270 30504 21326 30560
rect 21086 29688 21142 29744
rect 20626 28872 20682 28928
rect 20994 29416 21050 29472
rect 20994 29008 21050 29064
rect 20718 28192 20774 28248
rect 20534 27784 20590 27840
rect 20718 27104 20774 27160
rect 20718 26696 20774 26752
rect 20718 26424 20774 26480
rect 20810 25900 20866 25936
rect 20810 25880 20812 25900
rect 20812 25880 20864 25900
rect 20864 25880 20866 25900
rect 20810 24928 20866 24984
rect 20718 24384 20774 24440
rect 20810 24248 20866 24304
rect 20626 23840 20682 23896
rect 20626 23432 20682 23488
rect 20534 23316 20590 23352
rect 20534 23296 20536 23316
rect 20536 23296 20588 23316
rect 20588 23296 20590 23316
rect 20534 21528 20590 21584
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 1582 20032 1638 20088
rect 20902 23840 20958 23896
rect 20810 23296 20866 23352
rect 20718 22752 20774 22808
rect 20810 21800 20866 21856
rect 21454 30504 21510 30560
rect 21794 30490 21850 30492
rect 21874 30490 21930 30492
rect 21954 30490 22010 30492
rect 22034 30490 22090 30492
rect 21794 30438 21840 30490
rect 21840 30438 21850 30490
rect 21874 30438 21904 30490
rect 21904 30438 21916 30490
rect 21916 30438 21930 30490
rect 21954 30438 21968 30490
rect 21968 30438 21980 30490
rect 21980 30438 22010 30490
rect 22034 30438 22044 30490
rect 22044 30438 22090 30490
rect 21794 30436 21850 30438
rect 21874 30436 21930 30438
rect 21954 30436 22010 30438
rect 22034 30436 22090 30438
rect 22558 30368 22614 30424
rect 21794 29402 21850 29404
rect 21874 29402 21930 29404
rect 21954 29402 22010 29404
rect 22034 29402 22090 29404
rect 21794 29350 21840 29402
rect 21840 29350 21850 29402
rect 21874 29350 21904 29402
rect 21904 29350 21916 29402
rect 21916 29350 21930 29402
rect 21954 29350 21968 29402
rect 21968 29350 21980 29402
rect 21980 29350 22010 29402
rect 22034 29350 22044 29402
rect 22044 29350 22090 29402
rect 21794 29348 21850 29350
rect 21874 29348 21930 29350
rect 21954 29348 22010 29350
rect 22034 29348 22090 29350
rect 22282 29008 22338 29064
rect 21362 27240 21418 27296
rect 21178 26560 21234 26616
rect 21178 26152 21234 26208
rect 21454 26832 21510 26888
rect 21546 26016 21602 26072
rect 21454 25880 21510 25936
rect 21362 25472 21418 25528
rect 21794 28314 21850 28316
rect 21874 28314 21930 28316
rect 21954 28314 22010 28316
rect 22034 28314 22090 28316
rect 21794 28262 21840 28314
rect 21840 28262 21850 28314
rect 21874 28262 21904 28314
rect 21904 28262 21916 28314
rect 21916 28262 21930 28314
rect 21954 28262 21968 28314
rect 21968 28262 21980 28314
rect 21980 28262 22010 28314
rect 22034 28262 22044 28314
rect 22044 28262 22090 28314
rect 21794 28260 21850 28262
rect 21874 28260 21930 28262
rect 21954 28260 22010 28262
rect 22034 28260 22090 28262
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 22006 26968 22062 27024
rect 21730 26852 21786 26888
rect 22282 27784 22338 27840
rect 21730 26832 21732 26852
rect 21732 26832 21784 26852
rect 21784 26832 21786 26852
rect 22098 26560 22154 26616
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 22098 25472 22154 25528
rect 21638 25064 21694 25120
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 21178 24384 21234 24440
rect 21270 23976 21326 24032
rect 21270 23704 21326 23760
rect 21638 23976 21694 24032
rect 21178 23568 21234 23624
rect 21546 23704 21602 23760
rect 21362 23432 21418 23488
rect 21270 22072 21326 22128
rect 20994 21936 21050 21992
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 22190 23840 22246 23896
rect 21178 21256 21234 21312
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 1582 19352 1638 19408
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 22006 23604 22008 23624
rect 22008 23604 22060 23624
rect 22060 23604 22062 23624
rect 22006 23568 22062 23604
rect 22098 23432 22154 23488
rect 21822 23044 21878 23080
rect 21822 23024 21824 23044
rect 21824 23024 21876 23044
rect 21876 23024 21878 23044
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 21822 22636 21878 22672
rect 21822 22616 21824 22636
rect 21824 22616 21876 22636
rect 21876 22616 21878 22636
rect 22558 27648 22614 27704
rect 22926 29588 22928 29608
rect 22928 29588 22980 29608
rect 22980 29588 22982 29608
rect 22926 29552 22982 29588
rect 22926 29416 22982 29472
rect 22834 28736 22890 28792
rect 22742 27784 22798 27840
rect 22558 27104 22614 27160
rect 22558 26968 22614 27024
rect 22466 25472 22522 25528
rect 22190 22616 22246 22672
rect 22282 22380 22284 22400
rect 22284 22380 22336 22400
rect 22336 22380 22338 22400
rect 22282 22344 22338 22380
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 22466 22772 22522 22808
rect 22466 22752 22468 22772
rect 22468 22752 22520 22772
rect 22520 22752 22522 22772
rect 22466 22072 22522 22128
rect 22466 21564 22468 21584
rect 22468 21564 22520 21584
rect 22520 21564 22522 21584
rect 22466 21528 22522 21564
rect 23110 28872 23166 28928
rect 23018 28328 23074 28384
rect 23110 27648 23166 27704
rect 23110 27512 23166 27568
rect 22834 25064 22890 25120
rect 22834 24384 22890 24440
rect 23110 27104 23166 27160
rect 23570 28872 23626 28928
rect 23294 27784 23350 27840
rect 23662 28600 23718 28656
rect 23754 28328 23810 28384
rect 23386 26832 23442 26888
rect 23294 26560 23350 26616
rect 23110 26188 23112 26208
rect 23112 26188 23164 26208
rect 23164 26188 23166 26208
rect 23110 26152 23166 26188
rect 23386 26016 23442 26072
rect 23294 24928 23350 24984
rect 22834 24112 22890 24168
rect 23202 24112 23258 24168
rect 22834 23976 22890 24032
rect 23018 22888 23074 22944
rect 22650 21292 22652 21312
rect 22652 21292 22704 21312
rect 22704 21292 22706 21312
rect 22650 21256 22706 21292
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 1582 18028 1584 18048
rect 1584 18028 1636 18048
rect 1636 18028 1638 18048
rect 1582 17992 1638 18028
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 1582 17312 1638 17368
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 23018 22072 23074 22128
rect 23018 21956 23074 21992
rect 23018 21936 23020 21956
rect 23020 21936 23072 21956
rect 23072 21936 23074 21956
rect 23846 27820 23848 27840
rect 23848 27820 23900 27840
rect 23900 27820 23902 27840
rect 23846 27784 23902 27820
rect 23754 27512 23810 27568
rect 23662 26424 23718 26480
rect 23386 23296 23442 23352
rect 23294 22752 23350 22808
rect 23386 22480 23442 22536
rect 23570 22636 23626 22672
rect 23570 22616 23572 22636
rect 23572 22616 23624 22636
rect 23624 22616 23626 22636
rect 23202 22208 23258 22264
rect 23386 21936 23442 21992
rect 23294 21664 23350 21720
rect 23938 23432 23994 23488
rect 23938 22752 23994 22808
rect 24398 29280 24454 29336
rect 24582 30232 24638 30288
rect 24398 26968 24454 27024
rect 24122 24384 24178 24440
rect 24398 23568 24454 23624
rect 24306 23296 24362 23352
rect 23754 21256 23810 21312
rect 24582 26016 24638 26072
rect 24582 24556 24584 24576
rect 24584 24556 24636 24576
rect 24636 24556 24638 24576
rect 24582 24520 24638 24556
rect 25267 31034 25323 31036
rect 25347 31034 25403 31036
rect 25427 31034 25483 31036
rect 25507 31034 25563 31036
rect 25267 30982 25313 31034
rect 25313 30982 25323 31034
rect 25347 30982 25377 31034
rect 25377 30982 25389 31034
rect 25389 30982 25403 31034
rect 25427 30982 25441 31034
rect 25441 30982 25453 31034
rect 25453 30982 25483 31034
rect 25507 30982 25517 31034
rect 25517 30982 25563 31034
rect 25267 30980 25323 30982
rect 25347 30980 25403 30982
rect 25427 30980 25483 30982
rect 25507 30980 25563 30982
rect 25226 30232 25282 30288
rect 25134 30096 25190 30152
rect 25042 29996 25044 30016
rect 25044 29996 25096 30016
rect 25096 29996 25098 30016
rect 25042 29960 25098 29996
rect 25267 29946 25323 29948
rect 25347 29946 25403 29948
rect 25427 29946 25483 29948
rect 25507 29946 25563 29948
rect 25267 29894 25313 29946
rect 25313 29894 25323 29946
rect 25347 29894 25377 29946
rect 25377 29894 25389 29946
rect 25389 29894 25403 29946
rect 25427 29894 25441 29946
rect 25441 29894 25453 29946
rect 25453 29894 25483 29946
rect 25507 29894 25517 29946
rect 25517 29894 25563 29946
rect 25267 29892 25323 29894
rect 25347 29892 25403 29894
rect 25427 29892 25483 29894
rect 25507 29892 25563 29894
rect 24950 28872 25006 28928
rect 25042 27648 25098 27704
rect 25267 28858 25323 28860
rect 25347 28858 25403 28860
rect 25427 28858 25483 28860
rect 25507 28858 25563 28860
rect 25267 28806 25313 28858
rect 25313 28806 25323 28858
rect 25347 28806 25377 28858
rect 25377 28806 25389 28858
rect 25389 28806 25403 28858
rect 25427 28806 25441 28858
rect 25441 28806 25453 28858
rect 25453 28806 25483 28858
rect 25507 28806 25517 28858
rect 25517 28806 25563 28858
rect 25267 28804 25323 28806
rect 25347 28804 25403 28806
rect 25427 28804 25483 28806
rect 25507 28804 25563 28806
rect 25410 28500 25412 28520
rect 25412 28500 25464 28520
rect 25464 28500 25466 28520
rect 25410 28464 25466 28500
rect 25318 27920 25374 27976
rect 25502 27956 25504 27976
rect 25504 27956 25556 27976
rect 25556 27956 25558 27976
rect 25502 27920 25558 27956
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 25502 27104 25558 27160
rect 25226 26868 25228 26888
rect 25228 26868 25280 26888
rect 25280 26868 25282 26888
rect 25226 26832 25282 26868
rect 25686 27512 25742 27568
rect 25962 29280 26018 29336
rect 25870 27376 25926 27432
rect 25778 26832 25834 26888
rect 24950 26696 25006 26752
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 25686 26560 25742 26616
rect 26422 31184 26478 31240
rect 26422 30368 26478 30424
rect 25962 26560 26018 26616
rect 24858 25492 24914 25528
rect 24858 25472 24860 25492
rect 24860 25472 24912 25492
rect 24912 25472 24914 25492
rect 24950 25336 25006 25392
rect 24950 24656 25006 24712
rect 25134 26152 25190 26208
rect 25318 26152 25374 26208
rect 25226 26016 25282 26072
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25134 25472 25190 25528
rect 25226 25336 25282 25392
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25870 25472 25926 25528
rect 26146 26424 26202 26480
rect 25870 24928 25926 24984
rect 25778 24656 25834 24712
rect 25778 24384 25834 24440
rect 25134 24248 25190 24304
rect 25410 24248 25466 24304
rect 25134 23976 25190 24032
rect 25594 23840 25650 23896
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25410 22752 25466 22808
rect 25778 22772 25834 22808
rect 25778 22752 25780 22772
rect 25780 22752 25832 22772
rect 25832 22752 25834 22772
rect 25870 22616 25926 22672
rect 24674 22344 24730 22400
rect 24858 21392 24914 21448
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25870 22228 25926 22264
rect 25870 22208 25872 22228
rect 25872 22208 25924 22228
rect 25924 22208 25926 22228
rect 25594 20304 25650 20360
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 26422 26288 26478 26344
rect 26330 24928 26386 24984
rect 26698 27784 26754 27840
rect 26606 26852 26662 26888
rect 26606 26832 26608 26852
rect 26608 26832 26660 26852
rect 26660 26832 26662 26852
rect 26514 25880 26570 25936
rect 26606 25220 26662 25256
rect 26606 25200 26608 25220
rect 26608 25200 26660 25220
rect 26660 25200 26662 25220
rect 26238 23840 26294 23896
rect 26238 22888 26294 22944
rect 28170 31320 28226 31376
rect 27158 30776 27214 30832
rect 27342 28192 27398 28248
rect 27618 29008 27674 29064
rect 27526 28600 27582 28656
rect 27434 28056 27490 28112
rect 27158 26968 27214 27024
rect 27158 25764 27214 25800
rect 27158 25744 27160 25764
rect 27160 25744 27212 25764
rect 27212 25744 27214 25764
rect 27342 24928 27398 24984
rect 26882 23568 26938 23624
rect 27250 24248 27306 24304
rect 27158 24112 27214 24168
rect 27158 23976 27214 24032
rect 27066 23160 27122 23216
rect 26974 23024 27030 23080
rect 27618 26832 27674 26888
rect 27802 29164 27858 29200
rect 27802 29144 27804 29164
rect 27804 29144 27856 29164
rect 27856 29144 27858 29164
rect 27802 27920 27858 27976
rect 27710 26152 27766 26208
rect 27526 26016 27582 26072
rect 28170 28464 28226 28520
rect 28262 27240 28318 27296
rect 27894 25744 27950 25800
rect 27802 25336 27858 25392
rect 27526 25064 27582 25120
rect 27526 24248 27582 24304
rect 27710 24792 27766 24848
rect 27710 22072 27766 22128
rect 28170 24384 28226 24440
rect 28354 23724 28410 23760
rect 28354 23704 28356 23724
rect 28356 23704 28408 23724
rect 28408 23704 28410 23724
rect 28354 23060 28356 23080
rect 28356 23060 28408 23080
rect 28408 23060 28410 23080
rect 28354 23024 28410 23060
rect 28262 22344 28318 22400
rect 28354 21528 28410 21584
rect 28740 31578 28796 31580
rect 28820 31578 28876 31580
rect 28900 31578 28956 31580
rect 28980 31578 29036 31580
rect 28740 31526 28786 31578
rect 28786 31526 28796 31578
rect 28820 31526 28850 31578
rect 28850 31526 28862 31578
rect 28862 31526 28876 31578
rect 28900 31526 28914 31578
rect 28914 31526 28926 31578
rect 28926 31526 28956 31578
rect 28980 31526 28990 31578
rect 28990 31526 29036 31578
rect 28740 31524 28796 31526
rect 28820 31524 28876 31526
rect 28900 31524 28956 31526
rect 28980 31524 29036 31526
rect 28998 31184 29054 31240
rect 28740 30490 28796 30492
rect 28820 30490 28876 30492
rect 28900 30490 28956 30492
rect 28980 30490 29036 30492
rect 28740 30438 28786 30490
rect 28786 30438 28796 30490
rect 28820 30438 28850 30490
rect 28850 30438 28862 30490
rect 28862 30438 28876 30490
rect 28900 30438 28914 30490
rect 28914 30438 28926 30490
rect 28926 30438 28956 30490
rect 28980 30438 28990 30490
rect 28990 30438 29036 30490
rect 28740 30436 28796 30438
rect 28820 30436 28876 30438
rect 28900 30436 28956 30438
rect 28980 30436 29036 30438
rect 28538 29824 28594 29880
rect 28740 29402 28796 29404
rect 28820 29402 28876 29404
rect 28900 29402 28956 29404
rect 28980 29402 29036 29404
rect 28740 29350 28786 29402
rect 28786 29350 28796 29402
rect 28820 29350 28850 29402
rect 28850 29350 28862 29402
rect 28862 29350 28876 29402
rect 28900 29350 28914 29402
rect 28914 29350 28926 29402
rect 28926 29350 28956 29402
rect 28980 29350 28990 29402
rect 28990 29350 29036 29402
rect 28740 29348 28796 29350
rect 28820 29348 28876 29350
rect 28900 29348 28956 29350
rect 28980 29348 29036 29350
rect 28998 29144 29054 29200
rect 28740 28314 28796 28316
rect 28820 28314 28876 28316
rect 28900 28314 28956 28316
rect 28980 28314 29036 28316
rect 28740 28262 28786 28314
rect 28786 28262 28796 28314
rect 28820 28262 28850 28314
rect 28850 28262 28862 28314
rect 28862 28262 28876 28314
rect 28900 28262 28914 28314
rect 28914 28262 28926 28314
rect 28926 28262 28956 28314
rect 28980 28262 28990 28314
rect 28990 28262 29036 28314
rect 28740 28260 28796 28262
rect 28820 28260 28876 28262
rect 28900 28260 28956 28262
rect 28980 28260 29036 28262
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 28630 26968 28686 27024
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28354 20984 28410 21040
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28354 20304 28410 20360
rect 28354 19796 28356 19816
rect 28356 19796 28408 19816
rect 28408 19796 28410 19816
rect 28354 19760 28410 19796
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28354 18944 28410 19000
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28354 18300 28356 18320
rect 28356 18300 28408 18320
rect 28408 18300 28410 18320
rect 28354 18264 28410 18300
rect 28354 17620 28356 17640
rect 28356 17620 28408 17640
rect 28408 17620 28410 17640
rect 28354 17584 28410 17620
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28354 16940 28356 16960
rect 28356 16940 28408 16960
rect 28408 16940 28410 16960
rect 28354 16904 28410 16940
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 1582 15988 1584 16008
rect 1584 15988 1636 16008
rect 1636 15988 1638 16008
rect 1582 15952 1638 15988
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 28354 15544 28410 15600
rect 1582 15272 1638 15328
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 28354 14884 28410 14920
rect 28354 14864 28356 14884
rect 28356 14864 28408 14884
rect 28408 14864 28410 14884
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 1582 13912 1638 13968
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 28354 13504 28410 13560
rect 1582 13268 1584 13288
rect 1584 13268 1636 13288
rect 1636 13268 1638 13288
rect 1582 13232 1638 13268
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28354 12824 28410 12880
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 1582 11872 1638 11928
rect 28354 11500 28356 11520
rect 28356 11500 28408 11520
rect 28408 11500 28410 11520
rect 28354 11464 28410 11500
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 1582 11192 1638 11248
rect 28354 11092 28356 11112
rect 28356 11092 28408 11112
rect 28408 11092 28410 11112
rect 28354 11056 28410 11092
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 1582 9832 1638 9888
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28354 9444 28410 9480
rect 28354 9424 28356 9444
rect 28356 9424 28408 9444
rect 28408 9424 28410 9444
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 1582 9152 1638 9208
rect 28354 9052 28356 9072
rect 28356 9052 28408 9072
rect 28408 9052 28410 9072
rect 28354 9016 28410 9052
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 1582 7828 1584 7848
rect 1584 7828 1636 7848
rect 1636 7828 1638 7848
rect 1582 7792 1638 7828
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28354 7384 28410 7440
rect 1582 7148 1584 7168
rect 1584 7148 1636 7168
rect 1636 7148 1638 7168
rect 1582 7112 1638 7148
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 28354 6740 28356 6760
rect 28356 6740 28408 6760
rect 28408 6740 28410 6760
rect 28354 6704 28410 6740
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 1582 5752 1638 5808
rect 28354 5652 28356 5672
rect 28356 5652 28408 5672
rect 28408 5652 28410 5672
rect 28354 5616 28410 5652
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 1582 5108 1584 5128
rect 1584 5108 1636 5128
rect 1636 5108 1638 5128
rect 1582 5072 1638 5108
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 28354 4664 28410 4720
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 1582 3712 1638 3768
rect 28354 3612 28356 3632
rect 28356 3612 28408 3632
rect 28408 3612 28410 3632
rect 28354 3576 28410 3612
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 1582 3032 1638 3088
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 28354 2624 28410 2680
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
<< metal3 >>
rect 25998 31860 26004 31924
rect 26068 31922 26074 31924
rect 29200 31922 30000 31952
rect 26068 31862 30000 31922
rect 26068 31860 26074 31862
rect 29200 31832 30000 31862
rect 13537 31786 13603 31789
rect 23238 31786 23244 31788
rect 13537 31784 23244 31786
rect 13537 31728 13542 31784
rect 13598 31728 23244 31784
rect 13537 31726 23244 31728
rect 13537 31723 13603 31726
rect 23238 31724 23244 31726
rect 23308 31724 23314 31788
rect 17125 31650 17191 31653
rect 18229 31650 18295 31653
rect 17125 31648 18295 31650
rect 17125 31592 17130 31648
rect 17186 31592 18234 31648
rect 18290 31592 18295 31648
rect 17125 31590 18295 31592
rect 17125 31587 17191 31590
rect 18229 31587 18295 31590
rect 7892 31584 8208 31585
rect 7892 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8208 31584
rect 7892 31519 8208 31520
rect 14838 31584 15154 31585
rect 14838 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15154 31584
rect 14838 31519 15154 31520
rect 21784 31584 22100 31585
rect 21784 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22100 31584
rect 21784 31519 22100 31520
rect 28730 31584 29046 31585
rect 28730 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29046 31584
rect 28730 31519 29046 31520
rect 15653 31514 15719 31517
rect 21214 31514 21220 31516
rect 15653 31512 21220 31514
rect 15653 31456 15658 31512
rect 15714 31456 21220 31512
rect 15653 31454 21220 31456
rect 15653 31451 15719 31454
rect 21214 31452 21220 31454
rect 21284 31452 21290 31516
rect 11145 31378 11211 31381
rect 28165 31378 28231 31381
rect 11145 31376 28231 31378
rect 11145 31320 11150 31376
rect 11206 31320 28170 31376
rect 28226 31320 28231 31376
rect 11145 31318 28231 31320
rect 11145 31315 11211 31318
rect 28165 31315 28231 31318
rect 11973 31242 12039 31245
rect 26417 31242 26483 31245
rect 11973 31240 26483 31242
rect 11973 31184 11978 31240
rect 12034 31184 26422 31240
rect 26478 31184 26483 31240
rect 11973 31182 26483 31184
rect 11973 31179 12039 31182
rect 26417 31179 26483 31182
rect 28993 31242 29059 31245
rect 29200 31242 30000 31272
rect 28993 31240 30000 31242
rect 28993 31184 28998 31240
rect 29054 31184 30000 31240
rect 28993 31182 30000 31184
rect 28993 31179 29059 31182
rect 29200 31152 30000 31182
rect 11973 31106 12039 31109
rect 13353 31106 13419 31109
rect 11973 31104 13419 31106
rect 11973 31048 11978 31104
rect 12034 31048 13358 31104
rect 13414 31048 13419 31104
rect 11973 31046 13419 31048
rect 11973 31043 12039 31046
rect 13353 31043 13419 31046
rect 18822 31044 18828 31108
rect 18892 31106 18898 31108
rect 21725 31106 21791 31109
rect 18892 31104 21791 31106
rect 18892 31048 21730 31104
rect 21786 31048 21791 31104
rect 18892 31046 21791 31048
rect 18892 31044 18898 31046
rect 21725 31043 21791 31046
rect 4419 31040 4735 31041
rect 0 30880 800 31000
rect 4419 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4735 31040
rect 4419 30975 4735 30976
rect 11365 31040 11681 31041
rect 11365 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11681 31040
rect 11365 30975 11681 30976
rect 18311 31040 18627 31041
rect 18311 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18627 31040
rect 18311 30975 18627 30976
rect 25257 31040 25573 31041
rect 25257 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25573 31040
rect 25257 30975 25573 30976
rect 12065 30970 12131 30973
rect 17953 30970 18019 30973
rect 12065 30968 18019 30970
rect 12065 30912 12070 30968
rect 12126 30912 17958 30968
rect 18014 30912 18019 30968
rect 12065 30910 18019 30912
rect 12065 30907 12131 30910
rect 17953 30907 18019 30910
rect 18689 30970 18755 30973
rect 23422 30970 23428 30972
rect 18689 30968 23428 30970
rect 18689 30912 18694 30968
rect 18750 30912 23428 30968
rect 18689 30910 23428 30912
rect 18689 30907 18755 30910
rect 23422 30908 23428 30910
rect 23492 30908 23498 30972
rect 9305 30834 9371 30837
rect 27153 30834 27219 30837
rect 9305 30832 27219 30834
rect 9305 30776 9310 30832
rect 9366 30776 27158 30832
rect 27214 30776 27219 30832
rect 9305 30774 27219 30776
rect 9305 30771 9371 30774
rect 27153 30771 27219 30774
rect 5349 30698 5415 30701
rect 5349 30696 15946 30698
rect 5349 30640 5354 30696
rect 5410 30640 15946 30696
rect 5349 30638 15946 30640
rect 5349 30635 5415 30638
rect 15886 30562 15946 30638
rect 17350 30636 17356 30700
rect 17420 30698 17426 30700
rect 17493 30698 17559 30701
rect 17420 30696 17559 30698
rect 17420 30640 17498 30696
rect 17554 30640 17559 30696
rect 17420 30638 17559 30640
rect 17420 30636 17426 30638
rect 17493 30635 17559 30638
rect 17677 30698 17743 30701
rect 17902 30698 17908 30700
rect 17677 30696 17908 30698
rect 17677 30640 17682 30696
rect 17738 30640 17908 30696
rect 17677 30638 17908 30640
rect 17677 30635 17743 30638
rect 17902 30636 17908 30638
rect 17972 30636 17978 30700
rect 18137 30698 18203 30701
rect 23054 30698 23060 30700
rect 18137 30696 23060 30698
rect 18137 30640 18142 30696
rect 18198 30640 23060 30696
rect 18137 30638 23060 30640
rect 18137 30635 18203 30638
rect 23054 30636 23060 30638
rect 23124 30636 23130 30700
rect 19425 30562 19491 30565
rect 15886 30560 19491 30562
rect 15886 30504 19430 30560
rect 19486 30504 19491 30560
rect 15886 30502 19491 30504
rect 19425 30499 19491 30502
rect 19609 30562 19675 30565
rect 19926 30562 19932 30564
rect 19609 30560 19932 30562
rect 19609 30504 19614 30560
rect 19670 30504 19932 30560
rect 19609 30502 19932 30504
rect 19609 30499 19675 30502
rect 19926 30500 19932 30502
rect 19996 30500 20002 30564
rect 21265 30562 21331 30565
rect 21449 30562 21515 30565
rect 21265 30560 21515 30562
rect 21265 30504 21270 30560
rect 21326 30504 21454 30560
rect 21510 30504 21515 30560
rect 21265 30502 21515 30504
rect 21265 30499 21331 30502
rect 21449 30499 21515 30502
rect 7892 30496 8208 30497
rect 7892 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8208 30496
rect 7892 30431 8208 30432
rect 14838 30496 15154 30497
rect 14838 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15154 30496
rect 14838 30431 15154 30432
rect 21784 30496 22100 30497
rect 21784 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22100 30496
rect 21784 30431 22100 30432
rect 28730 30496 29046 30497
rect 28730 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29046 30496
rect 29200 30472 30000 30592
rect 28730 30431 29046 30432
rect 10041 30426 10107 30429
rect 9446 30424 10107 30426
rect 9446 30368 10046 30424
rect 10102 30368 10107 30424
rect 9446 30366 10107 30368
rect 0 30290 800 30320
rect 1577 30290 1643 30293
rect 0 30288 1643 30290
rect 0 30232 1582 30288
rect 1638 30232 1643 30288
rect 0 30230 1643 30232
rect 0 30200 800 30230
rect 1577 30227 1643 30230
rect 6545 30290 6611 30293
rect 9446 30290 9506 30366
rect 10041 30363 10107 30366
rect 11789 30426 11855 30429
rect 12014 30426 12020 30428
rect 11789 30424 12020 30426
rect 11789 30368 11794 30424
rect 11850 30368 12020 30424
rect 11789 30366 12020 30368
rect 11789 30363 11855 30366
rect 12014 30364 12020 30366
rect 12084 30364 12090 30428
rect 17585 30426 17651 30429
rect 19057 30426 19123 30429
rect 17585 30424 19123 30426
rect 17585 30368 17590 30424
rect 17646 30368 19062 30424
rect 19118 30368 19123 30424
rect 17585 30366 19123 30368
rect 17585 30363 17651 30366
rect 19057 30363 19123 30366
rect 19517 30426 19583 30429
rect 20478 30426 20484 30428
rect 19517 30424 20484 30426
rect 19517 30368 19522 30424
rect 19578 30368 20484 30424
rect 19517 30366 20484 30368
rect 19517 30363 19583 30366
rect 20478 30364 20484 30366
rect 20548 30364 20554 30428
rect 20621 30426 20687 30429
rect 22553 30426 22619 30429
rect 26417 30426 26483 30429
rect 20621 30424 21466 30426
rect 20621 30368 20626 30424
rect 20682 30368 21466 30424
rect 20621 30366 21466 30368
rect 20621 30363 20687 30366
rect 6545 30288 9506 30290
rect 6545 30232 6550 30288
rect 6606 30232 9506 30288
rect 6545 30230 9506 30232
rect 9581 30290 9647 30293
rect 14181 30290 14247 30293
rect 9581 30288 14247 30290
rect 9581 30232 9586 30288
rect 9642 30232 14186 30288
rect 14242 30232 14247 30288
rect 9581 30230 14247 30232
rect 6545 30227 6611 30230
rect 9581 30227 9647 30230
rect 14181 30227 14247 30230
rect 15285 30292 15351 30293
rect 15285 30288 15332 30292
rect 15396 30290 15402 30292
rect 17125 30290 17191 30293
rect 20989 30290 21055 30293
rect 15285 30232 15290 30288
rect 15285 30228 15332 30232
rect 15396 30230 15442 30290
rect 17125 30288 21055 30290
rect 17125 30232 17130 30288
rect 17186 30232 20994 30288
rect 21050 30232 21055 30288
rect 17125 30230 21055 30232
rect 21406 30290 21466 30366
rect 22553 30424 26483 30426
rect 22553 30368 22558 30424
rect 22614 30368 26422 30424
rect 26478 30368 26483 30424
rect 22553 30366 26483 30368
rect 22553 30363 22619 30366
rect 26417 30363 26483 30366
rect 24577 30290 24643 30293
rect 25221 30290 25287 30293
rect 21406 30288 25287 30290
rect 21406 30232 24582 30288
rect 24638 30232 25226 30288
rect 25282 30232 25287 30288
rect 21406 30230 25287 30232
rect 15396 30228 15402 30230
rect 15285 30227 15351 30228
rect 17125 30227 17191 30230
rect 20989 30227 21055 30230
rect 24577 30227 24643 30230
rect 25221 30227 25287 30230
rect 9765 30154 9831 30157
rect 9990 30154 9996 30156
rect 9765 30152 9996 30154
rect 9765 30096 9770 30152
rect 9826 30096 9996 30152
rect 9765 30094 9996 30096
rect 9765 30091 9831 30094
rect 9990 30092 9996 30094
rect 10060 30092 10066 30156
rect 11145 30154 11211 30157
rect 19149 30156 19215 30157
rect 19149 30154 19196 30156
rect 11145 30152 18890 30154
rect 11145 30096 11150 30152
rect 11206 30096 18890 30152
rect 11145 30094 18890 30096
rect 19104 30152 19196 30154
rect 19104 30096 19154 30152
rect 19104 30094 19196 30096
rect 11145 30091 11211 30094
rect 13261 30018 13327 30021
rect 15009 30018 15075 30021
rect 13261 30016 15075 30018
rect 13261 29960 13266 30016
rect 13322 29960 15014 30016
rect 15070 29960 15075 30016
rect 13261 29958 15075 29960
rect 13261 29955 13327 29958
rect 15009 29955 15075 29958
rect 16798 29956 16804 30020
rect 16868 30018 16874 30020
rect 17953 30018 18019 30021
rect 16868 30016 18019 30018
rect 16868 29960 17958 30016
rect 18014 29960 18019 30016
rect 16868 29958 18019 29960
rect 18830 30018 18890 30094
rect 19149 30092 19196 30094
rect 19260 30092 19266 30156
rect 19425 30154 19491 30157
rect 25129 30154 25195 30157
rect 19425 30152 25195 30154
rect 19425 30096 19430 30152
rect 19486 30096 25134 30152
rect 25190 30096 25195 30152
rect 19425 30094 25195 30096
rect 19149 30091 19215 30092
rect 19425 30091 19491 30094
rect 25129 30091 25195 30094
rect 25037 30020 25103 30021
rect 20662 30018 20668 30020
rect 18830 29958 20668 30018
rect 16868 29956 16874 29958
rect 17953 29955 18019 29958
rect 20662 29956 20668 29958
rect 20732 29956 20738 30020
rect 25037 30018 25084 30020
rect 23430 30016 25084 30018
rect 23430 29960 25042 30016
rect 23430 29958 25084 29960
rect 4419 29952 4735 29953
rect 4419 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4735 29952
rect 4419 29887 4735 29888
rect 11365 29952 11681 29953
rect 11365 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11681 29952
rect 11365 29887 11681 29888
rect 18311 29952 18627 29953
rect 18311 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18627 29952
rect 18311 29887 18627 29888
rect 14181 29882 14247 29885
rect 16205 29882 16271 29885
rect 17125 29882 17191 29885
rect 17309 29882 17375 29885
rect 14181 29880 17375 29882
rect 14181 29824 14186 29880
rect 14242 29824 16210 29880
rect 16266 29824 17130 29880
rect 17186 29824 17314 29880
rect 17370 29824 17375 29880
rect 14181 29822 17375 29824
rect 14181 29819 14247 29822
rect 16205 29819 16271 29822
rect 17125 29819 17191 29822
rect 17309 29819 17375 29822
rect 18045 29884 18111 29885
rect 18045 29880 18092 29884
rect 18156 29882 18162 29884
rect 19333 29882 19399 29885
rect 19793 29882 19859 29885
rect 23430 29882 23490 29958
rect 25037 29956 25084 29958
rect 25148 29956 25154 30020
rect 25037 29955 25103 29956
rect 25257 29952 25573 29953
rect 25257 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25573 29952
rect 25257 29887 25573 29888
rect 18045 29824 18050 29880
rect 18045 29820 18092 29824
rect 18156 29822 18202 29882
rect 19333 29880 23490 29882
rect 19333 29824 19338 29880
rect 19394 29824 19798 29880
rect 19854 29824 23490 29880
rect 19333 29822 23490 29824
rect 28533 29882 28599 29885
rect 29200 29882 30000 29912
rect 28533 29880 30000 29882
rect 28533 29824 28538 29880
rect 28594 29824 30000 29880
rect 28533 29822 30000 29824
rect 18156 29820 18162 29822
rect 18045 29819 18111 29820
rect 19333 29819 19399 29822
rect 19793 29819 19859 29822
rect 28533 29819 28599 29822
rect 29200 29792 30000 29822
rect 9765 29746 9831 29749
rect 11329 29746 11395 29749
rect 20846 29746 20852 29748
rect 9765 29744 11208 29746
rect 9765 29688 9770 29744
rect 9826 29688 11208 29744
rect 9765 29686 11208 29688
rect 9765 29683 9831 29686
rect 0 29610 800 29640
rect 1577 29610 1643 29613
rect 0 29608 1643 29610
rect 0 29552 1582 29608
rect 1638 29552 1643 29608
rect 0 29550 1643 29552
rect 11148 29610 11208 29686
rect 11329 29744 20852 29746
rect 11329 29688 11334 29744
rect 11390 29688 20852 29744
rect 11329 29686 20852 29688
rect 11329 29683 11395 29686
rect 20846 29684 20852 29686
rect 20916 29684 20922 29748
rect 21081 29746 21147 29749
rect 21081 29744 23122 29746
rect 21081 29688 21086 29744
rect 21142 29688 23122 29744
rect 21081 29686 23122 29688
rect 21081 29683 21147 29686
rect 13261 29610 13327 29613
rect 11148 29608 13327 29610
rect 11148 29552 13266 29608
rect 13322 29552 13327 29608
rect 11148 29550 13327 29552
rect 0 29520 800 29550
rect 1577 29547 1643 29550
rect 13261 29547 13327 29550
rect 13721 29610 13787 29613
rect 19374 29610 19380 29612
rect 13721 29608 19380 29610
rect 13721 29552 13726 29608
rect 13782 29552 19380 29608
rect 13721 29550 19380 29552
rect 13721 29547 13787 29550
rect 19374 29548 19380 29550
rect 19444 29548 19450 29612
rect 20621 29610 20687 29613
rect 22921 29610 22987 29613
rect 20621 29608 22987 29610
rect 20621 29552 20626 29608
rect 20682 29552 22926 29608
rect 22982 29552 22987 29608
rect 20621 29550 22987 29552
rect 20621 29547 20687 29550
rect 22921 29547 22987 29550
rect 12893 29474 12959 29477
rect 14089 29474 14155 29477
rect 12893 29472 14155 29474
rect 12893 29416 12898 29472
rect 12954 29416 14094 29472
rect 14150 29416 14155 29472
rect 12893 29414 14155 29416
rect 12893 29411 12959 29414
rect 14089 29411 14155 29414
rect 15745 29474 15811 29477
rect 15878 29474 15884 29476
rect 15745 29472 15884 29474
rect 15745 29416 15750 29472
rect 15806 29416 15884 29472
rect 15745 29414 15884 29416
rect 15745 29411 15811 29414
rect 15878 29412 15884 29414
rect 15948 29474 15954 29476
rect 17861 29474 17927 29477
rect 15948 29472 17927 29474
rect 15948 29416 17866 29472
rect 17922 29416 17927 29472
rect 15948 29414 17927 29416
rect 15948 29412 15954 29414
rect 17861 29411 17927 29414
rect 18086 29412 18092 29476
rect 18156 29474 18162 29476
rect 18689 29474 18755 29477
rect 20989 29474 21055 29477
rect 18156 29472 21055 29474
rect 18156 29416 18694 29472
rect 18750 29416 20994 29472
rect 21050 29416 21055 29472
rect 18156 29414 21055 29416
rect 18156 29412 18162 29414
rect 18689 29411 18755 29414
rect 20989 29411 21055 29414
rect 22921 29474 22987 29477
rect 23062 29474 23122 29686
rect 22921 29472 23122 29474
rect 22921 29416 22926 29472
rect 22982 29416 23122 29472
rect 22921 29414 23122 29416
rect 22921 29411 22987 29414
rect 7892 29408 8208 29409
rect 7892 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8208 29408
rect 7892 29343 8208 29344
rect 14838 29408 15154 29409
rect 14838 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15154 29408
rect 14838 29343 15154 29344
rect 21784 29408 22100 29409
rect 21784 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22100 29408
rect 21784 29343 22100 29344
rect 28730 29408 29046 29409
rect 28730 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29046 29408
rect 28730 29343 29046 29344
rect 8477 29338 8543 29341
rect 13353 29338 13419 29341
rect 8477 29336 13419 29338
rect 8477 29280 8482 29336
rect 8538 29280 13358 29336
rect 13414 29280 13419 29336
rect 8477 29278 13419 29280
rect 8477 29275 8543 29278
rect 13353 29275 13419 29278
rect 15745 29338 15811 29341
rect 16614 29338 16620 29340
rect 15745 29336 16620 29338
rect 15745 29280 15750 29336
rect 15806 29280 16620 29336
rect 15745 29278 16620 29280
rect 15745 29275 15811 29278
rect 16614 29276 16620 29278
rect 16684 29276 16690 29340
rect 16757 29338 16823 29341
rect 17718 29338 17724 29340
rect 16757 29336 17724 29338
rect 16757 29280 16762 29336
rect 16818 29280 17724 29336
rect 16757 29278 17724 29280
rect 16757 29275 16823 29278
rect 17718 29276 17724 29278
rect 17788 29276 17794 29340
rect 17953 29338 18019 29341
rect 18321 29338 18387 29341
rect 17953 29336 18387 29338
rect 17953 29280 17958 29336
rect 18014 29280 18326 29336
rect 18382 29280 18387 29336
rect 17953 29278 18387 29280
rect 17953 29275 18019 29278
rect 18321 29275 18387 29278
rect 18505 29338 18571 29341
rect 18822 29338 18828 29340
rect 18505 29336 18828 29338
rect 18505 29280 18510 29336
rect 18566 29280 18828 29336
rect 18505 29278 18828 29280
rect 18505 29275 18571 29278
rect 18822 29276 18828 29278
rect 18892 29276 18898 29340
rect 24393 29338 24459 29341
rect 25957 29338 26023 29341
rect 24393 29336 26023 29338
rect 24393 29280 24398 29336
rect 24454 29280 25962 29336
rect 26018 29280 26023 29336
rect 24393 29278 26023 29280
rect 24393 29275 24459 29278
rect 25957 29275 26023 29278
rect 11697 29202 11763 29205
rect 17861 29202 17927 29205
rect 27797 29202 27863 29205
rect 11697 29200 17740 29202
rect 11697 29144 11702 29200
rect 11758 29144 17740 29200
rect 11697 29142 17740 29144
rect 11697 29139 11763 29142
rect 9673 29066 9739 29069
rect 9990 29066 9996 29068
rect 9673 29064 9996 29066
rect 9673 29008 9678 29064
rect 9734 29008 9996 29064
rect 9673 29006 9996 29008
rect 9673 29003 9739 29006
rect 9990 29004 9996 29006
rect 10060 29004 10066 29068
rect 10593 29066 10659 29069
rect 10910 29066 10916 29068
rect 10593 29064 10916 29066
rect 10593 29008 10598 29064
rect 10654 29008 10916 29064
rect 10593 29006 10916 29008
rect 10593 29003 10659 29006
rect 10910 29004 10916 29006
rect 10980 29004 10986 29068
rect 11881 29066 11947 29069
rect 12198 29066 12204 29068
rect 11881 29064 12204 29066
rect 11881 29008 11886 29064
rect 11942 29008 12204 29064
rect 11881 29006 12204 29008
rect 11881 29003 11947 29006
rect 12198 29004 12204 29006
rect 12268 29004 12274 29068
rect 14457 29066 14523 29069
rect 14590 29066 14596 29068
rect 14457 29064 14596 29066
rect 14457 29008 14462 29064
rect 14518 29008 14596 29064
rect 14457 29006 14596 29008
rect 14457 29003 14523 29006
rect 14590 29004 14596 29006
rect 14660 29004 14666 29068
rect 17033 29066 17099 29069
rect 17401 29068 17467 29069
rect 17166 29066 17172 29068
rect 17033 29064 17172 29066
rect 17033 29008 17038 29064
rect 17094 29008 17172 29064
rect 17033 29006 17172 29008
rect 17033 29003 17099 29006
rect 17166 29004 17172 29006
rect 17236 29004 17242 29068
rect 17350 29004 17356 29068
rect 17420 29066 17467 29068
rect 17680 29066 17740 29142
rect 17861 29200 27863 29202
rect 17861 29144 17866 29200
rect 17922 29144 27802 29200
rect 27858 29144 27863 29200
rect 17861 29142 27863 29144
rect 17861 29139 17927 29142
rect 27797 29139 27863 29142
rect 28993 29202 29059 29205
rect 29200 29202 30000 29232
rect 28993 29200 30000 29202
rect 28993 29144 28998 29200
rect 29054 29144 30000 29200
rect 28993 29142 30000 29144
rect 28993 29139 29059 29142
rect 29200 29112 30000 29142
rect 20989 29066 21055 29069
rect 22277 29066 22343 29069
rect 27613 29066 27679 29069
rect 17420 29064 17512 29066
rect 17462 29008 17512 29064
rect 17420 29006 17512 29008
rect 17680 29064 22343 29066
rect 17680 29008 20994 29064
rect 21050 29008 22282 29064
rect 22338 29008 22343 29064
rect 17680 29006 22343 29008
rect 17420 29004 17467 29006
rect 17401 29003 17467 29004
rect 20989 29003 21055 29006
rect 22277 29003 22343 29006
rect 23430 29064 27679 29066
rect 23430 29008 27618 29064
rect 27674 29008 27679 29064
rect 23430 29006 27679 29008
rect 0 28840 800 28960
rect 14406 28868 14412 28932
rect 14476 28930 14482 28932
rect 15285 28930 15351 28933
rect 14476 28928 15351 28930
rect 14476 28872 15290 28928
rect 15346 28872 15351 28928
rect 14476 28870 15351 28872
rect 14476 28868 14482 28870
rect 15285 28867 15351 28870
rect 15745 28930 15811 28933
rect 17953 28930 18019 28933
rect 15745 28928 18019 28930
rect 15745 28872 15750 28928
rect 15806 28872 17958 28928
rect 18014 28872 18019 28928
rect 15745 28870 18019 28872
rect 15745 28867 15811 28870
rect 17953 28867 18019 28870
rect 18781 28930 18847 28933
rect 19425 28930 19491 28933
rect 18781 28928 19491 28930
rect 18781 28872 18786 28928
rect 18842 28872 19430 28928
rect 19486 28872 19491 28928
rect 18781 28870 19491 28872
rect 18781 28867 18847 28870
rect 19425 28867 19491 28870
rect 19701 28930 19767 28933
rect 20621 28930 20687 28933
rect 19701 28928 20687 28930
rect 19701 28872 19706 28928
rect 19762 28872 20626 28928
rect 20682 28872 20687 28928
rect 19701 28870 20687 28872
rect 19701 28867 19767 28870
rect 20621 28867 20687 28870
rect 22870 28868 22876 28932
rect 22940 28930 22946 28932
rect 23105 28930 23171 28933
rect 22940 28928 23171 28930
rect 22940 28872 23110 28928
rect 23166 28872 23171 28928
rect 22940 28870 23171 28872
rect 22940 28868 22946 28870
rect 23105 28867 23171 28870
rect 4419 28864 4735 28865
rect 4419 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4735 28864
rect 4419 28799 4735 28800
rect 11365 28864 11681 28865
rect 11365 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11681 28864
rect 11365 28799 11681 28800
rect 18311 28864 18627 28865
rect 18311 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18627 28864
rect 18311 28799 18627 28800
rect 17953 28794 18019 28797
rect 12390 28792 18019 28794
rect 12390 28736 17958 28792
rect 18014 28736 18019 28792
rect 12390 28734 18019 28736
rect 10869 28658 10935 28661
rect 12390 28658 12450 28734
rect 17953 28731 18019 28734
rect 19057 28794 19123 28797
rect 22829 28794 22895 28797
rect 19057 28792 22895 28794
rect 19057 28736 19062 28792
rect 19118 28736 22834 28792
rect 22890 28736 22895 28792
rect 19057 28734 22895 28736
rect 19057 28731 19123 28734
rect 22829 28731 22895 28734
rect 10869 28656 12450 28658
rect 10869 28600 10874 28656
rect 10930 28600 12450 28656
rect 10869 28598 12450 28600
rect 13261 28658 13327 28661
rect 23430 28658 23490 29006
rect 27613 29003 27679 29006
rect 23565 28930 23631 28933
rect 24945 28930 25011 28933
rect 23565 28928 25011 28930
rect 23565 28872 23570 28928
rect 23626 28872 24950 28928
rect 25006 28872 25011 28928
rect 23565 28870 25011 28872
rect 23565 28867 23631 28870
rect 24945 28867 25011 28870
rect 25257 28864 25573 28865
rect 25257 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25573 28864
rect 25257 28799 25573 28800
rect 13261 28656 23490 28658
rect 13261 28600 13266 28656
rect 13322 28600 23490 28656
rect 13261 28598 23490 28600
rect 23657 28658 23723 28661
rect 23790 28658 23796 28660
rect 23657 28656 23796 28658
rect 23657 28600 23662 28656
rect 23718 28600 23796 28656
rect 23657 28598 23796 28600
rect 10869 28595 10935 28598
rect 13261 28595 13327 28598
rect 23657 28595 23723 28598
rect 23790 28596 23796 28598
rect 23860 28658 23866 28660
rect 27521 28658 27587 28661
rect 23860 28656 27587 28658
rect 23860 28600 27526 28656
rect 27582 28600 27587 28656
rect 23860 28598 27587 28600
rect 23860 28596 23866 28598
rect 27521 28595 27587 28598
rect 12525 28522 12591 28525
rect 24710 28522 24716 28524
rect 12525 28520 24716 28522
rect 12525 28464 12530 28520
rect 12586 28464 24716 28520
rect 12525 28462 24716 28464
rect 12525 28459 12591 28462
rect 24710 28460 24716 28462
rect 24780 28460 24786 28524
rect 25405 28522 25471 28525
rect 25814 28522 25820 28524
rect 25405 28520 25820 28522
rect 25405 28464 25410 28520
rect 25466 28464 25820 28520
rect 25405 28462 25820 28464
rect 25405 28459 25471 28462
rect 25814 28460 25820 28462
rect 25884 28460 25890 28524
rect 28165 28522 28231 28525
rect 29200 28522 30000 28552
rect 28165 28520 30000 28522
rect 28165 28464 28170 28520
rect 28226 28464 30000 28520
rect 28165 28462 30000 28464
rect 28165 28459 28231 28462
rect 29200 28432 30000 28462
rect 11697 28386 11763 28389
rect 13813 28386 13879 28389
rect 11697 28384 13879 28386
rect 11697 28328 11702 28384
rect 11758 28328 13818 28384
rect 13874 28328 13879 28384
rect 11697 28326 13879 28328
rect 11697 28323 11763 28326
rect 13813 28323 13879 28326
rect 15469 28386 15535 28389
rect 16481 28386 16547 28389
rect 15469 28384 16547 28386
rect 15469 28328 15474 28384
rect 15530 28328 16486 28384
rect 16542 28328 16547 28384
rect 15469 28326 16547 28328
rect 15469 28323 15535 28326
rect 16481 28323 16547 28326
rect 17953 28386 18019 28389
rect 20069 28386 20135 28389
rect 17953 28384 20135 28386
rect 17953 28328 17958 28384
rect 18014 28328 20074 28384
rect 20130 28328 20135 28384
rect 17953 28326 20135 28328
rect 17953 28323 18019 28326
rect 20069 28323 20135 28326
rect 23013 28386 23079 28389
rect 23749 28386 23815 28389
rect 27470 28386 27476 28388
rect 23013 28384 27476 28386
rect 23013 28328 23018 28384
rect 23074 28328 23754 28384
rect 23810 28328 27476 28384
rect 23013 28326 27476 28328
rect 23013 28323 23079 28326
rect 23749 28323 23815 28326
rect 27470 28324 27476 28326
rect 27540 28324 27546 28388
rect 7892 28320 8208 28321
rect 0 28250 800 28280
rect 7892 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8208 28320
rect 7892 28255 8208 28256
rect 14838 28320 15154 28321
rect 14838 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15154 28320
rect 14838 28255 15154 28256
rect 21784 28320 22100 28321
rect 21784 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22100 28320
rect 21784 28255 22100 28256
rect 28730 28320 29046 28321
rect 28730 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29046 28320
rect 28730 28255 29046 28256
rect 1577 28250 1643 28253
rect 0 28248 1643 28250
rect 0 28192 1582 28248
rect 1638 28192 1643 28248
rect 0 28190 1643 28192
rect 0 28160 800 28190
rect 1577 28187 1643 28190
rect 12341 28250 12407 28253
rect 12985 28250 13051 28253
rect 12341 28248 13051 28250
rect 12341 28192 12346 28248
rect 12402 28192 12990 28248
rect 13046 28192 13051 28248
rect 12341 28190 13051 28192
rect 12341 28187 12407 28190
rect 12985 28187 13051 28190
rect 15377 28250 15443 28253
rect 15510 28250 15516 28252
rect 15377 28248 15516 28250
rect 15377 28192 15382 28248
rect 15438 28192 15516 28248
rect 15377 28190 15516 28192
rect 15377 28187 15443 28190
rect 15510 28188 15516 28190
rect 15580 28188 15586 28252
rect 16573 28250 16639 28253
rect 20253 28250 20319 28253
rect 20713 28250 20779 28253
rect 16573 28248 19442 28250
rect 16573 28192 16578 28248
rect 16634 28192 19442 28248
rect 16573 28190 19442 28192
rect 16573 28187 16639 28190
rect 11421 28114 11487 28117
rect 19241 28114 19307 28117
rect 11421 28112 19307 28114
rect 11421 28056 11426 28112
rect 11482 28056 19246 28112
rect 19302 28056 19307 28112
rect 11421 28054 19307 28056
rect 19382 28114 19442 28190
rect 20253 28248 20779 28250
rect 20253 28192 20258 28248
rect 20314 28192 20718 28248
rect 20774 28192 20779 28248
rect 20253 28190 20779 28192
rect 20253 28187 20319 28190
rect 20713 28187 20779 28190
rect 24526 28188 24532 28252
rect 24596 28250 24602 28252
rect 27337 28250 27403 28253
rect 24596 28248 27403 28250
rect 24596 28192 27342 28248
rect 27398 28192 27403 28248
rect 24596 28190 27403 28192
rect 24596 28188 24602 28190
rect 27337 28187 27403 28190
rect 27429 28114 27495 28117
rect 19382 28112 27495 28114
rect 19382 28056 27434 28112
rect 27490 28056 27495 28112
rect 19382 28054 27495 28056
rect 11421 28051 11487 28054
rect 19241 28051 19307 28054
rect 27429 28051 27495 28054
rect 13261 27978 13327 27981
rect 25313 27978 25379 27981
rect 13261 27976 24778 27978
rect 13261 27920 13266 27976
rect 13322 27920 24778 27976
rect 13261 27918 24778 27920
rect 13261 27915 13327 27918
rect 14457 27842 14523 27845
rect 17534 27842 17540 27844
rect 14457 27840 17540 27842
rect 14457 27784 14462 27840
rect 14518 27784 17540 27840
rect 14457 27782 17540 27784
rect 14457 27779 14523 27782
rect 17534 27780 17540 27782
rect 17604 27780 17610 27844
rect 18689 27842 18755 27845
rect 19333 27842 19399 27845
rect 20529 27842 20595 27845
rect 22277 27842 22343 27845
rect 18689 27840 19258 27842
rect 18689 27784 18694 27840
rect 18750 27784 19258 27840
rect 18689 27782 19258 27784
rect 18689 27779 18755 27782
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 12525 27706 12591 27709
rect 14181 27706 14247 27709
rect 12525 27704 14247 27706
rect 12525 27648 12530 27704
rect 12586 27648 14186 27704
rect 14242 27648 14247 27704
rect 12525 27646 14247 27648
rect 12525 27643 12591 27646
rect 14181 27643 14247 27646
rect 15193 27706 15259 27709
rect 15326 27706 15332 27708
rect 15193 27704 15332 27706
rect 15193 27648 15198 27704
rect 15254 27648 15332 27704
rect 15193 27646 15332 27648
rect 15193 27643 15259 27646
rect 15326 27644 15332 27646
rect 15396 27644 15402 27708
rect 15469 27706 15535 27709
rect 17493 27706 17559 27709
rect 15469 27704 17559 27706
rect 15469 27648 15474 27704
rect 15530 27648 17498 27704
rect 17554 27648 17559 27704
rect 15469 27646 17559 27648
rect 15469 27643 15535 27646
rect 17493 27643 17559 27646
rect 17769 27706 17835 27709
rect 17902 27706 17908 27708
rect 17769 27704 17908 27706
rect 17769 27648 17774 27704
rect 17830 27648 17908 27704
rect 17769 27646 17908 27648
rect 17769 27643 17835 27646
rect 17902 27644 17908 27646
rect 17972 27644 17978 27708
rect 19198 27706 19258 27782
rect 19333 27840 22343 27842
rect 19333 27784 19338 27840
rect 19394 27784 20534 27840
rect 20590 27784 22282 27840
rect 22338 27784 22343 27840
rect 19333 27782 22343 27784
rect 19333 27779 19399 27782
rect 20529 27779 20595 27782
rect 22277 27779 22343 27782
rect 22737 27842 22803 27845
rect 23289 27842 23355 27845
rect 23841 27842 23907 27845
rect 22737 27840 23907 27842
rect 22737 27784 22742 27840
rect 22798 27784 23294 27840
rect 23350 27784 23846 27840
rect 23902 27784 23907 27840
rect 22737 27782 23907 27784
rect 22737 27779 22803 27782
rect 23289 27779 23355 27782
rect 23841 27779 23907 27782
rect 19609 27706 19675 27709
rect 19198 27704 19675 27706
rect 19198 27648 19614 27704
rect 19670 27648 19675 27704
rect 19198 27646 19675 27648
rect 19609 27643 19675 27646
rect 20161 27706 20227 27709
rect 20294 27706 20300 27708
rect 20161 27704 20300 27706
rect 20161 27648 20166 27704
rect 20222 27648 20300 27704
rect 20161 27646 20300 27648
rect 20161 27643 20227 27646
rect 20294 27644 20300 27646
rect 20364 27644 20370 27708
rect 22553 27706 22619 27709
rect 20486 27704 22619 27706
rect 20486 27648 22558 27704
rect 22614 27648 22619 27704
rect 20486 27646 22619 27648
rect 0 27570 800 27600
rect 1577 27570 1643 27573
rect 0 27568 1643 27570
rect 0 27512 1582 27568
rect 1638 27512 1643 27568
rect 0 27510 1643 27512
rect 0 27480 800 27510
rect 1577 27507 1643 27510
rect 12065 27570 12131 27573
rect 20161 27570 20227 27573
rect 12065 27568 20227 27570
rect 12065 27512 12070 27568
rect 12126 27512 20166 27568
rect 20222 27512 20227 27568
rect 12065 27510 20227 27512
rect 12065 27507 12131 27510
rect 20161 27507 20227 27510
rect 20345 27570 20411 27573
rect 20486 27570 20546 27646
rect 22553 27643 22619 27646
rect 23105 27706 23171 27709
rect 23606 27706 23612 27708
rect 23105 27704 23612 27706
rect 23105 27648 23110 27704
rect 23166 27648 23612 27704
rect 23105 27646 23612 27648
rect 23105 27643 23171 27646
rect 23606 27644 23612 27646
rect 23676 27644 23682 27708
rect 20345 27568 20546 27570
rect 20345 27512 20350 27568
rect 20406 27512 20546 27568
rect 20345 27510 20546 27512
rect 20345 27507 20411 27510
rect 20662 27508 20668 27572
rect 20732 27570 20738 27572
rect 23105 27570 23171 27573
rect 20732 27568 23171 27570
rect 20732 27512 23110 27568
rect 23166 27512 23171 27568
rect 20732 27510 23171 27512
rect 20732 27508 20738 27510
rect 23105 27507 23171 27510
rect 23422 27508 23428 27572
rect 23492 27570 23498 27572
rect 23749 27570 23815 27573
rect 23492 27568 23815 27570
rect 23492 27512 23754 27568
rect 23810 27512 23815 27568
rect 23492 27510 23815 27512
rect 24718 27570 24778 27918
rect 25086 27976 25379 27978
rect 25086 27920 25318 27976
rect 25374 27920 25379 27976
rect 25086 27918 25379 27920
rect 25086 27709 25146 27918
rect 25313 27915 25379 27918
rect 25497 27978 25563 27981
rect 26182 27978 26188 27980
rect 25497 27976 26188 27978
rect 25497 27920 25502 27976
rect 25558 27920 26188 27976
rect 25497 27918 26188 27920
rect 25497 27915 25563 27918
rect 26182 27916 26188 27918
rect 26252 27916 26258 27980
rect 27470 27916 27476 27980
rect 27540 27978 27546 27980
rect 27797 27978 27863 27981
rect 27540 27976 27863 27978
rect 27540 27920 27802 27976
rect 27858 27920 27863 27976
rect 27540 27918 27863 27920
rect 27540 27916 27546 27918
rect 27797 27915 27863 27918
rect 26693 27842 26759 27845
rect 29200 27842 30000 27872
rect 26693 27840 30000 27842
rect 26693 27784 26698 27840
rect 26754 27784 30000 27840
rect 26693 27782 30000 27784
rect 26693 27779 26759 27782
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 29200 27752 30000 27782
rect 25257 27711 25573 27712
rect 25037 27704 25146 27709
rect 25037 27648 25042 27704
rect 25098 27648 25146 27704
rect 25037 27646 25146 27648
rect 25037 27643 25103 27646
rect 25681 27570 25747 27573
rect 24718 27568 25747 27570
rect 24718 27512 25686 27568
rect 25742 27512 25747 27568
rect 24718 27510 25747 27512
rect 23492 27508 23498 27510
rect 23749 27507 23815 27510
rect 25681 27507 25747 27510
rect 12433 27434 12499 27437
rect 25865 27434 25931 27437
rect 12433 27432 25931 27434
rect 12433 27376 12438 27432
rect 12494 27376 25870 27432
rect 25926 27376 25931 27432
rect 12433 27374 25931 27376
rect 12433 27371 12499 27374
rect 25865 27371 25931 27374
rect 13353 27298 13419 27301
rect 14457 27300 14523 27301
rect 13486 27298 13492 27300
rect 13353 27296 13492 27298
rect 13353 27240 13358 27296
rect 13414 27240 13492 27296
rect 13353 27238 13492 27240
rect 13353 27235 13419 27238
rect 13486 27236 13492 27238
rect 13556 27236 13562 27300
rect 14406 27236 14412 27300
rect 14476 27298 14523 27300
rect 15377 27298 15443 27301
rect 16021 27300 16087 27301
rect 15510 27298 15516 27300
rect 14476 27296 14568 27298
rect 14518 27240 14568 27296
rect 14476 27238 14568 27240
rect 15377 27296 15516 27298
rect 15377 27240 15382 27296
rect 15438 27240 15516 27296
rect 15377 27238 15516 27240
rect 14476 27236 14523 27238
rect 14457 27235 14523 27236
rect 15377 27235 15443 27238
rect 15510 27236 15516 27238
rect 15580 27236 15586 27300
rect 16021 27298 16068 27300
rect 15976 27296 16068 27298
rect 15976 27240 16026 27296
rect 15976 27238 16068 27240
rect 16021 27236 16068 27238
rect 16132 27236 16138 27300
rect 16614 27236 16620 27300
rect 16684 27298 16690 27300
rect 17401 27298 17467 27301
rect 16684 27296 17467 27298
rect 16684 27240 17406 27296
rect 17462 27240 17467 27296
rect 16684 27238 17467 27240
rect 16684 27236 16690 27238
rect 16021 27235 16087 27236
rect 17401 27235 17467 27238
rect 17677 27298 17743 27301
rect 20161 27298 20227 27301
rect 21357 27298 21423 27301
rect 17677 27296 21423 27298
rect 17677 27240 17682 27296
rect 17738 27240 20166 27296
rect 20222 27240 21362 27296
rect 21418 27240 21423 27296
rect 17677 27238 21423 27240
rect 17677 27235 17743 27238
rect 20161 27235 20227 27238
rect 21357 27235 21423 27238
rect 22686 27236 22692 27300
rect 22756 27298 22762 27300
rect 28257 27298 28323 27301
rect 22756 27296 28323 27298
rect 22756 27240 28262 27296
rect 28318 27240 28323 27296
rect 22756 27238 28323 27240
rect 22756 27236 22762 27238
rect 28257 27235 28323 27238
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 15878 27100 15884 27164
rect 15948 27162 15954 27164
rect 16297 27162 16363 27165
rect 15948 27160 16363 27162
rect 15948 27104 16302 27160
rect 16358 27104 16363 27160
rect 15948 27102 16363 27104
rect 15948 27100 15954 27102
rect 16297 27099 16363 27102
rect 16757 27162 16823 27165
rect 20713 27162 20779 27165
rect 16757 27160 20779 27162
rect 16757 27104 16762 27160
rect 16818 27104 20718 27160
rect 20774 27104 20779 27160
rect 16757 27102 20779 27104
rect 16757 27099 16823 27102
rect 20713 27099 20779 27102
rect 22318 27100 22324 27164
rect 22388 27162 22394 27164
rect 22553 27162 22619 27165
rect 22388 27160 22619 27162
rect 22388 27104 22558 27160
rect 22614 27104 22619 27160
rect 22388 27102 22619 27104
rect 22388 27100 22394 27102
rect 22553 27099 22619 27102
rect 23105 27162 23171 27165
rect 24894 27162 24900 27164
rect 23105 27160 24900 27162
rect 23105 27104 23110 27160
rect 23166 27104 24900 27160
rect 23105 27102 24900 27104
rect 23105 27099 23171 27102
rect 24894 27100 24900 27102
rect 24964 27162 24970 27164
rect 25497 27162 25563 27165
rect 24964 27160 25563 27162
rect 24964 27104 25502 27160
rect 25558 27104 25563 27160
rect 29200 27128 30000 27192
rect 24964 27102 25563 27104
rect 24964 27100 24970 27102
rect 25497 27099 25563 27102
rect 29134 27072 30000 27128
rect 29134 27068 29378 27072
rect 8293 27026 8359 27029
rect 9397 27026 9463 27029
rect 22001 27026 22067 27029
rect 22553 27026 22619 27029
rect 24393 27026 24459 27029
rect 8293 27024 24459 27026
rect 8293 26968 8298 27024
rect 8354 26968 9402 27024
rect 9458 26968 22006 27024
rect 22062 26968 22558 27024
rect 22614 26968 24398 27024
rect 24454 26968 24459 27024
rect 8293 26966 24459 26968
rect 8293 26963 8359 26966
rect 9397 26963 9463 26966
rect 22001 26963 22067 26966
rect 22553 26963 22619 26966
rect 24393 26963 24459 26966
rect 24710 26964 24716 27028
rect 24780 27026 24786 27028
rect 27153 27026 27219 27029
rect 24780 27024 27219 27026
rect 24780 26968 27158 27024
rect 27214 26968 27219 27024
rect 24780 26966 27219 26968
rect 24780 26964 24786 26966
rect 27153 26963 27219 26966
rect 28625 27026 28691 27029
rect 29134 27026 29194 27068
rect 28625 27024 29194 27026
rect 28625 26968 28630 27024
rect 28686 26968 29194 27024
rect 28625 26966 29194 26968
rect 28625 26963 28691 26966
rect 0 26800 800 26920
rect 14365 26890 14431 26893
rect 21449 26890 21515 26893
rect 14365 26888 21515 26890
rect 14365 26832 14370 26888
rect 14426 26832 21454 26888
rect 21510 26832 21515 26888
rect 14365 26830 21515 26832
rect 14365 26827 14431 26830
rect 21449 26827 21515 26830
rect 21725 26890 21791 26893
rect 23381 26890 23447 26893
rect 21725 26888 23447 26890
rect 21725 26832 21730 26888
rect 21786 26832 23386 26888
rect 23442 26832 23447 26888
rect 21725 26830 23447 26832
rect 21725 26827 21791 26830
rect 23381 26827 23447 26830
rect 25078 26828 25084 26892
rect 25148 26890 25154 26892
rect 25221 26890 25287 26893
rect 25148 26888 25287 26890
rect 25148 26832 25226 26888
rect 25282 26832 25287 26888
rect 25148 26830 25287 26832
rect 25148 26828 25154 26830
rect 25221 26827 25287 26830
rect 25630 26828 25636 26892
rect 25700 26890 25706 26892
rect 25773 26890 25839 26893
rect 25700 26888 25839 26890
rect 25700 26832 25778 26888
rect 25834 26832 25839 26888
rect 25700 26830 25839 26832
rect 25700 26828 25706 26830
rect 25773 26827 25839 26830
rect 26601 26890 26667 26893
rect 27613 26890 27679 26893
rect 26601 26888 27679 26890
rect 26601 26832 26606 26888
rect 26662 26832 27618 26888
rect 27674 26832 27679 26888
rect 26601 26830 27679 26832
rect 26601 26827 26667 26830
rect 27613 26827 27679 26830
rect 12985 26754 13051 26757
rect 14825 26754 14891 26757
rect 15285 26754 15351 26757
rect 12985 26752 15351 26754
rect 12985 26696 12990 26752
rect 13046 26696 14830 26752
rect 14886 26696 15290 26752
rect 15346 26696 15351 26752
rect 12985 26694 15351 26696
rect 12985 26691 13051 26694
rect 14825 26691 14891 26694
rect 15285 26691 15351 26694
rect 15929 26754 15995 26757
rect 17769 26754 17835 26757
rect 19241 26756 19307 26757
rect 20713 26756 20779 26757
rect 19190 26754 19196 26756
rect 15929 26752 17835 26754
rect 15929 26696 15934 26752
rect 15990 26696 17774 26752
rect 17830 26696 17835 26752
rect 15929 26694 17835 26696
rect 19150 26694 19196 26754
rect 19260 26752 19307 26756
rect 20662 26754 20668 26756
rect 19302 26696 19307 26752
rect 15929 26691 15995 26694
rect 17769 26691 17835 26694
rect 19190 26692 19196 26694
rect 19260 26692 19307 26696
rect 20586 26694 20668 26754
rect 20732 26754 20779 26756
rect 24945 26754 25011 26757
rect 20732 26752 25011 26754
rect 20774 26696 24950 26752
rect 25006 26696 25011 26752
rect 20662 26692 20668 26694
rect 20732 26694 25011 26696
rect 20732 26692 20779 26694
rect 19241 26691 19307 26692
rect 20713 26691 20779 26692
rect 24945 26691 25011 26694
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 15101 26618 15167 26621
rect 15469 26618 15535 26621
rect 15101 26616 15535 26618
rect 15101 26560 15106 26616
rect 15162 26560 15474 26616
rect 15530 26560 15535 26616
rect 15101 26558 15535 26560
rect 15101 26555 15167 26558
rect 15469 26555 15535 26558
rect 15929 26618 15995 26621
rect 16113 26618 16179 26621
rect 15929 26616 16179 26618
rect 15929 26560 15934 26616
rect 15990 26560 16118 26616
rect 16174 26560 16179 26616
rect 15929 26558 16179 26560
rect 15929 26555 15995 26558
rect 16113 26555 16179 26558
rect 16665 26618 16731 26621
rect 17861 26618 17927 26621
rect 16665 26616 17927 26618
rect 16665 26560 16670 26616
rect 16726 26560 17866 26616
rect 17922 26560 17927 26616
rect 16665 26558 17927 26560
rect 16665 26555 16731 26558
rect 17861 26555 17927 26558
rect 19701 26618 19767 26621
rect 21173 26618 21239 26621
rect 19701 26616 21239 26618
rect 19701 26560 19706 26616
rect 19762 26560 21178 26616
rect 21234 26560 21239 26616
rect 19701 26558 21239 26560
rect 19701 26555 19767 26558
rect 21173 26555 21239 26558
rect 22093 26618 22159 26621
rect 23289 26618 23355 26621
rect 22093 26616 23355 26618
rect 22093 26560 22098 26616
rect 22154 26560 23294 26616
rect 23350 26560 23355 26616
rect 22093 26558 23355 26560
rect 22093 26555 22159 26558
rect 23289 26555 23355 26558
rect 25681 26618 25747 26621
rect 25957 26618 26023 26621
rect 25681 26616 26023 26618
rect 25681 26560 25686 26616
rect 25742 26560 25962 26616
rect 26018 26560 26023 26616
rect 25681 26558 26023 26560
rect 25681 26555 25747 26558
rect 25957 26555 26023 26558
rect 10409 26482 10475 26485
rect 20713 26482 20779 26485
rect 10409 26480 20779 26482
rect 10409 26424 10414 26480
rect 10470 26424 20718 26480
rect 20774 26424 20779 26480
rect 10409 26422 20779 26424
rect 10409 26419 10475 26422
rect 20713 26419 20779 26422
rect 20846 26420 20852 26484
rect 20916 26482 20922 26484
rect 23657 26482 23723 26485
rect 20916 26480 23723 26482
rect 20916 26424 23662 26480
rect 23718 26424 23723 26480
rect 20916 26422 23723 26424
rect 20916 26420 20922 26422
rect 23657 26419 23723 26422
rect 24342 26420 24348 26484
rect 24412 26482 24418 26484
rect 26141 26482 26207 26485
rect 24412 26480 26207 26482
rect 24412 26424 26146 26480
rect 26202 26424 26207 26480
rect 24412 26422 26207 26424
rect 24412 26420 24418 26422
rect 26141 26419 26207 26422
rect 28022 26420 28028 26484
rect 28092 26482 28098 26484
rect 29200 26482 30000 26512
rect 28092 26422 30000 26482
rect 28092 26420 28098 26422
rect 29200 26392 30000 26422
rect 9857 26346 9923 26349
rect 13261 26346 13327 26349
rect 9857 26344 13327 26346
rect 9857 26288 9862 26344
rect 9918 26288 13266 26344
rect 13322 26288 13327 26344
rect 9857 26286 13327 26288
rect 9857 26283 9923 26286
rect 13261 26283 13327 26286
rect 14641 26346 14707 26349
rect 16614 26346 16620 26348
rect 14641 26344 16620 26346
rect 14641 26288 14646 26344
rect 14702 26288 16620 26344
rect 14641 26286 16620 26288
rect 14641 26283 14707 26286
rect 16614 26284 16620 26286
rect 16684 26284 16690 26348
rect 17493 26346 17559 26349
rect 17861 26346 17927 26349
rect 19057 26346 19123 26349
rect 17493 26344 17740 26346
rect 17493 26288 17498 26344
rect 17554 26288 17740 26344
rect 17493 26286 17740 26288
rect 17493 26283 17559 26286
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 16113 26212 16179 26213
rect 16062 26210 16068 26212
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 16022 26150 16068 26210
rect 16132 26208 16179 26212
rect 16174 26152 16179 26208
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 16062 26148 16068 26150
rect 16132 26148 16179 26152
rect 16113 26147 16179 26148
rect 16481 26210 16547 26213
rect 17493 26210 17559 26213
rect 16481 26208 17559 26210
rect 16481 26152 16486 26208
rect 16542 26152 17498 26208
rect 17554 26152 17559 26208
rect 16481 26150 17559 26152
rect 17680 26210 17740 26286
rect 17861 26344 19123 26346
rect 17861 26288 17866 26344
rect 17922 26288 19062 26344
rect 19118 26288 19123 26344
rect 17861 26286 19123 26288
rect 17861 26283 17927 26286
rect 19057 26283 19123 26286
rect 19793 26346 19859 26349
rect 26417 26346 26483 26349
rect 19793 26344 26483 26346
rect 19793 26288 19798 26344
rect 19854 26288 26422 26344
rect 26478 26288 26483 26344
rect 19793 26286 26483 26288
rect 19793 26283 19859 26286
rect 26417 26283 26483 26286
rect 21173 26210 21239 26213
rect 17680 26208 21239 26210
rect 17680 26152 21178 26208
rect 21234 26152 21239 26208
rect 17680 26150 21239 26152
rect 16481 26147 16547 26150
rect 17493 26147 17559 26150
rect 21173 26147 21239 26150
rect 23105 26210 23171 26213
rect 23790 26210 23796 26212
rect 23105 26208 23796 26210
rect 23105 26152 23110 26208
rect 23166 26152 23796 26208
rect 23105 26150 23796 26152
rect 23105 26147 23171 26150
rect 23790 26148 23796 26150
rect 23860 26148 23866 26212
rect 23974 26148 23980 26212
rect 24044 26210 24050 26212
rect 25129 26210 25195 26213
rect 24044 26208 25195 26210
rect 24044 26152 25134 26208
rect 25190 26152 25195 26208
rect 24044 26150 25195 26152
rect 24044 26148 24050 26150
rect 25129 26147 25195 26150
rect 25313 26210 25379 26213
rect 27705 26210 27771 26213
rect 25313 26208 27771 26210
rect 25313 26152 25318 26208
rect 25374 26152 27710 26208
rect 27766 26152 27771 26208
rect 25313 26150 27771 26152
rect 25313 26147 25379 26150
rect 27705 26147 27771 26150
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 16757 26074 16823 26077
rect 17217 26074 17283 26077
rect 16757 26072 17283 26074
rect 16757 26016 16762 26072
rect 16818 26016 17222 26072
rect 17278 26016 17283 26072
rect 16757 26014 17283 26016
rect 16757 26011 16823 26014
rect 17217 26011 17283 26014
rect 17534 26012 17540 26076
rect 17604 26074 17610 26076
rect 18689 26074 18755 26077
rect 17604 26072 18755 26074
rect 17604 26016 18694 26072
rect 18750 26016 18755 26072
rect 17604 26014 18755 26016
rect 17604 26012 17610 26014
rect 18689 26011 18755 26014
rect 19374 26012 19380 26076
rect 19444 26074 19450 26076
rect 19517 26074 19583 26077
rect 19444 26072 19583 26074
rect 19444 26016 19522 26072
rect 19578 26016 19583 26072
rect 19444 26014 19583 26016
rect 19444 26012 19450 26014
rect 19517 26011 19583 26014
rect 19742 26012 19748 26076
rect 19812 26074 19818 26076
rect 21541 26074 21607 26077
rect 19812 26072 21607 26074
rect 19812 26016 21546 26072
rect 21602 26016 21607 26072
rect 19812 26014 21607 26016
rect 19812 26012 19818 26014
rect 21541 26011 21607 26014
rect 23054 26012 23060 26076
rect 23124 26074 23130 26076
rect 23381 26074 23447 26077
rect 23124 26072 23447 26074
rect 23124 26016 23386 26072
rect 23442 26016 23447 26072
rect 23124 26014 23447 26016
rect 23124 26012 23130 26014
rect 23381 26011 23447 26014
rect 24577 26074 24643 26077
rect 25078 26074 25084 26076
rect 24577 26072 25084 26074
rect 24577 26016 24582 26072
rect 24638 26016 25084 26072
rect 24577 26014 25084 26016
rect 24577 26011 24643 26014
rect 25078 26012 25084 26014
rect 25148 26074 25154 26076
rect 25221 26074 25287 26077
rect 25148 26072 25287 26074
rect 25148 26016 25226 26072
rect 25282 26016 25287 26072
rect 25148 26014 25287 26016
rect 25148 26012 25154 26014
rect 25221 26011 25287 26014
rect 26366 26012 26372 26076
rect 26436 26074 26442 26076
rect 27521 26074 27587 26077
rect 26436 26072 27587 26074
rect 26436 26016 27526 26072
rect 27582 26016 27587 26072
rect 26436 26014 27587 26016
rect 26436 26012 26442 26014
rect 27521 26011 27587 26014
rect 12893 25938 12959 25941
rect 14733 25938 14799 25941
rect 12893 25936 14799 25938
rect 12893 25880 12898 25936
rect 12954 25880 14738 25936
rect 14794 25880 14799 25936
rect 12893 25878 14799 25880
rect 12893 25875 12959 25878
rect 14733 25875 14799 25878
rect 16849 25938 16915 25941
rect 16849 25936 19810 25938
rect 16849 25880 16854 25936
rect 16910 25880 19810 25936
rect 16849 25878 19810 25880
rect 16849 25875 16915 25878
rect 10910 25740 10916 25804
rect 10980 25802 10986 25804
rect 19057 25802 19123 25805
rect 19333 25802 19399 25805
rect 10980 25742 18890 25802
rect 10980 25740 10986 25742
rect 16389 25666 16455 25669
rect 17677 25666 17743 25669
rect 16389 25664 17743 25666
rect 16389 25608 16394 25664
rect 16450 25608 17682 25664
rect 17738 25608 17743 25664
rect 16389 25606 17743 25608
rect 18830 25666 18890 25742
rect 19057 25800 19399 25802
rect 19057 25744 19062 25800
rect 19118 25744 19338 25800
rect 19394 25744 19399 25800
rect 19057 25742 19399 25744
rect 19750 25802 19810 25878
rect 19926 25876 19932 25940
rect 19996 25938 20002 25940
rect 20069 25938 20135 25941
rect 19996 25936 20135 25938
rect 19996 25880 20074 25936
rect 20130 25880 20135 25936
rect 19996 25878 20135 25880
rect 19996 25876 20002 25878
rect 20069 25875 20135 25878
rect 20478 25876 20484 25940
rect 20548 25938 20554 25940
rect 20805 25938 20871 25941
rect 20548 25936 20871 25938
rect 20548 25880 20810 25936
rect 20866 25880 20871 25936
rect 20548 25878 20871 25880
rect 20548 25876 20554 25878
rect 20805 25875 20871 25878
rect 21449 25938 21515 25941
rect 26509 25938 26575 25941
rect 21449 25936 26575 25938
rect 21449 25880 21454 25936
rect 21510 25880 26514 25936
rect 26570 25880 26575 25936
rect 21449 25878 26575 25880
rect 21449 25875 21515 25878
rect 26509 25875 26575 25878
rect 27153 25802 27219 25805
rect 19750 25800 27219 25802
rect 19750 25744 27158 25800
rect 27214 25744 27219 25800
rect 19750 25742 27219 25744
rect 19057 25739 19123 25742
rect 19333 25739 19399 25742
rect 27153 25739 27219 25742
rect 27889 25802 27955 25805
rect 29200 25802 30000 25832
rect 27889 25800 30000 25802
rect 27889 25744 27894 25800
rect 27950 25744 30000 25800
rect 27889 25742 30000 25744
rect 27889 25739 27955 25742
rect 29200 25712 30000 25742
rect 25078 25666 25084 25668
rect 18830 25606 25084 25666
rect 16389 25603 16455 25606
rect 17677 25603 17743 25606
rect 25078 25604 25084 25606
rect 25148 25604 25154 25668
rect 4419 25600 4735 25601
rect 0 25530 800 25560
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 1577 25530 1643 25533
rect 0 25528 1643 25530
rect 0 25472 1582 25528
rect 1638 25472 1643 25528
rect 0 25470 1643 25472
rect 0 25440 800 25470
rect 1577 25467 1643 25470
rect 17493 25530 17559 25533
rect 17769 25530 17835 25533
rect 17493 25528 17835 25530
rect 17493 25472 17498 25528
rect 17554 25472 17774 25528
rect 17830 25472 17835 25528
rect 17493 25470 17835 25472
rect 17493 25467 17559 25470
rect 17769 25467 17835 25470
rect 18689 25530 18755 25533
rect 21357 25530 21423 25533
rect 18689 25528 21423 25530
rect 18689 25472 18694 25528
rect 18750 25472 21362 25528
rect 21418 25472 21423 25528
rect 18689 25470 21423 25472
rect 18689 25467 18755 25470
rect 21357 25467 21423 25470
rect 22093 25530 22159 25533
rect 22461 25530 22527 25533
rect 22093 25528 22527 25530
rect 22093 25472 22098 25528
rect 22154 25472 22466 25528
rect 22522 25472 22527 25528
rect 22093 25470 22527 25472
rect 22093 25467 22159 25470
rect 22461 25467 22527 25470
rect 24853 25530 24919 25533
rect 25129 25530 25195 25533
rect 24853 25528 25195 25530
rect 24853 25472 24858 25528
rect 24914 25472 25134 25528
rect 25190 25472 25195 25528
rect 24853 25470 25195 25472
rect 24853 25467 24919 25470
rect 25129 25467 25195 25470
rect 25865 25530 25931 25533
rect 25998 25530 26004 25532
rect 25865 25528 26004 25530
rect 25865 25472 25870 25528
rect 25926 25472 26004 25528
rect 25865 25470 26004 25472
rect 25865 25467 25931 25470
rect 25998 25468 26004 25470
rect 26068 25468 26074 25532
rect 14590 25332 14596 25396
rect 14660 25394 14666 25396
rect 24945 25394 25011 25397
rect 14660 25392 25011 25394
rect 14660 25336 24950 25392
rect 25006 25336 25011 25392
rect 14660 25334 25011 25336
rect 14660 25332 14666 25334
rect 24945 25331 25011 25334
rect 25221 25394 25287 25397
rect 25814 25394 25820 25396
rect 25221 25392 25820 25394
rect 25221 25336 25226 25392
rect 25282 25336 25820 25392
rect 25221 25334 25820 25336
rect 25221 25331 25287 25334
rect 25814 25332 25820 25334
rect 25884 25332 25890 25396
rect 26182 25332 26188 25396
rect 26252 25394 26258 25396
rect 27797 25394 27863 25397
rect 26252 25392 27863 25394
rect 26252 25336 27802 25392
rect 27858 25336 27863 25392
rect 26252 25334 27863 25336
rect 26252 25332 26258 25334
rect 27797 25331 27863 25334
rect 13997 25258 14063 25261
rect 17217 25258 17283 25261
rect 26601 25258 26667 25261
rect 13997 25256 15394 25258
rect 13997 25200 14002 25256
rect 14058 25200 15394 25256
rect 13997 25198 15394 25200
rect 13997 25195 14063 25198
rect 15334 25122 15394 25198
rect 17217 25256 26667 25258
rect 17217 25200 17222 25256
rect 17278 25200 26606 25256
rect 26662 25200 26667 25256
rect 17217 25198 26667 25200
rect 17217 25195 17283 25198
rect 26601 25195 26667 25198
rect 19701 25122 19767 25125
rect 19977 25124 20043 25125
rect 19926 25122 19932 25124
rect 15334 25120 19767 25122
rect 15334 25064 19706 25120
rect 19762 25064 19767 25120
rect 15334 25062 19767 25064
rect 19886 25062 19932 25122
rect 19996 25120 20043 25124
rect 20038 25064 20043 25120
rect 19701 25059 19767 25062
rect 19926 25060 19932 25062
rect 19996 25060 20043 25064
rect 19977 25059 20043 25060
rect 20161 25122 20227 25125
rect 21633 25122 21699 25125
rect 20161 25120 21699 25122
rect 20161 25064 20166 25120
rect 20222 25064 21638 25120
rect 21694 25064 21699 25120
rect 20161 25062 21699 25064
rect 20161 25059 20227 25062
rect 21633 25059 21699 25062
rect 22829 25122 22895 25125
rect 27521 25122 27587 25125
rect 22829 25120 27587 25122
rect 22829 25064 22834 25120
rect 22890 25064 27526 25120
rect 27582 25064 27587 25120
rect 22829 25062 27587 25064
rect 22829 25059 22895 25062
rect 27521 25059 27587 25062
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 29200 25032 30000 25152
rect 28730 24991 29046 24992
rect 16614 24924 16620 24988
rect 16684 24986 16690 24988
rect 20805 24986 20871 24989
rect 23289 24988 23355 24989
rect 16684 24984 20871 24986
rect 16684 24928 20810 24984
rect 20866 24928 20871 24984
rect 16684 24926 20871 24928
rect 16684 24924 16690 24926
rect 20805 24923 20871 24926
rect 23238 24924 23244 24988
rect 23308 24986 23355 24988
rect 23308 24984 23400 24986
rect 23350 24928 23400 24984
rect 23308 24926 23400 24928
rect 25865 24984 25931 24989
rect 25865 24928 25870 24984
rect 25926 24928 25931 24984
rect 23308 24924 23355 24926
rect 23289 24923 23355 24924
rect 25865 24923 25931 24928
rect 26325 24986 26391 24989
rect 27337 24986 27403 24989
rect 26325 24984 27403 24986
rect 26325 24928 26330 24984
rect 26386 24928 27342 24984
rect 27398 24928 27403 24984
rect 26325 24926 27403 24928
rect 26325 24923 26391 24926
rect 27337 24923 27403 24926
rect 0 24760 800 24880
rect 14089 24850 14155 24853
rect 17677 24850 17743 24853
rect 14089 24848 17743 24850
rect 14089 24792 14094 24848
rect 14150 24792 17682 24848
rect 17738 24792 17743 24848
rect 14089 24790 17743 24792
rect 14089 24787 14155 24790
rect 17677 24787 17743 24790
rect 18689 24850 18755 24853
rect 18822 24850 18828 24852
rect 18689 24848 18828 24850
rect 18689 24792 18694 24848
rect 18750 24792 18828 24848
rect 18689 24790 18828 24792
rect 18689 24787 18755 24790
rect 18822 24788 18828 24790
rect 18892 24788 18898 24852
rect 19057 24850 19123 24853
rect 24526 24850 24532 24852
rect 19057 24848 24532 24850
rect 19057 24792 19062 24848
rect 19118 24792 24532 24848
rect 19057 24790 24532 24792
rect 19057 24787 19123 24790
rect 24526 24788 24532 24790
rect 24596 24788 24602 24852
rect 25868 24850 25928 24923
rect 29502 24870 29562 25032
rect 25998 24850 26004 24852
rect 25868 24790 26004 24850
rect 25998 24788 26004 24790
rect 26068 24788 26074 24852
rect 27705 24850 27771 24853
rect 29134 24850 29562 24870
rect 27705 24848 29562 24850
rect 27705 24792 27710 24848
rect 27766 24810 29562 24848
rect 27766 24792 29194 24810
rect 27705 24790 29194 24792
rect 27705 24787 27771 24790
rect 16573 24714 16639 24717
rect 17217 24714 17283 24717
rect 16573 24712 17283 24714
rect 16573 24656 16578 24712
rect 16634 24656 17222 24712
rect 17278 24656 17283 24712
rect 16573 24654 17283 24656
rect 16573 24651 16639 24654
rect 17217 24651 17283 24654
rect 17718 24652 17724 24716
rect 17788 24714 17794 24716
rect 18045 24714 18111 24717
rect 17788 24712 18111 24714
rect 17788 24656 18050 24712
rect 18106 24656 18111 24712
rect 17788 24654 18111 24656
rect 17788 24652 17794 24654
rect 18045 24651 18111 24654
rect 18505 24714 18571 24717
rect 24945 24714 25011 24717
rect 18505 24712 25011 24714
rect 18505 24656 18510 24712
rect 18566 24656 24950 24712
rect 25006 24656 25011 24712
rect 18505 24654 25011 24656
rect 18505 24651 18571 24654
rect 24945 24651 25011 24654
rect 25078 24652 25084 24716
rect 25148 24714 25154 24716
rect 25773 24714 25839 24717
rect 25148 24712 25839 24714
rect 25148 24656 25778 24712
rect 25834 24656 25839 24712
rect 25148 24654 25839 24656
rect 25148 24652 25154 24654
rect 25773 24651 25839 24654
rect 16481 24578 16547 24581
rect 17585 24578 17651 24581
rect 19742 24578 19748 24580
rect 16481 24576 17651 24578
rect 16481 24520 16486 24576
rect 16542 24520 17590 24576
rect 17646 24520 17651 24576
rect 16481 24518 17651 24520
rect 16481 24515 16547 24518
rect 17585 24515 17651 24518
rect 19566 24518 19748 24578
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 19425 24442 19491 24445
rect 19566 24442 19626 24518
rect 19742 24516 19748 24518
rect 19812 24516 19818 24580
rect 20069 24578 20135 24581
rect 24577 24578 24643 24581
rect 20069 24576 24643 24578
rect 20069 24520 20074 24576
rect 20130 24520 24582 24576
rect 24638 24520 24643 24576
rect 20069 24518 24643 24520
rect 20069 24515 20135 24518
rect 24577 24515 24643 24518
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 19425 24440 19626 24442
rect 19425 24384 19430 24440
rect 19486 24384 19626 24440
rect 19425 24382 19626 24384
rect 19793 24442 19859 24445
rect 20713 24442 20779 24445
rect 19793 24440 20779 24442
rect 19793 24384 19798 24440
rect 19854 24384 20718 24440
rect 20774 24384 20779 24440
rect 19793 24382 20779 24384
rect 19425 24379 19491 24382
rect 19793 24379 19859 24382
rect 20713 24379 20779 24382
rect 21173 24442 21239 24445
rect 22829 24442 22895 24445
rect 24117 24442 24183 24445
rect 25773 24442 25839 24445
rect 21173 24440 22754 24442
rect 21173 24384 21178 24440
rect 21234 24384 22754 24440
rect 21173 24382 22754 24384
rect 21173 24379 21239 24382
rect 13077 24306 13143 24309
rect 20805 24306 20871 24309
rect 13077 24304 20871 24306
rect 13077 24248 13082 24304
rect 13138 24248 20810 24304
rect 20866 24248 20871 24304
rect 13077 24246 20871 24248
rect 22694 24306 22754 24382
rect 22829 24440 24183 24442
rect 22829 24384 22834 24440
rect 22890 24384 24122 24440
rect 24178 24384 24183 24440
rect 22829 24382 24183 24384
rect 22829 24379 22895 24382
rect 24117 24379 24183 24382
rect 25638 24440 25839 24442
rect 25638 24384 25778 24440
rect 25834 24384 25839 24440
rect 25638 24382 25839 24384
rect 25129 24306 25195 24309
rect 22694 24304 25195 24306
rect 22694 24248 25134 24304
rect 25190 24248 25195 24304
rect 22694 24246 25195 24248
rect 13077 24243 13143 24246
rect 20805 24243 20871 24246
rect 25129 24243 25195 24246
rect 25405 24306 25471 24309
rect 25638 24306 25698 24382
rect 25773 24379 25839 24382
rect 28165 24442 28231 24445
rect 29200 24442 30000 24472
rect 28165 24440 30000 24442
rect 28165 24384 28170 24440
rect 28226 24384 30000 24440
rect 28165 24382 30000 24384
rect 28165 24379 28231 24382
rect 29200 24352 30000 24382
rect 25405 24304 25698 24306
rect 25405 24248 25410 24304
rect 25466 24248 25698 24304
rect 25405 24246 25698 24248
rect 27245 24306 27311 24309
rect 27521 24308 27587 24309
rect 27245 24304 27354 24306
rect 27245 24248 27250 24304
rect 27306 24248 27354 24304
rect 25405 24243 25471 24246
rect 27245 24243 27354 24248
rect 27470 24244 27476 24308
rect 27540 24306 27587 24308
rect 27540 24304 27632 24306
rect 27582 24248 27632 24304
rect 27540 24246 27632 24248
rect 27540 24244 27587 24246
rect 27521 24243 27587 24244
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 14457 24170 14523 24173
rect 20253 24170 20319 24173
rect 22829 24170 22895 24173
rect 14457 24168 20319 24170
rect 14457 24112 14462 24168
rect 14518 24112 20258 24168
rect 20314 24112 20319 24168
rect 14457 24110 20319 24112
rect 14457 24107 14523 24110
rect 20253 24107 20319 24110
rect 20486 24168 22895 24170
rect 20486 24112 22834 24168
rect 22890 24112 22895 24168
rect 20486 24110 22895 24112
rect 16113 24034 16179 24037
rect 20345 24034 20411 24037
rect 16113 24032 20411 24034
rect 16113 23976 16118 24032
rect 16174 23976 20350 24032
rect 20406 23976 20411 24032
rect 16113 23974 20411 23976
rect 16113 23971 16179 23974
rect 20345 23971 20411 23974
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 20110 23898 20116 23900
rect 15334 23838 20116 23898
rect 13486 23700 13492 23764
rect 13556 23762 13562 23764
rect 15334 23762 15394 23838
rect 20110 23836 20116 23838
rect 20180 23898 20186 23900
rect 20486 23898 20546 24110
rect 22829 24107 22895 24110
rect 23197 24170 23263 24173
rect 27153 24170 27219 24173
rect 23197 24168 27219 24170
rect 23197 24112 23202 24168
rect 23258 24112 27158 24168
rect 27214 24112 27219 24168
rect 23197 24110 27219 24112
rect 23197 24107 23263 24110
rect 27153 24107 27219 24110
rect 21265 24034 21331 24037
rect 21633 24034 21699 24037
rect 21265 24032 21699 24034
rect 21265 23976 21270 24032
rect 21326 23976 21638 24032
rect 21694 23976 21699 24032
rect 21265 23974 21699 23976
rect 21265 23971 21331 23974
rect 21633 23971 21699 23974
rect 22686 23972 22692 24036
rect 22756 24034 22762 24036
rect 22829 24034 22895 24037
rect 25129 24036 25195 24037
rect 22756 24032 22895 24034
rect 22756 23976 22834 24032
rect 22890 23976 22895 24032
rect 22756 23974 22895 23976
rect 22756 23972 22762 23974
rect 22829 23971 22895 23974
rect 25078 23972 25084 24036
rect 25148 24034 25195 24036
rect 26366 24034 26372 24036
rect 25148 24032 25240 24034
rect 25190 23976 25240 24032
rect 25148 23974 25240 23976
rect 25316 23974 26372 24034
rect 25148 23972 25195 23974
rect 25129 23971 25195 23972
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 20180 23838 20546 23898
rect 20621 23898 20687 23901
rect 20897 23898 20963 23901
rect 20621 23896 20963 23898
rect 20621 23840 20626 23896
rect 20682 23840 20902 23896
rect 20958 23840 20963 23896
rect 20621 23838 20963 23840
rect 20180 23836 20186 23838
rect 20621 23835 20687 23838
rect 20897 23835 20963 23838
rect 22185 23898 22251 23901
rect 25316 23898 25376 23974
rect 26366 23972 26372 23974
rect 26436 23972 26442 24036
rect 27153 24034 27219 24037
rect 27294 24034 27354 24243
rect 27153 24032 27354 24034
rect 27153 23976 27158 24032
rect 27214 23976 27354 24032
rect 27153 23974 27354 23976
rect 27153 23971 27219 23974
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 22185 23896 25376 23898
rect 22185 23840 22190 23896
rect 22246 23840 25376 23896
rect 22185 23838 25376 23840
rect 25589 23898 25655 23901
rect 26233 23900 26299 23901
rect 25814 23898 25820 23900
rect 25589 23896 25820 23898
rect 25589 23840 25594 23896
rect 25650 23840 25820 23896
rect 25589 23838 25820 23840
rect 22185 23835 22251 23838
rect 25589 23835 25655 23838
rect 25814 23836 25820 23838
rect 25884 23836 25890 23900
rect 26182 23836 26188 23900
rect 26252 23898 26299 23900
rect 26252 23896 26344 23898
rect 26294 23840 26344 23896
rect 26252 23838 26344 23840
rect 26252 23836 26299 23838
rect 26233 23835 26299 23836
rect 13556 23702 15394 23762
rect 17033 23762 17099 23765
rect 21265 23764 21331 23765
rect 17033 23760 21098 23762
rect 17033 23704 17038 23760
rect 17094 23704 21098 23760
rect 17033 23702 21098 23704
rect 13556 23700 13562 23702
rect 17033 23699 17099 23702
rect 15653 23626 15719 23629
rect 19609 23626 19675 23629
rect 19926 23626 19932 23628
rect 15653 23624 19932 23626
rect 15653 23568 15658 23624
rect 15714 23568 19614 23624
rect 19670 23568 19932 23624
rect 15653 23566 19932 23568
rect 15653 23563 15719 23566
rect 19609 23563 19675 23566
rect 19926 23564 19932 23566
rect 19996 23564 20002 23628
rect 21038 23626 21098 23702
rect 21214 23700 21220 23764
rect 21284 23762 21331 23764
rect 21541 23762 21607 23765
rect 28349 23762 28415 23765
rect 29200 23762 30000 23792
rect 21284 23760 21376 23762
rect 21326 23704 21376 23760
rect 21284 23702 21376 23704
rect 21541 23760 24870 23762
rect 21541 23704 21546 23760
rect 21602 23704 24870 23760
rect 21541 23702 24870 23704
rect 21284 23700 21331 23702
rect 21265 23699 21331 23700
rect 21541 23699 21607 23702
rect 21173 23626 21239 23629
rect 21038 23624 21239 23626
rect 21038 23568 21178 23624
rect 21234 23568 21239 23624
rect 21038 23566 21239 23568
rect 21173 23563 21239 23566
rect 22001 23626 22067 23629
rect 24393 23626 24459 23629
rect 22001 23624 24459 23626
rect 22001 23568 22006 23624
rect 22062 23568 24398 23624
rect 24454 23568 24459 23624
rect 22001 23566 24459 23568
rect 24810 23626 24870 23702
rect 28349 23760 30000 23762
rect 28349 23704 28354 23760
rect 28410 23704 30000 23760
rect 28349 23702 30000 23704
rect 28349 23699 28415 23702
rect 29200 23672 30000 23702
rect 26877 23626 26943 23629
rect 24810 23624 26943 23626
rect 24810 23568 26882 23624
rect 26938 23568 26943 23624
rect 24810 23566 26943 23568
rect 22001 23563 22067 23566
rect 24393 23563 24459 23566
rect 26877 23563 26943 23566
rect 0 23490 800 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 800 23430
rect 1577 23427 1643 23430
rect 18045 23492 18111 23493
rect 18045 23488 18092 23492
rect 18156 23490 18162 23492
rect 19517 23490 19583 23493
rect 20621 23490 20687 23493
rect 21357 23490 21423 23493
rect 18045 23432 18050 23488
rect 18045 23428 18092 23432
rect 18156 23430 18202 23490
rect 19517 23488 21423 23490
rect 19517 23432 19522 23488
rect 19578 23432 20626 23488
rect 20682 23432 21362 23488
rect 21418 23432 21423 23488
rect 19517 23430 21423 23432
rect 18156 23428 18162 23430
rect 18045 23427 18111 23428
rect 19517 23427 19583 23430
rect 20621 23427 20687 23430
rect 21357 23427 21423 23430
rect 22093 23490 22159 23493
rect 23933 23490 23999 23493
rect 22093 23488 23999 23490
rect 22093 23432 22098 23488
rect 22154 23432 23938 23488
rect 23994 23432 23999 23488
rect 22093 23430 23999 23432
rect 22093 23427 22159 23430
rect 23933 23427 23999 23430
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 19701 23354 19767 23357
rect 20529 23354 20595 23357
rect 19701 23352 20595 23354
rect 19701 23296 19706 23352
rect 19762 23296 20534 23352
rect 20590 23296 20595 23352
rect 19701 23294 20595 23296
rect 19701 23291 19767 23294
rect 20529 23291 20595 23294
rect 20805 23354 20871 23357
rect 23381 23354 23447 23357
rect 24301 23354 24367 23357
rect 20805 23352 24367 23354
rect 20805 23296 20810 23352
rect 20866 23296 23386 23352
rect 23442 23296 24306 23352
rect 24362 23296 24367 23352
rect 20805 23294 24367 23296
rect 20805 23291 20871 23294
rect 23381 23291 23447 23294
rect 24301 23291 24367 23294
rect 17902 23156 17908 23220
rect 17972 23218 17978 23220
rect 27061 23218 27127 23221
rect 17972 23216 27127 23218
rect 17972 23160 27066 23216
rect 27122 23160 27127 23216
rect 17972 23158 27127 23160
rect 17972 23156 17978 23158
rect 27061 23155 27127 23158
rect 12198 23020 12204 23084
rect 12268 23082 12274 23084
rect 19517 23082 19583 23085
rect 21817 23082 21883 23085
rect 26969 23082 27035 23085
rect 12268 23080 19583 23082
rect 12268 23024 19522 23080
rect 19578 23024 19583 23080
rect 12268 23022 19583 23024
rect 12268 23020 12274 23022
rect 19517 23019 19583 23022
rect 19704 23080 27035 23082
rect 19704 23024 21822 23080
rect 21878 23024 26974 23080
rect 27030 23024 27035 23080
rect 19704 23022 27035 23024
rect 17309 22946 17375 22949
rect 17677 22946 17743 22949
rect 19704 22946 19764 23022
rect 21817 23019 21883 23022
rect 26969 23019 27035 23022
rect 28349 23082 28415 23085
rect 29200 23082 30000 23112
rect 28349 23080 30000 23082
rect 28349 23024 28354 23080
rect 28410 23024 30000 23080
rect 28349 23022 30000 23024
rect 28349 23019 28415 23022
rect 29200 22992 30000 23022
rect 17309 22944 19764 22946
rect 17309 22888 17314 22944
rect 17370 22888 17682 22944
rect 17738 22888 19764 22944
rect 17309 22886 19764 22888
rect 23013 22946 23079 22949
rect 26233 22946 26299 22949
rect 23013 22944 26299 22946
rect 23013 22888 23018 22944
rect 23074 22888 26238 22944
rect 26294 22888 26299 22944
rect 23013 22886 26299 22888
rect 17309 22883 17375 22886
rect 17677 22883 17743 22886
rect 23013 22883 23079 22886
rect 26233 22883 26299 22886
rect 7892 22880 8208 22881
rect 0 22720 800 22840
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 18229 22810 18295 22813
rect 19977 22810 20043 22813
rect 20713 22812 20779 22813
rect 18229 22808 20043 22810
rect 18229 22752 18234 22808
rect 18290 22752 19982 22808
rect 20038 22752 20043 22808
rect 18229 22750 20043 22752
rect 18229 22747 18295 22750
rect 19977 22747 20043 22750
rect 20662 22748 20668 22812
rect 20732 22810 20779 22812
rect 22461 22810 22527 22813
rect 20732 22808 20824 22810
rect 20774 22752 20824 22808
rect 20732 22750 20824 22752
rect 22188 22808 22527 22810
rect 22188 22752 22466 22808
rect 22522 22752 22527 22808
rect 22188 22750 22527 22752
rect 20732 22748 20779 22750
rect 20713 22747 20779 22748
rect 22188 22677 22248 22750
rect 22461 22747 22527 22750
rect 23289 22810 23355 22813
rect 23933 22810 23999 22813
rect 23289 22808 23999 22810
rect 23289 22752 23294 22808
rect 23350 22752 23938 22808
rect 23994 22752 23999 22808
rect 23289 22750 23999 22752
rect 23289 22747 23355 22750
rect 23933 22747 23999 22750
rect 25078 22748 25084 22812
rect 25148 22810 25154 22812
rect 25405 22810 25471 22813
rect 25148 22808 25471 22810
rect 25148 22752 25410 22808
rect 25466 22752 25471 22808
rect 25148 22750 25471 22752
rect 25148 22748 25154 22750
rect 25405 22747 25471 22750
rect 25630 22748 25636 22812
rect 25700 22810 25706 22812
rect 25773 22810 25839 22813
rect 25700 22808 25839 22810
rect 25700 22752 25778 22808
rect 25834 22752 25839 22808
rect 25700 22750 25839 22752
rect 25700 22748 25706 22750
rect 25773 22747 25839 22750
rect 12014 22612 12020 22676
rect 12084 22674 12090 22676
rect 21817 22674 21883 22677
rect 12084 22672 21883 22674
rect 12084 22616 21822 22672
rect 21878 22616 21883 22672
rect 12084 22614 21883 22616
rect 12084 22612 12090 22614
rect 21817 22611 21883 22614
rect 22185 22672 22251 22677
rect 22185 22616 22190 22672
rect 22246 22616 22251 22672
rect 22185 22611 22251 22616
rect 23565 22674 23631 22677
rect 25865 22674 25931 22677
rect 23565 22672 25931 22674
rect 23565 22616 23570 22672
rect 23626 22616 25870 22672
rect 25926 22616 25931 22672
rect 23565 22614 25931 22616
rect 23565 22611 23631 22614
rect 25865 22611 25931 22614
rect 17861 22538 17927 22541
rect 23381 22538 23447 22541
rect 17861 22536 23447 22538
rect 17861 22480 17866 22536
rect 17922 22480 23386 22536
rect 23442 22480 23447 22536
rect 17861 22478 23447 22480
rect 17861 22475 17927 22478
rect 23381 22475 23447 22478
rect 22277 22402 22343 22405
rect 24669 22402 24735 22405
rect 22277 22400 24735 22402
rect 22277 22344 22282 22400
rect 22338 22344 24674 22400
rect 24730 22344 24735 22400
rect 22277 22342 24735 22344
rect 22277 22339 22343 22342
rect 24669 22339 24735 22342
rect 28257 22402 28323 22405
rect 29200 22402 30000 22432
rect 28257 22400 30000 22402
rect 28257 22344 28262 22400
rect 28318 22344 30000 22400
rect 28257 22342 30000 22344
rect 28257 22339 28323 22342
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 29200 22312 30000 22342
rect 25257 22271 25573 22272
rect 20161 22266 20227 22269
rect 23197 22266 23263 22269
rect 20161 22264 23263 22266
rect 20161 22208 20166 22264
rect 20222 22208 23202 22264
rect 23258 22208 23263 22264
rect 20161 22206 23263 22208
rect 20161 22203 20227 22206
rect 23197 22203 23263 22206
rect 25865 22266 25931 22269
rect 25998 22266 26004 22268
rect 25865 22264 26004 22266
rect 25865 22208 25870 22264
rect 25926 22208 26004 22264
rect 25865 22206 26004 22208
rect 25865 22203 25931 22206
rect 25998 22204 26004 22206
rect 26068 22204 26074 22268
rect 0 22130 800 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 800 22070
rect 1577 22067 1643 22070
rect 21265 22130 21331 22133
rect 22318 22130 22324 22132
rect 21265 22128 22324 22130
rect 21265 22072 21270 22128
rect 21326 22072 22324 22128
rect 21265 22070 22324 22072
rect 21265 22067 21331 22070
rect 22318 22068 22324 22070
rect 22388 22068 22394 22132
rect 22461 22130 22527 22133
rect 22870 22130 22876 22132
rect 22461 22128 22876 22130
rect 22461 22072 22466 22128
rect 22522 22072 22876 22128
rect 22461 22070 22876 22072
rect 22461 22067 22527 22070
rect 22870 22068 22876 22070
rect 22940 22068 22946 22132
rect 23013 22130 23079 22133
rect 24342 22130 24348 22132
rect 23013 22128 24348 22130
rect 23013 22072 23018 22128
rect 23074 22072 24348 22128
rect 23013 22070 24348 22072
rect 23013 22067 23079 22070
rect 24342 22068 24348 22070
rect 24412 22068 24418 22132
rect 27705 22130 27771 22133
rect 28022 22130 28028 22132
rect 27705 22128 28028 22130
rect 27705 22072 27710 22128
rect 27766 22072 28028 22128
rect 27705 22070 28028 22072
rect 27705 22067 27771 22070
rect 28022 22068 28028 22070
rect 28092 22068 28098 22132
rect 20989 21994 21055 21997
rect 23013 21994 23079 21997
rect 20989 21992 23079 21994
rect 20989 21936 20994 21992
rect 21050 21936 23018 21992
rect 23074 21936 23079 21992
rect 20989 21934 23079 21936
rect 20989 21931 21055 21934
rect 23013 21931 23079 21934
rect 23381 21994 23447 21997
rect 23606 21994 23612 21996
rect 23381 21992 23612 21994
rect 23381 21936 23386 21992
rect 23442 21936 23612 21992
rect 23381 21934 23612 21936
rect 23381 21931 23447 21934
rect 23606 21932 23612 21934
rect 23676 21932 23682 21996
rect 19425 21858 19491 21861
rect 20805 21858 20871 21861
rect 19425 21856 20871 21858
rect 19425 21800 19430 21856
rect 19486 21800 20810 21856
rect 20866 21800 20871 21856
rect 19425 21798 20871 21800
rect 19425 21795 19491 21798
rect 20805 21795 20871 21798
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 28730 21727 29046 21728
rect 17166 21660 17172 21724
rect 17236 21722 17242 21724
rect 17236 21662 20730 21722
rect 17236 21660 17242 21662
rect 20294 21524 20300 21588
rect 20364 21586 20370 21588
rect 20529 21586 20595 21589
rect 20364 21584 20595 21586
rect 20364 21528 20534 21584
rect 20590 21528 20595 21584
rect 20364 21526 20595 21528
rect 20670 21586 20730 21662
rect 23054 21660 23060 21724
rect 23124 21722 23130 21724
rect 23289 21722 23355 21725
rect 23124 21720 23355 21722
rect 23124 21664 23294 21720
rect 23350 21664 23355 21720
rect 29200 21688 30000 21752
rect 23124 21662 23355 21664
rect 23124 21660 23130 21662
rect 23289 21659 23355 21662
rect 29134 21632 30000 21688
rect 29134 21628 29378 21632
rect 22461 21586 22527 21589
rect 20670 21584 22527 21586
rect 20670 21528 22466 21584
rect 22522 21528 22527 21584
rect 20670 21526 22527 21528
rect 20364 21524 20370 21526
rect 20529 21523 20595 21526
rect 22461 21523 22527 21526
rect 28349 21586 28415 21589
rect 29134 21586 29194 21628
rect 28349 21584 29194 21586
rect 28349 21528 28354 21584
rect 28410 21528 29194 21584
rect 28349 21526 29194 21528
rect 28349 21523 28415 21526
rect 0 21450 800 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 800 21390
rect 1577 21387 1643 21390
rect 24853 21450 24919 21453
rect 25814 21450 25820 21452
rect 24853 21448 25820 21450
rect 24853 21392 24858 21448
rect 24914 21392 25820 21448
rect 24853 21390 25820 21392
rect 24853 21387 24919 21390
rect 25814 21388 25820 21390
rect 25884 21388 25890 21452
rect 21173 21314 21239 21317
rect 22645 21314 22711 21317
rect 21173 21312 22711 21314
rect 21173 21256 21178 21312
rect 21234 21256 22650 21312
rect 22706 21256 22711 21312
rect 21173 21254 22711 21256
rect 21173 21251 21239 21254
rect 22645 21251 22711 21254
rect 23749 21314 23815 21317
rect 23974 21314 23980 21316
rect 23749 21312 23980 21314
rect 23749 21256 23754 21312
rect 23810 21256 23980 21312
rect 23749 21254 23980 21256
rect 23749 21251 23815 21254
rect 23974 21252 23980 21254
rect 24044 21252 24050 21316
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 28349 21042 28415 21045
rect 29200 21042 30000 21072
rect 28349 21040 30000 21042
rect 28349 20984 28354 21040
rect 28410 20984 30000 21040
rect 28349 20982 30000 20984
rect 28349 20979 28415 20982
rect 29200 20952 30000 20982
rect 0 20680 800 20800
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 19977 20634 20043 20637
rect 20110 20634 20116 20636
rect 19977 20632 20116 20634
rect 19977 20576 19982 20632
rect 20038 20576 20116 20632
rect 19977 20574 20116 20576
rect 19977 20571 20043 20574
rect 20110 20572 20116 20574
rect 20180 20572 20186 20636
rect 24894 20300 24900 20364
rect 24964 20362 24970 20364
rect 25589 20362 25655 20365
rect 24964 20360 25655 20362
rect 24964 20304 25594 20360
rect 25650 20304 25655 20360
rect 24964 20302 25655 20304
rect 24964 20300 24970 20302
rect 25589 20299 25655 20302
rect 28349 20362 28415 20365
rect 29200 20362 30000 20392
rect 28349 20360 30000 20362
rect 28349 20304 28354 20360
rect 28410 20304 30000 20360
rect 28349 20302 30000 20304
rect 28349 20299 28415 20302
rect 29200 20272 30000 20302
rect 4419 20160 4735 20161
rect 0 20090 800 20120
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 28349 19818 28415 19821
rect 28349 19816 29194 19818
rect 28349 19760 28354 19816
rect 28410 19760 29194 19816
rect 28349 19758 29194 19760
rect 28349 19755 28415 19758
rect 29134 19716 29194 19758
rect 29134 19712 29378 19716
rect 29134 19656 30000 19712
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 29200 19592 30000 19656
rect 28730 19551 29046 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 28349 19002 28415 19005
rect 29200 19002 30000 19032
rect 28349 19000 30000 19002
rect 28349 18944 28354 19000
rect 28410 18944 30000 19000
rect 28349 18942 30000 18944
rect 28349 18939 28415 18942
rect 29200 18912 30000 18942
rect 0 18640 800 18760
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 28730 18463 29046 18464
rect 28349 18322 28415 18325
rect 29200 18322 30000 18352
rect 28349 18320 30000 18322
rect 28349 18264 28354 18320
rect 28410 18264 30000 18320
rect 28349 18262 30000 18264
rect 28349 18259 28415 18262
rect 29200 18232 30000 18262
rect 0 18050 800 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 800 17990
rect 1577 17987 1643 17990
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 28349 17642 28415 17645
rect 29200 17642 30000 17672
rect 28349 17640 30000 17642
rect 28349 17584 28354 17640
rect 28410 17584 30000 17640
rect 28349 17582 30000 17584
rect 28349 17579 28415 17582
rect 29200 17552 30000 17582
rect 7892 17440 8208 17441
rect 0 17370 800 17400
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 28349 16962 28415 16965
rect 29200 16962 30000 16992
rect 28349 16960 30000 16962
rect 28349 16904 28354 16960
rect 28410 16904 30000 16960
rect 28349 16902 30000 16904
rect 28349 16899 28415 16902
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 29200 16872 30000 16902
rect 25257 16831 25573 16832
rect 0 16600 800 16720
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 29200 16192 30000 16312
rect 0 16010 800 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 800 15950
rect 1577 15947 1643 15950
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 28349 15602 28415 15605
rect 29200 15602 30000 15632
rect 28349 15600 30000 15602
rect 28349 15544 28354 15600
rect 28410 15544 30000 15600
rect 28349 15542 30000 15544
rect 28349 15539 28415 15542
rect 29200 15512 30000 15542
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 28730 15199 29046 15200
rect 28349 14922 28415 14925
rect 29200 14922 30000 14952
rect 28349 14920 30000 14922
rect 28349 14864 28354 14920
rect 28410 14864 30000 14920
rect 28349 14862 30000 14864
rect 28349 14859 28415 14862
rect 29200 14832 30000 14862
rect 4419 14720 4735 14721
rect 0 14560 800 14680
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 29200 14152 30000 14272
rect 28730 14111 29046 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 28349 13562 28415 13565
rect 29200 13562 30000 13592
rect 28349 13560 30000 13562
rect 28349 13504 28354 13560
rect 28410 13504 30000 13560
rect 28349 13502 30000 13504
rect 28349 13499 28415 13502
rect 29200 13472 30000 13502
rect 0 13290 800 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 800 13230
rect 1577 13227 1643 13230
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 28349 12882 28415 12885
rect 29200 12882 30000 12912
rect 28349 12880 30000 12882
rect 28349 12824 28354 12880
rect 28410 12824 30000 12880
rect 28349 12822 30000 12824
rect 28349 12819 28415 12822
rect 29200 12792 30000 12822
rect 0 12520 800 12640
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 29200 12112 30000 12232
rect 7892 12000 8208 12001
rect 0 11930 800 11960
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 28730 11935 29046 11936
rect 1577 11930 1643 11933
rect 0 11928 1643 11930
rect 0 11872 1582 11928
rect 1638 11872 1643 11928
rect 0 11870 1643 11872
rect 0 11840 800 11870
rect 1577 11867 1643 11870
rect 28349 11522 28415 11525
rect 29200 11522 30000 11552
rect 28349 11520 30000 11522
rect 28349 11464 28354 11520
rect 28410 11464 30000 11520
rect 28349 11462 30000 11464
rect 28349 11459 28415 11462
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 29200 11432 30000 11462
rect 25257 11391 25573 11392
rect 0 11250 800 11280
rect 1577 11250 1643 11253
rect 0 11248 1643 11250
rect 0 11192 1582 11248
rect 1638 11192 1643 11248
rect 0 11190 1643 11192
rect 0 11160 800 11190
rect 1577 11187 1643 11190
rect 28349 11114 28415 11117
rect 28349 11112 29378 11114
rect 28349 11056 28354 11112
rect 28410 11056 29378 11112
rect 28349 11054 29378 11056
rect 28349 11051 28415 11054
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 29318 10872 29378 11054
rect 28730 10847 29046 10848
rect 29200 10752 30000 10872
rect 0 10480 800 10600
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 29200 10072 30000 10192
rect 0 9890 800 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 800 9830
rect 1577 9827 1643 9830
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 28349 9482 28415 9485
rect 29200 9482 30000 9512
rect 28349 9480 30000 9482
rect 28349 9424 28354 9480
rect 28410 9424 30000 9480
rect 28349 9422 30000 9424
rect 28349 9419 28415 9422
rect 29200 9392 30000 9422
rect 4419 9280 4735 9281
rect 0 9210 800 9240
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 1577 9210 1643 9213
rect 0 9208 1643 9210
rect 0 9152 1582 9208
rect 1638 9152 1643 9208
rect 0 9150 1643 9152
rect 0 9120 800 9150
rect 1577 9147 1643 9150
rect 28349 9074 28415 9077
rect 28349 9072 29378 9074
rect 28349 9016 28354 9072
rect 28410 9016 29378 9072
rect 28349 9014 29378 9016
rect 28349 9011 28415 9014
rect 29318 8832 29378 9014
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 29200 8712 30000 8832
rect 28730 8671 29046 8672
rect 0 8440 800 8560
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 29200 8032 30000 8152
rect 0 7850 800 7880
rect 1577 7850 1643 7853
rect 0 7848 1643 7850
rect 0 7792 1582 7848
rect 1638 7792 1643 7848
rect 0 7790 1643 7792
rect 0 7760 800 7790
rect 1577 7787 1643 7790
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 28349 7442 28415 7445
rect 29200 7442 30000 7472
rect 28349 7440 30000 7442
rect 28349 7384 28354 7440
rect 28410 7384 30000 7440
rect 28349 7382 30000 7384
rect 28349 7379 28415 7382
rect 29200 7352 30000 7382
rect 0 7170 800 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 800 7110
rect 1577 7107 1643 7110
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 28349 6762 28415 6765
rect 29200 6762 30000 6792
rect 28349 6760 30000 6762
rect 28349 6704 28354 6760
rect 28410 6704 30000 6760
rect 28349 6702 30000 6704
rect 28349 6699 28415 6702
rect 29200 6672 30000 6702
rect 7892 6560 8208 6561
rect 0 6400 800 6520
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 29200 5992 30000 6112
rect 25257 5951 25573 5952
rect 0 5810 800 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 800 5750
rect 1577 5747 1643 5750
rect 28349 5674 28415 5677
rect 28349 5672 29378 5674
rect 28349 5616 28354 5672
rect 28410 5616 29378 5672
rect 28349 5614 29378 5616
rect 28349 5611 28415 5614
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 29318 5432 29378 5614
rect 28730 5407 29046 5408
rect 29200 5312 30000 5432
rect 0 5130 800 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 800 5070
rect 1577 5067 1643 5070
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 28349 4722 28415 4725
rect 29200 4722 30000 4752
rect 28349 4720 30000 4722
rect 28349 4664 28354 4720
rect 28410 4664 30000 4720
rect 28349 4662 30000 4664
rect 28349 4659 28415 4662
rect 29200 4632 30000 4662
rect 0 4360 800 4480
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 29200 3952 30000 4072
rect 4419 3840 4735 3841
rect 0 3770 800 3800
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 28349 3634 28415 3637
rect 28349 3632 29378 3634
rect 28349 3576 28354 3632
rect 28410 3576 29378 3632
rect 28349 3574 29378 3576
rect 28349 3571 28415 3574
rect 29318 3392 29378 3574
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 29200 3272 30000 3392
rect 28730 3231 29046 3232
rect 0 3090 800 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 800 3030
rect 1577 3027 1643 3030
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 28349 2682 28415 2685
rect 29200 2682 30000 2712
rect 28349 2680 30000 2682
rect 28349 2624 28354 2680
rect 28410 2624 30000 2680
rect 28349 2622 30000 2624
rect 28349 2619 28415 2622
rect 29200 2592 30000 2622
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 28730 2143 29046 2144
rect 29200 1912 30000 2032
<< via3 >>
rect 26004 31860 26068 31924
rect 23244 31724 23308 31788
rect 7898 31580 7962 31584
rect 7898 31524 7902 31580
rect 7902 31524 7958 31580
rect 7958 31524 7962 31580
rect 7898 31520 7962 31524
rect 7978 31580 8042 31584
rect 7978 31524 7982 31580
rect 7982 31524 8038 31580
rect 8038 31524 8042 31580
rect 7978 31520 8042 31524
rect 8058 31580 8122 31584
rect 8058 31524 8062 31580
rect 8062 31524 8118 31580
rect 8118 31524 8122 31580
rect 8058 31520 8122 31524
rect 8138 31580 8202 31584
rect 8138 31524 8142 31580
rect 8142 31524 8198 31580
rect 8198 31524 8202 31580
rect 8138 31520 8202 31524
rect 14844 31580 14908 31584
rect 14844 31524 14848 31580
rect 14848 31524 14904 31580
rect 14904 31524 14908 31580
rect 14844 31520 14908 31524
rect 14924 31580 14988 31584
rect 14924 31524 14928 31580
rect 14928 31524 14984 31580
rect 14984 31524 14988 31580
rect 14924 31520 14988 31524
rect 15004 31580 15068 31584
rect 15004 31524 15008 31580
rect 15008 31524 15064 31580
rect 15064 31524 15068 31580
rect 15004 31520 15068 31524
rect 15084 31580 15148 31584
rect 15084 31524 15088 31580
rect 15088 31524 15144 31580
rect 15144 31524 15148 31580
rect 15084 31520 15148 31524
rect 21790 31580 21854 31584
rect 21790 31524 21794 31580
rect 21794 31524 21850 31580
rect 21850 31524 21854 31580
rect 21790 31520 21854 31524
rect 21870 31580 21934 31584
rect 21870 31524 21874 31580
rect 21874 31524 21930 31580
rect 21930 31524 21934 31580
rect 21870 31520 21934 31524
rect 21950 31580 22014 31584
rect 21950 31524 21954 31580
rect 21954 31524 22010 31580
rect 22010 31524 22014 31580
rect 21950 31520 22014 31524
rect 22030 31580 22094 31584
rect 22030 31524 22034 31580
rect 22034 31524 22090 31580
rect 22090 31524 22094 31580
rect 22030 31520 22094 31524
rect 28736 31580 28800 31584
rect 28736 31524 28740 31580
rect 28740 31524 28796 31580
rect 28796 31524 28800 31580
rect 28736 31520 28800 31524
rect 28816 31580 28880 31584
rect 28816 31524 28820 31580
rect 28820 31524 28876 31580
rect 28876 31524 28880 31580
rect 28816 31520 28880 31524
rect 28896 31580 28960 31584
rect 28896 31524 28900 31580
rect 28900 31524 28956 31580
rect 28956 31524 28960 31580
rect 28896 31520 28960 31524
rect 28976 31580 29040 31584
rect 28976 31524 28980 31580
rect 28980 31524 29036 31580
rect 29036 31524 29040 31580
rect 28976 31520 29040 31524
rect 21220 31452 21284 31516
rect 18828 31044 18892 31108
rect 4425 31036 4489 31040
rect 4425 30980 4429 31036
rect 4429 30980 4485 31036
rect 4485 30980 4489 31036
rect 4425 30976 4489 30980
rect 4505 31036 4569 31040
rect 4505 30980 4509 31036
rect 4509 30980 4565 31036
rect 4565 30980 4569 31036
rect 4505 30976 4569 30980
rect 4585 31036 4649 31040
rect 4585 30980 4589 31036
rect 4589 30980 4645 31036
rect 4645 30980 4649 31036
rect 4585 30976 4649 30980
rect 4665 31036 4729 31040
rect 4665 30980 4669 31036
rect 4669 30980 4725 31036
rect 4725 30980 4729 31036
rect 4665 30976 4729 30980
rect 11371 31036 11435 31040
rect 11371 30980 11375 31036
rect 11375 30980 11431 31036
rect 11431 30980 11435 31036
rect 11371 30976 11435 30980
rect 11451 31036 11515 31040
rect 11451 30980 11455 31036
rect 11455 30980 11511 31036
rect 11511 30980 11515 31036
rect 11451 30976 11515 30980
rect 11531 31036 11595 31040
rect 11531 30980 11535 31036
rect 11535 30980 11591 31036
rect 11591 30980 11595 31036
rect 11531 30976 11595 30980
rect 11611 31036 11675 31040
rect 11611 30980 11615 31036
rect 11615 30980 11671 31036
rect 11671 30980 11675 31036
rect 11611 30976 11675 30980
rect 18317 31036 18381 31040
rect 18317 30980 18321 31036
rect 18321 30980 18377 31036
rect 18377 30980 18381 31036
rect 18317 30976 18381 30980
rect 18397 31036 18461 31040
rect 18397 30980 18401 31036
rect 18401 30980 18457 31036
rect 18457 30980 18461 31036
rect 18397 30976 18461 30980
rect 18477 31036 18541 31040
rect 18477 30980 18481 31036
rect 18481 30980 18537 31036
rect 18537 30980 18541 31036
rect 18477 30976 18541 30980
rect 18557 31036 18621 31040
rect 18557 30980 18561 31036
rect 18561 30980 18617 31036
rect 18617 30980 18621 31036
rect 18557 30976 18621 30980
rect 25263 31036 25327 31040
rect 25263 30980 25267 31036
rect 25267 30980 25323 31036
rect 25323 30980 25327 31036
rect 25263 30976 25327 30980
rect 25343 31036 25407 31040
rect 25343 30980 25347 31036
rect 25347 30980 25403 31036
rect 25403 30980 25407 31036
rect 25343 30976 25407 30980
rect 25423 31036 25487 31040
rect 25423 30980 25427 31036
rect 25427 30980 25483 31036
rect 25483 30980 25487 31036
rect 25423 30976 25487 30980
rect 25503 31036 25567 31040
rect 25503 30980 25507 31036
rect 25507 30980 25563 31036
rect 25563 30980 25567 31036
rect 25503 30976 25567 30980
rect 23428 30908 23492 30972
rect 17356 30636 17420 30700
rect 17908 30636 17972 30700
rect 23060 30636 23124 30700
rect 19932 30500 19996 30564
rect 7898 30492 7962 30496
rect 7898 30436 7902 30492
rect 7902 30436 7958 30492
rect 7958 30436 7962 30492
rect 7898 30432 7962 30436
rect 7978 30492 8042 30496
rect 7978 30436 7982 30492
rect 7982 30436 8038 30492
rect 8038 30436 8042 30492
rect 7978 30432 8042 30436
rect 8058 30492 8122 30496
rect 8058 30436 8062 30492
rect 8062 30436 8118 30492
rect 8118 30436 8122 30492
rect 8058 30432 8122 30436
rect 8138 30492 8202 30496
rect 8138 30436 8142 30492
rect 8142 30436 8198 30492
rect 8198 30436 8202 30492
rect 8138 30432 8202 30436
rect 14844 30492 14908 30496
rect 14844 30436 14848 30492
rect 14848 30436 14904 30492
rect 14904 30436 14908 30492
rect 14844 30432 14908 30436
rect 14924 30492 14988 30496
rect 14924 30436 14928 30492
rect 14928 30436 14984 30492
rect 14984 30436 14988 30492
rect 14924 30432 14988 30436
rect 15004 30492 15068 30496
rect 15004 30436 15008 30492
rect 15008 30436 15064 30492
rect 15064 30436 15068 30492
rect 15004 30432 15068 30436
rect 15084 30492 15148 30496
rect 15084 30436 15088 30492
rect 15088 30436 15144 30492
rect 15144 30436 15148 30492
rect 15084 30432 15148 30436
rect 21790 30492 21854 30496
rect 21790 30436 21794 30492
rect 21794 30436 21850 30492
rect 21850 30436 21854 30492
rect 21790 30432 21854 30436
rect 21870 30492 21934 30496
rect 21870 30436 21874 30492
rect 21874 30436 21930 30492
rect 21930 30436 21934 30492
rect 21870 30432 21934 30436
rect 21950 30492 22014 30496
rect 21950 30436 21954 30492
rect 21954 30436 22010 30492
rect 22010 30436 22014 30492
rect 21950 30432 22014 30436
rect 22030 30492 22094 30496
rect 22030 30436 22034 30492
rect 22034 30436 22090 30492
rect 22090 30436 22094 30492
rect 22030 30432 22094 30436
rect 28736 30492 28800 30496
rect 28736 30436 28740 30492
rect 28740 30436 28796 30492
rect 28796 30436 28800 30492
rect 28736 30432 28800 30436
rect 28816 30492 28880 30496
rect 28816 30436 28820 30492
rect 28820 30436 28876 30492
rect 28876 30436 28880 30492
rect 28816 30432 28880 30436
rect 28896 30492 28960 30496
rect 28896 30436 28900 30492
rect 28900 30436 28956 30492
rect 28956 30436 28960 30492
rect 28896 30432 28960 30436
rect 28976 30492 29040 30496
rect 28976 30436 28980 30492
rect 28980 30436 29036 30492
rect 29036 30436 29040 30492
rect 28976 30432 29040 30436
rect 12020 30364 12084 30428
rect 20484 30364 20548 30428
rect 15332 30288 15396 30292
rect 15332 30232 15346 30288
rect 15346 30232 15396 30288
rect 15332 30228 15396 30232
rect 9996 30092 10060 30156
rect 19196 30152 19260 30156
rect 19196 30096 19210 30152
rect 19210 30096 19260 30152
rect 16804 29956 16868 30020
rect 19196 30092 19260 30096
rect 20668 29956 20732 30020
rect 25084 30016 25148 30020
rect 25084 29960 25098 30016
rect 25098 29960 25148 30016
rect 4425 29948 4489 29952
rect 4425 29892 4429 29948
rect 4429 29892 4485 29948
rect 4485 29892 4489 29948
rect 4425 29888 4489 29892
rect 4505 29948 4569 29952
rect 4505 29892 4509 29948
rect 4509 29892 4565 29948
rect 4565 29892 4569 29948
rect 4505 29888 4569 29892
rect 4585 29948 4649 29952
rect 4585 29892 4589 29948
rect 4589 29892 4645 29948
rect 4645 29892 4649 29948
rect 4585 29888 4649 29892
rect 4665 29948 4729 29952
rect 4665 29892 4669 29948
rect 4669 29892 4725 29948
rect 4725 29892 4729 29948
rect 4665 29888 4729 29892
rect 11371 29948 11435 29952
rect 11371 29892 11375 29948
rect 11375 29892 11431 29948
rect 11431 29892 11435 29948
rect 11371 29888 11435 29892
rect 11451 29948 11515 29952
rect 11451 29892 11455 29948
rect 11455 29892 11511 29948
rect 11511 29892 11515 29948
rect 11451 29888 11515 29892
rect 11531 29948 11595 29952
rect 11531 29892 11535 29948
rect 11535 29892 11591 29948
rect 11591 29892 11595 29948
rect 11531 29888 11595 29892
rect 11611 29948 11675 29952
rect 11611 29892 11615 29948
rect 11615 29892 11671 29948
rect 11671 29892 11675 29948
rect 11611 29888 11675 29892
rect 18317 29948 18381 29952
rect 18317 29892 18321 29948
rect 18321 29892 18377 29948
rect 18377 29892 18381 29948
rect 18317 29888 18381 29892
rect 18397 29948 18461 29952
rect 18397 29892 18401 29948
rect 18401 29892 18457 29948
rect 18457 29892 18461 29948
rect 18397 29888 18461 29892
rect 18477 29948 18541 29952
rect 18477 29892 18481 29948
rect 18481 29892 18537 29948
rect 18537 29892 18541 29948
rect 18477 29888 18541 29892
rect 18557 29948 18621 29952
rect 18557 29892 18561 29948
rect 18561 29892 18617 29948
rect 18617 29892 18621 29948
rect 18557 29888 18621 29892
rect 18092 29880 18156 29884
rect 25084 29956 25148 29960
rect 25263 29948 25327 29952
rect 25263 29892 25267 29948
rect 25267 29892 25323 29948
rect 25323 29892 25327 29948
rect 25263 29888 25327 29892
rect 25343 29948 25407 29952
rect 25343 29892 25347 29948
rect 25347 29892 25403 29948
rect 25403 29892 25407 29948
rect 25343 29888 25407 29892
rect 25423 29948 25487 29952
rect 25423 29892 25427 29948
rect 25427 29892 25483 29948
rect 25483 29892 25487 29948
rect 25423 29888 25487 29892
rect 25503 29948 25567 29952
rect 25503 29892 25507 29948
rect 25507 29892 25563 29948
rect 25563 29892 25567 29948
rect 25503 29888 25567 29892
rect 18092 29824 18106 29880
rect 18106 29824 18156 29880
rect 18092 29820 18156 29824
rect 20852 29684 20916 29748
rect 19380 29548 19444 29612
rect 15884 29412 15948 29476
rect 18092 29412 18156 29476
rect 7898 29404 7962 29408
rect 7898 29348 7902 29404
rect 7902 29348 7958 29404
rect 7958 29348 7962 29404
rect 7898 29344 7962 29348
rect 7978 29404 8042 29408
rect 7978 29348 7982 29404
rect 7982 29348 8038 29404
rect 8038 29348 8042 29404
rect 7978 29344 8042 29348
rect 8058 29404 8122 29408
rect 8058 29348 8062 29404
rect 8062 29348 8118 29404
rect 8118 29348 8122 29404
rect 8058 29344 8122 29348
rect 8138 29404 8202 29408
rect 8138 29348 8142 29404
rect 8142 29348 8198 29404
rect 8198 29348 8202 29404
rect 8138 29344 8202 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 21790 29404 21854 29408
rect 21790 29348 21794 29404
rect 21794 29348 21850 29404
rect 21850 29348 21854 29404
rect 21790 29344 21854 29348
rect 21870 29404 21934 29408
rect 21870 29348 21874 29404
rect 21874 29348 21930 29404
rect 21930 29348 21934 29404
rect 21870 29344 21934 29348
rect 21950 29404 22014 29408
rect 21950 29348 21954 29404
rect 21954 29348 22010 29404
rect 22010 29348 22014 29404
rect 21950 29344 22014 29348
rect 22030 29404 22094 29408
rect 22030 29348 22034 29404
rect 22034 29348 22090 29404
rect 22090 29348 22094 29404
rect 22030 29344 22094 29348
rect 28736 29404 28800 29408
rect 28736 29348 28740 29404
rect 28740 29348 28796 29404
rect 28796 29348 28800 29404
rect 28736 29344 28800 29348
rect 28816 29404 28880 29408
rect 28816 29348 28820 29404
rect 28820 29348 28876 29404
rect 28876 29348 28880 29404
rect 28816 29344 28880 29348
rect 28896 29404 28960 29408
rect 28896 29348 28900 29404
rect 28900 29348 28956 29404
rect 28956 29348 28960 29404
rect 28896 29344 28960 29348
rect 28976 29404 29040 29408
rect 28976 29348 28980 29404
rect 28980 29348 29036 29404
rect 29036 29348 29040 29404
rect 28976 29344 29040 29348
rect 16620 29276 16684 29340
rect 17724 29276 17788 29340
rect 18828 29276 18892 29340
rect 9996 29004 10060 29068
rect 10916 29004 10980 29068
rect 12204 29004 12268 29068
rect 14596 29004 14660 29068
rect 17172 29004 17236 29068
rect 17356 29064 17420 29068
rect 17356 29008 17406 29064
rect 17406 29008 17420 29064
rect 17356 29004 17420 29008
rect 14412 28868 14476 28932
rect 22876 28868 22940 28932
rect 4425 28860 4489 28864
rect 4425 28804 4429 28860
rect 4429 28804 4485 28860
rect 4485 28804 4489 28860
rect 4425 28800 4489 28804
rect 4505 28860 4569 28864
rect 4505 28804 4509 28860
rect 4509 28804 4565 28860
rect 4565 28804 4569 28860
rect 4505 28800 4569 28804
rect 4585 28860 4649 28864
rect 4585 28804 4589 28860
rect 4589 28804 4645 28860
rect 4645 28804 4649 28860
rect 4585 28800 4649 28804
rect 4665 28860 4729 28864
rect 4665 28804 4669 28860
rect 4669 28804 4725 28860
rect 4725 28804 4729 28860
rect 4665 28800 4729 28804
rect 11371 28860 11435 28864
rect 11371 28804 11375 28860
rect 11375 28804 11431 28860
rect 11431 28804 11435 28860
rect 11371 28800 11435 28804
rect 11451 28860 11515 28864
rect 11451 28804 11455 28860
rect 11455 28804 11511 28860
rect 11511 28804 11515 28860
rect 11451 28800 11515 28804
rect 11531 28860 11595 28864
rect 11531 28804 11535 28860
rect 11535 28804 11591 28860
rect 11591 28804 11595 28860
rect 11531 28800 11595 28804
rect 11611 28860 11675 28864
rect 11611 28804 11615 28860
rect 11615 28804 11671 28860
rect 11671 28804 11675 28860
rect 11611 28800 11675 28804
rect 18317 28860 18381 28864
rect 18317 28804 18321 28860
rect 18321 28804 18377 28860
rect 18377 28804 18381 28860
rect 18317 28800 18381 28804
rect 18397 28860 18461 28864
rect 18397 28804 18401 28860
rect 18401 28804 18457 28860
rect 18457 28804 18461 28860
rect 18397 28800 18461 28804
rect 18477 28860 18541 28864
rect 18477 28804 18481 28860
rect 18481 28804 18537 28860
rect 18537 28804 18541 28860
rect 18477 28800 18541 28804
rect 18557 28860 18621 28864
rect 18557 28804 18561 28860
rect 18561 28804 18617 28860
rect 18617 28804 18621 28860
rect 18557 28800 18621 28804
rect 25263 28860 25327 28864
rect 25263 28804 25267 28860
rect 25267 28804 25323 28860
rect 25323 28804 25327 28860
rect 25263 28800 25327 28804
rect 25343 28860 25407 28864
rect 25343 28804 25347 28860
rect 25347 28804 25403 28860
rect 25403 28804 25407 28860
rect 25343 28800 25407 28804
rect 25423 28860 25487 28864
rect 25423 28804 25427 28860
rect 25427 28804 25483 28860
rect 25483 28804 25487 28860
rect 25423 28800 25487 28804
rect 25503 28860 25567 28864
rect 25503 28804 25507 28860
rect 25507 28804 25563 28860
rect 25563 28804 25567 28860
rect 25503 28800 25567 28804
rect 23796 28596 23860 28660
rect 24716 28460 24780 28524
rect 25820 28460 25884 28524
rect 27476 28324 27540 28388
rect 7898 28316 7962 28320
rect 7898 28260 7902 28316
rect 7902 28260 7958 28316
rect 7958 28260 7962 28316
rect 7898 28256 7962 28260
rect 7978 28316 8042 28320
rect 7978 28260 7982 28316
rect 7982 28260 8038 28316
rect 8038 28260 8042 28316
rect 7978 28256 8042 28260
rect 8058 28316 8122 28320
rect 8058 28260 8062 28316
rect 8062 28260 8118 28316
rect 8118 28260 8122 28316
rect 8058 28256 8122 28260
rect 8138 28316 8202 28320
rect 8138 28260 8142 28316
rect 8142 28260 8198 28316
rect 8198 28260 8202 28316
rect 8138 28256 8202 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 21790 28316 21854 28320
rect 21790 28260 21794 28316
rect 21794 28260 21850 28316
rect 21850 28260 21854 28316
rect 21790 28256 21854 28260
rect 21870 28316 21934 28320
rect 21870 28260 21874 28316
rect 21874 28260 21930 28316
rect 21930 28260 21934 28316
rect 21870 28256 21934 28260
rect 21950 28316 22014 28320
rect 21950 28260 21954 28316
rect 21954 28260 22010 28316
rect 22010 28260 22014 28316
rect 21950 28256 22014 28260
rect 22030 28316 22094 28320
rect 22030 28260 22034 28316
rect 22034 28260 22090 28316
rect 22090 28260 22094 28316
rect 22030 28256 22094 28260
rect 28736 28316 28800 28320
rect 28736 28260 28740 28316
rect 28740 28260 28796 28316
rect 28796 28260 28800 28316
rect 28736 28256 28800 28260
rect 28816 28316 28880 28320
rect 28816 28260 28820 28316
rect 28820 28260 28876 28316
rect 28876 28260 28880 28316
rect 28816 28256 28880 28260
rect 28896 28316 28960 28320
rect 28896 28260 28900 28316
rect 28900 28260 28956 28316
rect 28956 28260 28960 28316
rect 28896 28256 28960 28260
rect 28976 28316 29040 28320
rect 28976 28260 28980 28316
rect 28980 28260 29036 28316
rect 29036 28260 29040 28316
rect 28976 28256 29040 28260
rect 15516 28188 15580 28252
rect 24532 28188 24596 28252
rect 17540 27780 17604 27844
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 15332 27644 15396 27708
rect 17908 27644 17972 27708
rect 20300 27644 20364 27708
rect 23612 27644 23676 27708
rect 20668 27508 20732 27572
rect 23428 27508 23492 27572
rect 26188 27916 26252 27980
rect 27476 27916 27540 27980
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 13492 27236 13556 27300
rect 14412 27296 14476 27300
rect 14412 27240 14462 27296
rect 14462 27240 14476 27296
rect 14412 27236 14476 27240
rect 15516 27236 15580 27300
rect 16068 27296 16132 27300
rect 16068 27240 16082 27296
rect 16082 27240 16132 27296
rect 16068 27236 16132 27240
rect 16620 27236 16684 27300
rect 22692 27236 22756 27300
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 15884 27100 15948 27164
rect 22324 27100 22388 27164
rect 24900 27100 24964 27164
rect 24716 26964 24780 27028
rect 25084 26828 25148 26892
rect 25636 26828 25700 26892
rect 19196 26752 19260 26756
rect 19196 26696 19246 26752
rect 19246 26696 19260 26752
rect 19196 26692 19260 26696
rect 20668 26752 20732 26756
rect 20668 26696 20718 26752
rect 20718 26696 20732 26752
rect 20668 26692 20732 26696
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 20852 26420 20916 26484
rect 24348 26420 24412 26484
rect 28028 26420 28092 26484
rect 16620 26284 16684 26348
rect 16068 26208 16132 26212
rect 16068 26152 16118 26208
rect 16118 26152 16132 26208
rect 16068 26148 16132 26152
rect 23796 26148 23860 26212
rect 23980 26148 24044 26212
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 17540 26012 17604 26076
rect 19380 26012 19444 26076
rect 19748 26012 19812 26076
rect 23060 26012 23124 26076
rect 25084 26012 25148 26076
rect 26372 26012 26436 26076
rect 10916 25740 10980 25804
rect 19932 25876 19996 25940
rect 20484 25876 20548 25940
rect 25084 25604 25148 25668
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 26004 25468 26068 25532
rect 14596 25332 14660 25396
rect 25820 25332 25884 25396
rect 26188 25332 26252 25396
rect 19932 25120 19996 25124
rect 19932 25064 19982 25120
rect 19982 25064 19996 25120
rect 19932 25060 19996 25064
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 16620 24924 16684 24988
rect 23244 24984 23308 24988
rect 23244 24928 23294 24984
rect 23294 24928 23308 24984
rect 23244 24924 23308 24928
rect 18828 24788 18892 24852
rect 24532 24788 24596 24852
rect 26004 24788 26068 24852
rect 17724 24652 17788 24716
rect 25084 24652 25148 24716
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 19748 24516 19812 24580
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 27476 24304 27540 24308
rect 27476 24248 27526 24304
rect 27526 24248 27540 24304
rect 27476 24244 27540 24248
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 13492 23700 13556 23764
rect 20116 23836 20180 23900
rect 22692 23972 22756 24036
rect 25084 24032 25148 24036
rect 25084 23976 25134 24032
rect 25134 23976 25148 24032
rect 25084 23972 25148 23976
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 26372 23972 26436 24036
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 25820 23836 25884 23900
rect 26188 23896 26252 23900
rect 26188 23840 26238 23896
rect 26238 23840 26252 23896
rect 26188 23836 26252 23840
rect 19932 23564 19996 23628
rect 21220 23760 21284 23764
rect 21220 23704 21270 23760
rect 21270 23704 21284 23760
rect 21220 23700 21284 23704
rect 18092 23488 18156 23492
rect 18092 23432 18106 23488
rect 18106 23432 18156 23488
rect 18092 23428 18156 23432
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 17908 23156 17972 23220
rect 12204 23020 12268 23084
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 20668 22808 20732 22812
rect 20668 22752 20718 22808
rect 20718 22752 20732 22808
rect 20668 22748 20732 22752
rect 25084 22748 25148 22812
rect 25636 22748 25700 22812
rect 12020 22612 12084 22676
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 26004 22204 26068 22268
rect 22324 22068 22388 22132
rect 22876 22068 22940 22132
rect 24348 22068 24412 22132
rect 28028 22068 28092 22132
rect 23612 21932 23676 21996
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 17172 21660 17236 21724
rect 20300 21524 20364 21588
rect 23060 21660 23124 21724
rect 25820 21388 25884 21452
rect 23980 21252 24044 21316
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 20116 20572 20180 20636
rect 24900 20300 24964 20364
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 26003 31924 26069 31925
rect 26003 31860 26004 31924
rect 26068 31860 26069 31924
rect 26003 31859 26069 31860
rect 23243 31788 23309 31789
rect 23243 31724 23244 31788
rect 23308 31724 23309 31788
rect 23243 31723 23309 31724
rect 4417 31040 4737 31600
rect 4417 30976 4425 31040
rect 4489 30976 4505 31040
rect 4569 30976 4585 31040
rect 4649 30976 4665 31040
rect 4729 30976 4737 31040
rect 4417 29952 4737 30976
rect 4417 29888 4425 29952
rect 4489 29888 4505 29952
rect 4569 29888 4585 29952
rect 4649 29888 4665 29952
rect 4729 29888 4737 29952
rect 4417 28864 4737 29888
rect 4417 28800 4425 28864
rect 4489 28800 4505 28864
rect 4569 28800 4585 28864
rect 4649 28800 4665 28864
rect 4729 28800 4737 28864
rect 4417 27776 4737 28800
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 31584 8210 31600
rect 7890 31520 7898 31584
rect 7962 31520 7978 31584
rect 8042 31520 8058 31584
rect 8122 31520 8138 31584
rect 8202 31520 8210 31584
rect 7890 30496 8210 31520
rect 7890 30432 7898 30496
rect 7962 30432 7978 30496
rect 8042 30432 8058 30496
rect 8122 30432 8138 30496
rect 8202 30432 8210 30496
rect 7890 29408 8210 30432
rect 11363 31040 11683 31600
rect 11363 30976 11371 31040
rect 11435 30976 11451 31040
rect 11515 30976 11531 31040
rect 11595 30976 11611 31040
rect 11675 30976 11683 31040
rect 9995 30156 10061 30157
rect 9995 30092 9996 30156
rect 10060 30092 10061 30156
rect 9995 30091 10061 30092
rect 7890 29344 7898 29408
rect 7962 29344 7978 29408
rect 8042 29344 8058 29408
rect 8122 29344 8138 29408
rect 8202 29344 8210 29408
rect 7890 28320 8210 29344
rect 9998 29069 10058 30091
rect 11363 29952 11683 30976
rect 14836 31584 15156 31600
rect 14836 31520 14844 31584
rect 14908 31520 14924 31584
rect 14988 31520 15004 31584
rect 15068 31520 15084 31584
rect 15148 31520 15156 31584
rect 14836 30496 15156 31520
rect 18309 31040 18629 31600
rect 21782 31584 22102 31600
rect 21782 31520 21790 31584
rect 21854 31520 21870 31584
rect 21934 31520 21950 31584
rect 22014 31520 22030 31584
rect 22094 31520 22102 31584
rect 21219 31516 21285 31517
rect 21219 31452 21220 31516
rect 21284 31452 21285 31516
rect 21219 31451 21285 31452
rect 18827 31108 18893 31109
rect 18827 31044 18828 31108
rect 18892 31044 18893 31108
rect 18827 31043 18893 31044
rect 18309 30976 18317 31040
rect 18381 30976 18397 31040
rect 18461 30976 18477 31040
rect 18541 30976 18557 31040
rect 18621 30976 18629 31040
rect 17355 30700 17421 30701
rect 17355 30636 17356 30700
rect 17420 30636 17421 30700
rect 17355 30635 17421 30636
rect 17907 30700 17973 30701
rect 17907 30636 17908 30700
rect 17972 30636 17973 30700
rect 17907 30635 17973 30636
rect 14836 30432 14844 30496
rect 14908 30432 14924 30496
rect 14988 30432 15004 30496
rect 15068 30432 15084 30496
rect 15148 30432 15156 30496
rect 12019 30428 12085 30429
rect 12019 30364 12020 30428
rect 12084 30364 12085 30428
rect 12019 30363 12085 30364
rect 11363 29888 11371 29952
rect 11435 29888 11451 29952
rect 11515 29888 11531 29952
rect 11595 29888 11611 29952
rect 11675 29888 11683 29952
rect 9995 29068 10061 29069
rect 9995 29004 9996 29068
rect 10060 29004 10061 29068
rect 9995 29003 10061 29004
rect 10915 29068 10981 29069
rect 10915 29004 10916 29068
rect 10980 29004 10981 29068
rect 10915 29003 10981 29004
rect 7890 28256 7898 28320
rect 7962 28256 7978 28320
rect 8042 28256 8058 28320
rect 8122 28256 8138 28320
rect 8202 28256 8210 28320
rect 7890 27232 8210 28256
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 10918 25805 10978 29003
rect 11363 28864 11683 29888
rect 11363 28800 11371 28864
rect 11435 28800 11451 28864
rect 11515 28800 11531 28864
rect 11595 28800 11611 28864
rect 11675 28800 11683 28864
rect 11363 27776 11683 28800
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 10915 25804 10981 25805
rect 10915 25740 10916 25804
rect 10980 25740 10981 25804
rect 10915 25739 10981 25740
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 12022 22677 12082 30363
rect 14836 29408 15156 30432
rect 15331 30292 15397 30293
rect 15331 30228 15332 30292
rect 15396 30228 15397 30292
rect 15331 30227 15397 30228
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 12203 29068 12269 29069
rect 12203 29004 12204 29068
rect 12268 29004 12269 29068
rect 12203 29003 12269 29004
rect 14595 29068 14661 29069
rect 14595 29004 14596 29068
rect 14660 29004 14661 29068
rect 14595 29003 14661 29004
rect 12206 23085 12266 29003
rect 14411 28932 14477 28933
rect 14411 28868 14412 28932
rect 14476 28868 14477 28932
rect 14411 28867 14477 28868
rect 14414 27301 14474 28867
rect 13491 27300 13557 27301
rect 13491 27236 13492 27300
rect 13556 27236 13557 27300
rect 13491 27235 13557 27236
rect 14411 27300 14477 27301
rect 14411 27236 14412 27300
rect 14476 27236 14477 27300
rect 14411 27235 14477 27236
rect 13494 23765 13554 27235
rect 14598 25397 14658 29003
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 15334 27709 15394 30227
rect 16803 30020 16869 30021
rect 16803 29956 16804 30020
rect 16868 29956 16869 30020
rect 16803 29955 16869 29956
rect 15883 29476 15949 29477
rect 15883 29412 15884 29476
rect 15948 29412 15949 29476
rect 15883 29411 15949 29412
rect 15515 28252 15581 28253
rect 15515 28188 15516 28252
rect 15580 28188 15581 28252
rect 15515 28187 15581 28188
rect 15331 27708 15397 27709
rect 15331 27644 15332 27708
rect 15396 27644 15397 27708
rect 15331 27643 15397 27644
rect 15518 27301 15578 28187
rect 15515 27300 15581 27301
rect 15515 27236 15516 27300
rect 15580 27236 15581 27300
rect 15515 27235 15581 27236
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 15886 27165 15946 29411
rect 16619 29340 16685 29341
rect 16619 29276 16620 29340
rect 16684 29338 16685 29340
rect 16806 29338 16866 29955
rect 16684 29278 16866 29338
rect 16684 29276 16685 29278
rect 16619 29275 16685 29276
rect 17358 29069 17418 30635
rect 17910 30290 17970 30635
rect 17910 30230 18154 30290
rect 18094 29885 18154 30230
rect 18309 29952 18629 30976
rect 18309 29888 18317 29952
rect 18381 29888 18397 29952
rect 18461 29888 18477 29952
rect 18541 29888 18557 29952
rect 18621 29888 18629 29952
rect 18091 29884 18157 29885
rect 18091 29820 18092 29884
rect 18156 29820 18157 29884
rect 18091 29819 18157 29820
rect 18091 29476 18157 29477
rect 18091 29412 18092 29476
rect 18156 29412 18157 29476
rect 18091 29411 18157 29412
rect 17723 29340 17789 29341
rect 17723 29276 17724 29340
rect 17788 29276 17789 29340
rect 17723 29275 17789 29276
rect 17171 29068 17237 29069
rect 17171 29004 17172 29068
rect 17236 29004 17237 29068
rect 17171 29003 17237 29004
rect 17355 29068 17421 29069
rect 17355 29004 17356 29068
rect 17420 29004 17421 29068
rect 17355 29003 17421 29004
rect 16067 27300 16133 27301
rect 16067 27236 16068 27300
rect 16132 27236 16133 27300
rect 16067 27235 16133 27236
rect 16619 27300 16685 27301
rect 16619 27236 16620 27300
rect 16684 27236 16685 27300
rect 16619 27235 16685 27236
rect 15883 27164 15949 27165
rect 15883 27100 15884 27164
rect 15948 27100 15949 27164
rect 15883 27099 15949 27100
rect 16070 26213 16130 27235
rect 16622 26349 16682 27235
rect 16619 26348 16685 26349
rect 16619 26284 16620 26348
rect 16684 26284 16685 26348
rect 16619 26283 16685 26284
rect 16067 26212 16133 26213
rect 16067 26148 16068 26212
rect 16132 26148 16133 26212
rect 16067 26147 16133 26148
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14595 25396 14661 25397
rect 14595 25332 14596 25396
rect 14660 25332 14661 25396
rect 14595 25331 14661 25332
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 16622 24989 16682 26283
rect 16619 24988 16685 24989
rect 16619 24924 16620 24988
rect 16684 24924 16685 24988
rect 16619 24923 16685 24924
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 13491 23764 13557 23765
rect 13491 23700 13492 23764
rect 13556 23700 13557 23764
rect 13491 23699 13557 23700
rect 12203 23084 12269 23085
rect 12203 23020 12204 23084
rect 12268 23020 12269 23084
rect 12203 23019 12269 23020
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 12019 22676 12085 22677
rect 12019 22612 12020 22676
rect 12084 22612 12085 22676
rect 12019 22611 12085 22612
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 17174 21725 17234 29003
rect 17539 27844 17605 27845
rect 17539 27780 17540 27844
rect 17604 27780 17605 27844
rect 17539 27779 17605 27780
rect 17542 26077 17602 27779
rect 17539 26076 17605 26077
rect 17539 26012 17540 26076
rect 17604 26012 17605 26076
rect 17539 26011 17605 26012
rect 17726 24717 17786 29275
rect 17907 27708 17973 27709
rect 17907 27644 17908 27708
rect 17972 27644 17973 27708
rect 17907 27643 17973 27644
rect 17723 24716 17789 24717
rect 17723 24652 17724 24716
rect 17788 24652 17789 24716
rect 17723 24651 17789 24652
rect 17910 23221 17970 27643
rect 18094 23493 18154 29411
rect 18309 28864 18629 29888
rect 18830 29341 18890 31043
rect 19931 30564 19997 30565
rect 19931 30500 19932 30564
rect 19996 30500 19997 30564
rect 19931 30499 19997 30500
rect 19195 30156 19261 30157
rect 19195 30092 19196 30156
rect 19260 30092 19261 30156
rect 19195 30091 19261 30092
rect 18827 29340 18893 29341
rect 18827 29276 18828 29340
rect 18892 29276 18893 29340
rect 18827 29275 18893 29276
rect 18309 28800 18317 28864
rect 18381 28800 18397 28864
rect 18461 28800 18477 28864
rect 18541 28800 18557 28864
rect 18621 28800 18629 28864
rect 18309 27776 18629 28800
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18830 24853 18890 29275
rect 19198 26757 19258 30091
rect 19379 29612 19445 29613
rect 19379 29548 19380 29612
rect 19444 29548 19445 29612
rect 19379 29547 19445 29548
rect 19195 26756 19261 26757
rect 19195 26692 19196 26756
rect 19260 26692 19261 26756
rect 19195 26691 19261 26692
rect 19382 26077 19442 29547
rect 19379 26076 19445 26077
rect 19379 26012 19380 26076
rect 19444 26012 19445 26076
rect 19379 26011 19445 26012
rect 19747 26076 19813 26077
rect 19747 26012 19748 26076
rect 19812 26012 19813 26076
rect 19747 26011 19813 26012
rect 18827 24852 18893 24853
rect 18827 24788 18828 24852
rect 18892 24788 18893 24852
rect 18827 24787 18893 24788
rect 19750 24581 19810 26011
rect 19934 25941 19994 30499
rect 20483 30428 20549 30429
rect 20483 30364 20484 30428
rect 20548 30364 20549 30428
rect 20483 30363 20549 30364
rect 20299 27708 20365 27709
rect 20299 27644 20300 27708
rect 20364 27644 20365 27708
rect 20299 27643 20365 27644
rect 19931 25940 19997 25941
rect 19931 25876 19932 25940
rect 19996 25876 19997 25940
rect 19931 25875 19997 25876
rect 19931 25124 19997 25125
rect 19931 25060 19932 25124
rect 19996 25060 19997 25124
rect 19931 25059 19997 25060
rect 19747 24580 19813 24581
rect 19747 24516 19748 24580
rect 19812 24516 19813 24580
rect 19747 24515 19813 24516
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18091 23492 18157 23493
rect 18091 23428 18092 23492
rect 18156 23428 18157 23492
rect 18091 23427 18157 23428
rect 18309 23424 18629 24448
rect 19934 23629 19994 25059
rect 20115 23900 20181 23901
rect 20115 23836 20116 23900
rect 20180 23836 20181 23900
rect 20115 23835 20181 23836
rect 19931 23628 19997 23629
rect 19931 23564 19932 23628
rect 19996 23564 19997 23628
rect 19931 23563 19997 23564
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 17907 23220 17973 23221
rect 17907 23156 17908 23220
rect 17972 23156 17973 23220
rect 17907 23155 17973 23156
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 17171 21724 17237 21725
rect 17171 21660 17172 21724
rect 17236 21660 17237 21724
rect 17171 21659 17237 21660
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 20118 20637 20178 23835
rect 20302 21589 20362 27643
rect 20486 25941 20546 30363
rect 20667 30020 20733 30021
rect 20667 29956 20668 30020
rect 20732 29956 20733 30020
rect 20667 29955 20733 29956
rect 20670 27573 20730 29955
rect 20851 29748 20917 29749
rect 20851 29684 20852 29748
rect 20916 29684 20917 29748
rect 20851 29683 20917 29684
rect 20667 27572 20733 27573
rect 20667 27508 20668 27572
rect 20732 27508 20733 27572
rect 20667 27507 20733 27508
rect 20667 26756 20733 26757
rect 20667 26692 20668 26756
rect 20732 26692 20733 26756
rect 20667 26691 20733 26692
rect 20483 25940 20549 25941
rect 20483 25876 20484 25940
rect 20548 25876 20549 25940
rect 20483 25875 20549 25876
rect 20670 22813 20730 26691
rect 20854 26485 20914 29683
rect 20851 26484 20917 26485
rect 20851 26420 20852 26484
rect 20916 26420 20917 26484
rect 20851 26419 20917 26420
rect 21222 23765 21282 31451
rect 21782 30496 22102 31520
rect 23059 30700 23125 30701
rect 23059 30636 23060 30700
rect 23124 30636 23125 30700
rect 23059 30635 23125 30636
rect 21782 30432 21790 30496
rect 21854 30432 21870 30496
rect 21934 30432 21950 30496
rect 22014 30432 22030 30496
rect 22094 30432 22102 30496
rect 21782 29408 22102 30432
rect 21782 29344 21790 29408
rect 21854 29344 21870 29408
rect 21934 29344 21950 29408
rect 22014 29344 22030 29408
rect 22094 29344 22102 29408
rect 21782 28320 22102 29344
rect 22875 28932 22941 28933
rect 22875 28868 22876 28932
rect 22940 28868 22941 28932
rect 22875 28867 22941 28868
rect 21782 28256 21790 28320
rect 21854 28256 21870 28320
rect 21934 28256 21950 28320
rect 22014 28256 22030 28320
rect 22094 28256 22102 28320
rect 21782 27232 22102 28256
rect 22691 27300 22757 27301
rect 22691 27236 22692 27300
rect 22756 27236 22757 27300
rect 22691 27235 22757 27236
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 22323 27164 22389 27165
rect 22323 27100 22324 27164
rect 22388 27100 22389 27164
rect 22323 27099 22389 27100
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21219 23764 21285 23765
rect 21219 23700 21220 23764
rect 21284 23700 21285 23764
rect 21219 23699 21285 23700
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 20667 22812 20733 22813
rect 20667 22748 20668 22812
rect 20732 22748 20733 22812
rect 20667 22747 20733 22748
rect 21782 21792 22102 22816
rect 22326 22133 22386 27099
rect 22694 24037 22754 27235
rect 22691 24036 22757 24037
rect 22691 23972 22692 24036
rect 22756 23972 22757 24036
rect 22691 23971 22757 23972
rect 22878 22133 22938 28867
rect 23062 26077 23122 30635
rect 23059 26076 23125 26077
rect 23059 26012 23060 26076
rect 23124 26012 23125 26076
rect 23059 26011 23125 26012
rect 22323 22132 22389 22133
rect 22323 22068 22324 22132
rect 22388 22068 22389 22132
rect 22323 22067 22389 22068
rect 22875 22132 22941 22133
rect 22875 22068 22876 22132
rect 22940 22068 22941 22132
rect 22875 22067 22941 22068
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 20299 21588 20365 21589
rect 20299 21524 20300 21588
rect 20364 21524 20365 21588
rect 20299 21523 20365 21524
rect 21782 20704 22102 21728
rect 23062 21725 23122 26011
rect 23246 24989 23306 31723
rect 25255 31040 25575 31600
rect 25255 30976 25263 31040
rect 25327 30976 25343 31040
rect 25407 30976 25423 31040
rect 25487 30976 25503 31040
rect 25567 30976 25575 31040
rect 23427 30972 23493 30973
rect 23427 30908 23428 30972
rect 23492 30908 23493 30972
rect 23427 30907 23493 30908
rect 23430 27573 23490 30907
rect 25083 30020 25149 30021
rect 25083 29956 25084 30020
rect 25148 29956 25149 30020
rect 25083 29955 25149 29956
rect 23795 28660 23861 28661
rect 23795 28596 23796 28660
rect 23860 28596 23861 28660
rect 23795 28595 23861 28596
rect 23611 27708 23677 27709
rect 23611 27644 23612 27708
rect 23676 27644 23677 27708
rect 23611 27643 23677 27644
rect 23427 27572 23493 27573
rect 23427 27508 23428 27572
rect 23492 27508 23493 27572
rect 23427 27507 23493 27508
rect 23243 24988 23309 24989
rect 23243 24924 23244 24988
rect 23308 24924 23309 24988
rect 23243 24923 23309 24924
rect 23614 21997 23674 27643
rect 23798 26213 23858 28595
rect 24715 28524 24781 28525
rect 24715 28460 24716 28524
rect 24780 28460 24781 28524
rect 24715 28459 24781 28460
rect 24531 28252 24597 28253
rect 24531 28188 24532 28252
rect 24596 28188 24597 28252
rect 24531 28187 24597 28188
rect 24347 26484 24413 26485
rect 24347 26420 24348 26484
rect 24412 26420 24413 26484
rect 24347 26419 24413 26420
rect 23795 26212 23861 26213
rect 23795 26148 23796 26212
rect 23860 26148 23861 26212
rect 23795 26147 23861 26148
rect 23979 26212 24045 26213
rect 23979 26148 23980 26212
rect 24044 26148 24045 26212
rect 23979 26147 24045 26148
rect 23611 21996 23677 21997
rect 23611 21932 23612 21996
rect 23676 21932 23677 21996
rect 23611 21931 23677 21932
rect 23059 21724 23125 21725
rect 23059 21660 23060 21724
rect 23124 21660 23125 21724
rect 23059 21659 23125 21660
rect 23982 21317 24042 26147
rect 24350 22133 24410 26419
rect 24534 24853 24594 28187
rect 24718 27029 24778 28459
rect 24899 27164 24965 27165
rect 24899 27100 24900 27164
rect 24964 27100 24965 27164
rect 24899 27099 24965 27100
rect 24715 27028 24781 27029
rect 24715 26964 24716 27028
rect 24780 26964 24781 27028
rect 24715 26963 24781 26964
rect 24531 24852 24597 24853
rect 24531 24788 24532 24852
rect 24596 24788 24597 24852
rect 24531 24787 24597 24788
rect 24347 22132 24413 22133
rect 24347 22068 24348 22132
rect 24412 22068 24413 22132
rect 24347 22067 24413 22068
rect 23979 21316 24045 21317
rect 23979 21252 23980 21316
rect 24044 21252 24045 21316
rect 23979 21251 24045 21252
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 20115 20636 20181 20637
rect 20115 20572 20116 20636
rect 20180 20572 20181 20636
rect 20115 20571 20181 20572
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 19616 22102 20640
rect 24902 20365 24962 27099
rect 25086 26893 25146 29955
rect 25255 29952 25575 30976
rect 25255 29888 25263 29952
rect 25327 29888 25343 29952
rect 25407 29888 25423 29952
rect 25487 29888 25503 29952
rect 25567 29888 25575 29952
rect 25255 28864 25575 29888
rect 25255 28800 25263 28864
rect 25327 28800 25343 28864
rect 25407 28800 25423 28864
rect 25487 28800 25503 28864
rect 25567 28800 25575 28864
rect 25255 27776 25575 28800
rect 25819 28524 25885 28525
rect 25819 28460 25820 28524
rect 25884 28460 25885 28524
rect 25819 28459 25885 28460
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25083 26892 25149 26893
rect 25083 26828 25084 26892
rect 25148 26828 25149 26892
rect 25083 26827 25149 26828
rect 25086 26077 25146 26827
rect 25255 26688 25575 27712
rect 25635 26892 25701 26893
rect 25635 26828 25636 26892
rect 25700 26828 25701 26892
rect 25635 26827 25701 26828
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25083 26076 25149 26077
rect 25083 26012 25084 26076
rect 25148 26012 25149 26076
rect 25083 26011 25149 26012
rect 25083 25668 25149 25669
rect 25083 25604 25084 25668
rect 25148 25604 25149 25668
rect 25083 25603 25149 25604
rect 25086 24717 25146 25603
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25083 24716 25149 24717
rect 25083 24652 25084 24716
rect 25148 24652 25149 24716
rect 25083 24651 25149 24652
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25083 24036 25149 24037
rect 25083 23972 25084 24036
rect 25148 23972 25149 24036
rect 25083 23971 25149 23972
rect 25086 22813 25146 23971
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25083 22812 25149 22813
rect 25083 22748 25084 22812
rect 25148 22748 25149 22812
rect 25083 22747 25149 22748
rect 25255 22336 25575 23360
rect 25638 22813 25698 26827
rect 25822 25397 25882 28459
rect 26006 25533 26066 31859
rect 28728 31584 29048 31600
rect 28728 31520 28736 31584
rect 28800 31520 28816 31584
rect 28880 31520 28896 31584
rect 28960 31520 28976 31584
rect 29040 31520 29048 31584
rect 28728 30496 29048 31520
rect 28728 30432 28736 30496
rect 28800 30432 28816 30496
rect 28880 30432 28896 30496
rect 28960 30432 28976 30496
rect 29040 30432 29048 30496
rect 28728 29408 29048 30432
rect 28728 29344 28736 29408
rect 28800 29344 28816 29408
rect 28880 29344 28896 29408
rect 28960 29344 28976 29408
rect 29040 29344 29048 29408
rect 27475 28388 27541 28389
rect 27475 28324 27476 28388
rect 27540 28324 27541 28388
rect 27475 28323 27541 28324
rect 27478 27981 27538 28323
rect 28728 28320 29048 29344
rect 28728 28256 28736 28320
rect 28800 28256 28816 28320
rect 28880 28256 28896 28320
rect 28960 28256 28976 28320
rect 29040 28256 29048 28320
rect 26187 27980 26253 27981
rect 26187 27916 26188 27980
rect 26252 27916 26253 27980
rect 26187 27915 26253 27916
rect 27475 27980 27541 27981
rect 27475 27916 27476 27980
rect 27540 27916 27541 27980
rect 27475 27915 27541 27916
rect 26003 25532 26069 25533
rect 26003 25468 26004 25532
rect 26068 25468 26069 25532
rect 26003 25467 26069 25468
rect 26190 25397 26250 27915
rect 26371 26076 26437 26077
rect 26371 26012 26372 26076
rect 26436 26012 26437 26076
rect 26371 26011 26437 26012
rect 25819 25396 25885 25397
rect 25819 25332 25820 25396
rect 25884 25332 25885 25396
rect 25819 25331 25885 25332
rect 26187 25396 26253 25397
rect 26187 25332 26188 25396
rect 26252 25332 26253 25396
rect 26187 25331 26253 25332
rect 26003 24852 26069 24853
rect 26003 24788 26004 24852
rect 26068 24788 26069 24852
rect 26003 24787 26069 24788
rect 25819 23900 25885 23901
rect 25819 23836 25820 23900
rect 25884 23836 25885 23900
rect 25819 23835 25885 23836
rect 25635 22812 25701 22813
rect 25635 22748 25636 22812
rect 25700 22748 25701 22812
rect 25635 22747 25701 22748
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25822 21453 25882 23835
rect 26006 22269 26066 24787
rect 26190 23901 26250 25331
rect 26374 24037 26434 26011
rect 27478 24309 27538 27915
rect 28728 27232 29048 28256
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28027 26484 28093 26485
rect 28027 26420 28028 26484
rect 28092 26420 28093 26484
rect 28027 26419 28093 26420
rect 27475 24308 27541 24309
rect 27475 24244 27476 24308
rect 27540 24244 27541 24308
rect 27475 24243 27541 24244
rect 26371 24036 26437 24037
rect 26371 23972 26372 24036
rect 26436 23972 26437 24036
rect 26371 23971 26437 23972
rect 26187 23900 26253 23901
rect 26187 23836 26188 23900
rect 26252 23836 26253 23900
rect 26187 23835 26253 23836
rect 26003 22268 26069 22269
rect 26003 22204 26004 22268
rect 26068 22204 26069 22268
rect 26003 22203 26069 22204
rect 28030 22133 28090 26419
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28027 22132 28093 22133
rect 28027 22068 28028 22132
rect 28092 22068 28093 22132
rect 28027 22067 28093 22068
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 25819 21452 25885 21453
rect 25819 21388 25820 21452
rect 25884 21388 25885 21452
rect 25819 21387 25885 21388
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 24899 20364 24965 20365
rect 24899 20300 24900 20364
rect 24964 20300 24965 20364
rect 24899 20299 24965 20300
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1666464484
transform 1 0 22632 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__B
timestamp 1666464484
transform -1 0 27140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__C
timestamp 1666464484
transform -1 0 27324 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A2
timestamp 1666464484
transform 1 0 15272 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__B1
timestamp 1666464484
transform 1 0 15088 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1666464484
transform -1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1666464484
transform -1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1666464484
transform -1 0 10580 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__B
timestamp 1666464484
transform 1 0 4600 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__C
timestamp 1666464484
transform 1 0 9752 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A2
timestamp 1666464484
transform 1 0 25852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__B1
timestamp 1666464484
transform -1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__C1
timestamp 1666464484
transform -1 0 26588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A1
timestamp 1666464484
transform -1 0 5244 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A2
timestamp 1666464484
transform 1 0 6164 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__B
timestamp 1666464484
transform 1 0 19596 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__C
timestamp 1666464484
transform 1 0 19780 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A2
timestamp 1666464484
transform 1 0 13616 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__B
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__C
timestamp 1666464484
transform 1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A2
timestamp 1666464484
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__B1
timestamp 1666464484
transform 1 0 15640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__B
timestamp 1666464484
transform 1 0 11040 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__C
timestamp 1666464484
transform 1 0 12052 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A2
timestamp 1666464484
transform -1 0 5796 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__B1
timestamp 1666464484
transform -1 0 6900 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__B
timestamp 1666464484
transform 1 0 20700 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__C
timestamp 1666464484
transform 1 0 20884 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A2
timestamp 1666464484
transform 1 0 13524 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__B1
timestamp 1666464484
transform 1 0 14076 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__B
timestamp 1666464484
transform 1 0 19688 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__C
timestamp 1666464484
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A2
timestamp 1666464484
transform 1 0 7728 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__B1
timestamp 1666464484
transform 1 0 9384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A1
timestamp 1666464484
transform 1 0 6808 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A2
timestamp 1666464484
transform 1 0 8464 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__B
timestamp 1666464484
transform -1 0 22172 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__C
timestamp 1666464484
transform -1 0 21620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A1
timestamp 1666464484
transform 1 0 25300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A2
timestamp 1666464484
transform -1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__B
timestamp 1666464484
transform 1 0 11040 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__C
timestamp 1666464484
transform 1 0 11960 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A2
timestamp 1666464484
transform 1 0 7360 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__B1
timestamp 1666464484
transform -1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__B
timestamp 1666464484
transform 1 0 23644 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__C
timestamp 1666464484
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A1
timestamp 1666464484
transform 1 0 19412 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A2
timestamp 1666464484
transform 1 0 17112 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__B1
timestamp 1666464484
transform 1 0 17204 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__B
timestamp 1666464484
transform -1 0 25300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__C
timestamp 1666464484
transform -1 0 26128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A2
timestamp 1666464484
transform -1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__B1
timestamp 1666464484
transform 1 0 20516 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A1
timestamp 1666464484
transform 1 0 18216 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A2
timestamp 1666464484
transform 1 0 16100 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__B
timestamp 1666464484
transform 1 0 10304 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__C
timestamp 1666464484
transform 1 0 6716 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A1
timestamp 1666464484
transform 1 0 8464 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__B
timestamp 1666464484
transform 1 0 26220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__C
timestamp 1666464484
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A2
timestamp 1666464484
transform 1 0 14628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__B1
timestamp 1666464484
transform 1 0 12420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__B
timestamp 1666464484
transform -1 0 26404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__C
timestamp 1666464484
transform -1 0 26220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A2
timestamp 1666464484
transform -1 0 27324 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__B1
timestamp 1666464484
transform -1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__B
timestamp 1666464484
transform 1 0 14628 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__C
timestamp 1666464484
transform 1 0 16192 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A2
timestamp 1666464484
transform -1 0 7452 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__B1
timestamp 1666464484
transform -1 0 8004 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A1
timestamp 1666464484
transform 1 0 9844 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A2
timestamp 1666464484
transform 1 0 9384 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__B
timestamp 1666464484
transform -1 0 4416 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__C
timestamp 1666464484
transform -1 0 5336 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A1
timestamp 1666464484
transform 1 0 25300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A3
timestamp 1666464484
transform -1 0 25668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__B
timestamp 1666464484
transform 1 0 23736 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__C
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A2
timestamp 1666464484
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__B1
timestamp 1666464484
transform 1 0 14720 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__B
timestamp 1666464484
transform -1 0 4692 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__C
timestamp 1666464484
transform -1 0 6440 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A2
timestamp 1666464484
transform 1 0 11868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__B1
timestamp 1666464484
transform 1 0 9936 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__B
timestamp 1666464484
transform 1 0 17756 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__C
timestamp 1666464484
transform 1 0 17940 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A2
timestamp 1666464484
transform 1 0 9476 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__B1
timestamp 1666464484
transform 1 0 9568 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A1
timestamp 1666464484
transform 1 0 14996 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A2
timestamp 1666464484
transform 1 0 14444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__B
timestamp 1666464484
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__C
timestamp 1666464484
transform 1 0 25116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A1
timestamp 1666464484
transform 1 0 16836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__B
timestamp 1666464484
transform 1 0 12512 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__C
timestamp 1666464484
transform 1 0 13064 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A2
timestamp 1666464484
transform 1 0 16192 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__B1
timestamp 1666464484
transform 1 0 13616 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__B
timestamp 1666464484
transform 1 0 17848 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__C
timestamp 1666464484
transform 1 0 18308 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A2
timestamp 1666464484
transform -1 0 5520 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B1
timestamp 1666464484
transform 1 0 6532 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__B
timestamp 1666464484
transform 1 0 18952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__C
timestamp 1666464484
transform 1 0 15824 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A2
timestamp 1666464484
transform 1 0 23368 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__B1
timestamp 1666464484
transform 1 0 24564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A1
timestamp 1666464484
transform 1 0 7084 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A2
timestamp 1666464484
transform -1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__B
timestamp 1666464484
transform 1 0 18768 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__C
timestamp 1666464484
transform 1 0 16652 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A1
timestamp 1666464484
transform 1 0 22908 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__B
timestamp 1666464484
transform -1 0 4140 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__C
timestamp 1666464484
transform -1 0 4968 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A2
timestamp 1666464484
transform -1 0 24472 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__B1
timestamp 1666464484
transform -1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__C1
timestamp 1666464484
transform -1 0 23368 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__B
timestamp 1666464484
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__C
timestamp 1666464484
transform 1 0 25668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A2
timestamp 1666464484
transform 1 0 26220 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__B1
timestamp 1666464484
transform 1 0 26772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__B
timestamp 1666464484
transform 1 0 16928 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__C
timestamp 1666464484
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A2
timestamp 1666464484
transform 1 0 8280 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__B1
timestamp 1666464484
transform 1 0 8464 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A1
timestamp 1666464484
transform 1 0 12144 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A2
timestamp 1666464484
transform 1 0 12696 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__B
timestamp 1666464484
transform 1 0 22264 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__C
timestamp 1666464484
transform 1 0 25024 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A1
timestamp 1666464484
transform -1 0 19596 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__B
timestamp 1666464484
transform 1 0 10856 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__C
timestamp 1666464484
transform 1 0 8832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A2
timestamp 1666464484
transform -1 0 20608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__B1
timestamp 1666464484
transform 1 0 21068 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__B
timestamp 1666464484
transform 1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__C
timestamp 1666464484
transform 1 0 24840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A2
timestamp 1666464484
transform 1 0 20976 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__B1
timestamp 1666464484
transform 1 0 26496 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1666464484
transform -1 0 10580 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1666464484
transform 1 0 10488 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__C
timestamp 1666464484
transform 1 0 11408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A2
timestamp 1666464484
transform 1 0 10948 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__B1
timestamp 1666464484
transform 1 0 11500 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A1
timestamp 1666464484
transform 1 0 7360 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A2
timestamp 1666464484
transform 1 0 7912 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__B
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__C
timestamp 1666464484
transform 1 0 19228 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A1
timestamp 1666464484
transform -1 0 27140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__CLK
timestamp 1666464484
transform 1 0 24748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__CLK
timestamp 1666464484
transform 1 0 13064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__CLK
timestamp 1666464484
transform 1 0 13892 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__CLK
timestamp 1666464484
transform 1 0 8924 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__CLK
timestamp 1666464484
transform -1 0 6716 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__CLK
timestamp 1666464484
transform 1 0 12972 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__CLK
timestamp 1666464484
transform 1 0 24472 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__CLK
timestamp 1666464484
transform 1 0 12052 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__CLK
timestamp 1666464484
transform 1 0 21988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__CLK
timestamp 1666464484
transform 1 0 23460 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__CLK
timestamp 1666464484
transform -1 0 26220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__CLK
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__CLK
timestamp 1666464484
transform 1 0 10488 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__CLK
timestamp 1666464484
transform -1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__CLK
timestamp 1666464484
transform -1 0 25208 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__CLK
timestamp 1666464484
transform -1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__CLK
timestamp 1666464484
transform 1 0 5888 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__CLK
timestamp 1666464484
transform 1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__CLK
timestamp 1666464484
transform -1 0 28428 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__CLK
timestamp 1666464484
transform 1 0 10120 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__CLK
timestamp 1666464484
transform -1 0 5888 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__CLK
timestamp 1666464484
transform -1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__CLK
timestamp 1666464484
transform -1 0 25668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__CLK
timestamp 1666464484
transform -1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__CLK
timestamp 1666464484
transform -1 0 24104 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__CLK
timestamp 1666464484
transform -1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__CLK
timestamp 1666464484
transform 1 0 17664 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__CLK
timestamp 1666464484
transform 1 0 8188 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__CLK
timestamp 1666464484
transform 1 0 22356 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__D
timestamp 1666464484
transform -1 0 20056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__D
timestamp 1666464484
transform -1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__CLK
timestamp 1666464484
transform 1 0 7912 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__CLK
timestamp 1666464484
transform -1 0 3496 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__CLK
timestamp 1666464484
transform 1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__CLK
timestamp 1666464484
transform -1 0 26404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__CLK
timestamp 1666464484
transform 1 0 7820 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__CLK
timestamp 1666464484
transform 1 0 18676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__CLK
timestamp 1666464484
transform 1 0 11040 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__CLK
timestamp 1666464484
transform -1 0 7820 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__D
timestamp 1666464484
transform -1 0 8556 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__CLK
timestamp 1666464484
transform -1 0 6992 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1666464484
transform -1 0 6440 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1666464484
transform -1 0 7360 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout17_A
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout18_A
timestamp 1666464484
transform 1 0 15548 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout19_A
timestamp 1666464484
transform -1 0 23920 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout20_A
timestamp 1666464484
transform 1 0 9292 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout21_A
timestamp 1666464484
transform 1 0 9936 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout22_A
timestamp 1666464484
transform -1 0 27784 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout23_A
timestamp 1666464484
transform -1 0 8096 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 27784 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 27876 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 27232 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 27784 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 27324 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 28428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 27784 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1666464484
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_293
timestamp 1666464484
transform 1 0 28060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1666464484
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1666464484
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1666464484
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1666464484
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1666464484
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1666464484
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1666464484
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1666464484
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1666464484
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1666464484
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_293
timestamp 1666464484
transform 1 0 28060 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1666464484
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_8
timestamp 1666464484
transform 1 0 1840 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_20
timestamp 1666464484
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1666464484
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1666464484
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_293
timestamp 1666464484
transform 1 0 28060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp 1666464484
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1666464484
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1666464484
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1666464484
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1666464484
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666464484
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1666464484
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1666464484
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666464484
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1666464484
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666464484
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1666464484
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_293
timestamp 1666464484
transform 1 0 28060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp 1666464484
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1666464484
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1666464484
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1666464484
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_293
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1666464484
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1666464484
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1666464484
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1666464484
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1666464484
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp 1666464484
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1666464484
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1666464484
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1666464484
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1666464484
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1666464484
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_293
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1666464484
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_8
timestamp 1666464484
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1666464484
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1666464484
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1666464484
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666464484
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1666464484
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1666464484
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_293
timestamp 1666464484
transform 1 0 28060 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1666464484
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1666464484
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1666464484
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1666464484
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666464484
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666464484
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1666464484
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1666464484
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666464484
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666464484
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666464484
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1666464484
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_8
timestamp 1666464484
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1666464484
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666464484
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666464484
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666464484
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666464484
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1666464484
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1666464484
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1666464484
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1666464484
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1666464484
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666464484
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666464484
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1666464484
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_290
timestamp 1666464484
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1666464484
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666464484
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_265
timestamp 1666464484
transform 1 0 25484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_275
timestamp 1666464484
transform 1 0 26404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_283
timestamp 1666464484
transform 1 0 27140 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_289
timestamp 1666464484
transform 1 0 27692 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_292
timestamp 1666464484
transform 1 0 27968 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1666464484
transform 1 0 28520 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_249
timestamp 1666464484
transform 1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_257
timestamp 1666464484
transform 1 0 24748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1666464484
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_267
timestamp 1666464484
transform 1 0 25668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666464484
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_285
timestamp 1666464484
transform 1 0 27324 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1666464484
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_8
timestamp 1666464484
transform 1 0 1840 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1666464484
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_257
timestamp 1666464484
transform 1 0 24748 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_267
timestamp 1666464484
transform 1 0 25668 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_275
timestamp 1666464484
transform 1 0 26404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_283
timestamp 1666464484
transform 1 0 27140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_287
timestamp 1666464484
transform 1 0 27508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_290
timestamp 1666464484
transform 1 0 27784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1666464484
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1666464484
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1666464484
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1666464484
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1666464484
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_245
timestamp 1666464484
transform 1 0 23644 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_248
timestamp 1666464484
transform 1 0 23920 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_256
timestamp 1666464484
transform 1 0 24656 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1666464484
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_271
timestamp 1666464484
transform 1 0 26036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1666464484
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_285
timestamp 1666464484
transform 1 0 27324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_291
timestamp 1666464484
transform 1 0 27876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_297
timestamp 1666464484
transform 1 0 28428 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_229
timestamp 1666464484
transform 1 0 22172 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1666464484
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1666464484
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666464484
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666464484
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_259
timestamp 1666464484
transform 1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1666464484
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_275
timestamp 1666464484
transform 1 0 26404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_281
timestamp 1666464484
transform 1 0 26956 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1666464484
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_229
timestamp 1666464484
transform 1 0 22172 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_235
timestamp 1666464484
transform 1 0 22724 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1666464484
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_244
timestamp 1666464484
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_250
timestamp 1666464484
transform 1 0 24104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_256
timestamp 1666464484
transform 1 0 24656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_262
timestamp 1666464484
transform 1 0 25208 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_270
timestamp 1666464484
transform 1 0 25944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666464484
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_287
timestamp 1666464484
transform 1 0 27508 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_290
timestamp 1666464484
transform 1 0 27784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1666464484
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_8
timestamp 1666464484
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1666464484
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1666464484
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1666464484
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_225
timestamp 1666464484
transform 1 0 21804 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_229
timestamp 1666464484
transform 1 0 22172 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_232
timestamp 1666464484
transform 1 0 22448 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_238
timestamp 1666464484
transform 1 0 23000 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_241
timestamp 1666464484
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1666464484
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_257
timestamp 1666464484
transform 1 0 24748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_263
timestamp 1666464484
transform 1 0 25300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_269
timestamp 1666464484
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_275
timestamp 1666464484
transform 1 0 26404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_281
timestamp 1666464484
transform 1 0 26956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1666464484
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_290
timestamp 1666464484
transform 1 0 27784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1666464484
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1666464484
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1666464484
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1666464484
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_201
timestamp 1666464484
transform 1 0 19596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1666464484
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_212
timestamp 1666464484
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1666464484
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1666464484
transform 1 0 22172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_233
timestamp 1666464484
transform 1 0 22540 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1666464484
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_242
timestamp 1666464484
transform 1 0 23368 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_248
timestamp 1666464484
transform 1 0 23920 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1666464484
transform 1 0 24472 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_260
timestamp 1666464484
transform 1 0 25024 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_266
timestamp 1666464484
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1666464484
transform 1 0 26128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1666464484
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_285
timestamp 1666464484
transform 1 0 27324 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1666464484
transform 1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_205
timestamp 1666464484
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1666464484
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 1666464484
transform 1 0 21068 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_223
timestamp 1666464484
transform 1 0 21620 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_229
timestamp 1666464484
transform 1 0 22172 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1666464484
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp 1666464484
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1666464484
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_257
timestamp 1666464484
transform 1 0 24748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_263
timestamp 1666464484
transform 1 0 25300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_269
timestamp 1666464484
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_275
timestamp 1666464484
transform 1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_279
timestamp 1666464484
transform 1 0 26772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_283
timestamp 1666464484
transform 1 0 27140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1666464484
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_8
timestamp 1666464484
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_20
timestamp 1666464484
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_32
timestamp 1666464484
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_44
timestamp 1666464484
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 1666464484
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_199
timestamp 1666464484
transform 1 0 19412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1666464484
transform 1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_219
timestamp 1666464484
transform 1 0 21252 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_233
timestamp 1666464484
transform 1 0 22540 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_242
timestamp 1666464484
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_249
timestamp 1666464484
transform 1 0 24012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1666464484
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1666464484
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_268
timestamp 1666464484
transform 1 0 25760 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_274
timestamp 1666464484
transform 1 0 26312 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1666464484
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_286
timestamp 1666464484
transform 1 0 27416 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_182
timestamp 1666464484
transform 1 0 17848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_188
timestamp 1666464484
transform 1 0 18400 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_203
timestamp 1666464484
transform 1 0 19780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1666464484
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_239
timestamp 1666464484
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1666464484
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_258
timestamp 1666464484
transform 1 0 24840 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_269
timestamp 1666464484
transform 1 0 25852 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_276
timestamp 1666464484
transform 1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_283
timestamp 1666464484
transform 1 0 27140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_290
timestamp 1666464484
transform 1 0 27784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1666464484
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1666464484
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1666464484
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_32
timestamp 1666464484
transform 1 0 4048 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_44
timestamp 1666464484
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1666464484
transform 1 0 17020 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1666464484
transform 1 0 17572 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_185
timestamp 1666464484
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_196
timestamp 1666464484
transform 1 0 19136 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1666464484
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1666464484
transform 1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1666464484
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_234
timestamp 1666464484
transform 1 0 22632 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_245
timestamp 1666464484
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_254
timestamp 1666464484
transform 1 0 24472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_263
timestamp 1666464484
transform 1 0 25300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_271
timestamp 1666464484
transform 1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1666464484
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_290
timestamp 1666464484
transform 1 0 27784 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_297
timestamp 1666464484
transform 1 0 28428 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_161
timestamp 1666464484
transform 1 0 15916 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1666464484
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1666464484
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1666464484
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_214
timestamp 1666464484
transform 1 0 20792 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_225
timestamp 1666464484
transform 1 0 21804 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666464484
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666464484
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_260
timestamp 1666464484
transform 1 0 25024 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_269
timestamp 1666464484
transform 1 0 25852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_276
timestamp 1666464484
transform 1 0 26496 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_283
timestamp 1666464484
transform 1 0 27140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_290
timestamp 1666464484
transform 1 0 27784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1666464484
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_8
timestamp 1666464484
transform 1 0 1840 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_20
timestamp 1666464484
transform 1 0 2944 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_32
timestamp 1666464484
transform 1 0 4048 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_44
timestamp 1666464484
transform 1 0 5152 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1666464484
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_160
timestamp 1666464484
transform 1 0 15824 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1666464484
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1666464484
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_176
timestamp 1666464484
transform 1 0 17296 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_184
timestamp 1666464484
transform 1 0 18032 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_192
timestamp 1666464484
transform 1 0 18768 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_201
timestamp 1666464484
transform 1 0 19596 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_211
timestamp 1666464484
transform 1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1666464484
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_243
timestamp 1666464484
transform 1 0 23460 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_263
timestamp 1666464484
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_272
timestamp 1666464484
transform 1 0 26128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1666464484
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_290
timestamp 1666464484
transform 1 0 27784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_297
timestamp 1666464484
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1666464484
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1666464484
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1666464484
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_150
timestamp 1666464484
transform 1 0 14904 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_156
timestamp 1666464484
transform 1 0 15456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_162
timestamp 1666464484
transform 1 0 16008 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_168
timestamp 1666464484
transform 1 0 16560 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_174
timestamp 1666464484
transform 1 0 17112 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1666464484
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_204
timestamp 1666464484
transform 1 0 19872 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1666464484
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_235
timestamp 1666464484
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1666464484
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1666464484
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_280
timestamp 1666464484
transform 1 0 26864 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_288
timestamp 1666464484
transform 1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_292
timestamp 1666464484
transform 1 0 27968 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp 1666464484
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1666464484
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_141
timestamp 1666464484
transform 1 0 14076 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_147
timestamp 1666464484
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_153
timestamp 1666464484
transform 1 0 15180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_159
timestamp 1666464484
transform 1 0 15732 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_163
timestamp 1666464484
transform 1 0 16100 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1666464484
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_175
timestamp 1666464484
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_191
timestamp 1666464484
transform 1 0 18676 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1666464484
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_243
timestamp 1666464484
transform 1 0 23460 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_263
timestamp 1666464484
transform 1 0 25300 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1666464484
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_288
timestamp 1666464484
transform 1 0 27600 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_296
timestamp 1666464484
transform 1 0 28336 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1666464484
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_129
timestamp 1666464484
transform 1 0 12972 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_132
timestamp 1666464484
transform 1 0 13248 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1666464484
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_149
timestamp 1666464484
transform 1 0 14812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_155
timestamp 1666464484
transform 1 0 15364 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_163
timestamp 1666464484
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_172
timestamp 1666464484
transform 1 0 16928 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_183
timestamp 1666464484
transform 1 0 17940 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1666464484
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_215
timestamp 1666464484
transform 1 0 20884 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_235
timestamp 1666464484
transform 1 0 22724 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_246
timestamp 1666464484
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1666464484
transform 1 0 26036 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_282
timestamp 1666464484
transform 1 0 27048 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_292
timestamp 1666464484
transform 1 0 27968 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_298
timestamp 1666464484
transform 1 0 28520 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_8
timestamp 1666464484
transform 1 0 1840 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_20
timestamp 1666464484
transform 1 0 2944 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_32
timestamp 1666464484
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_44
timestamp 1666464484
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_103
timestamp 1666464484
transform 1 0 10580 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_107
timestamp 1666464484
transform 1 0 10948 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1666464484
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_119
timestamp 1666464484
transform 1 0 12052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_131
timestamp 1666464484
transform 1 0 13156 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1666464484
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_157
timestamp 1666464484
transform 1 0 15548 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1666464484
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1666464484
transform 1 0 17848 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1666464484
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1666464484
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_243
timestamp 1666464484
transform 1 0 23460 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_263
timestamp 1666464484
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1666464484
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_290
timestamp 1666464484
transform 1 0 27784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1666464484
transform 1 0 28428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1666464484
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1666464484
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_93
timestamp 1666464484
transform 1 0 9660 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_96
timestamp 1666464484
transform 1 0 9936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1666464484
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_108
timestamp 1666464484
transform 1 0 11040 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1666464484
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_120
timestamp 1666464484
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1666464484
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_132
timestamp 1666464484
transform 1 0 13248 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1666464484
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_152
timestamp 1666464484
transform 1 0 15088 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_163
timestamp 1666464484
transform 1 0 16100 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_174
timestamp 1666464484
transform 1 0 17112 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_216
timestamp 1666464484
transform 1 0 20976 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_236
timestamp 1666464484
transform 1 0 22816 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1666464484
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_271
timestamp 1666464484
transform 1 0 26036 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_291
timestamp 1666464484
transform 1 0 27876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1666464484
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1666464484
transform 1 0 9016 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_92
timestamp 1666464484
transform 1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_98
timestamp 1666464484
transform 1 0 10120 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_104
timestamp 1666464484
transform 1 0 10672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1666464484
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_119
timestamp 1666464484
transform 1 0 12052 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_122
timestamp 1666464484
transform 1 0 12328 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_128
timestamp 1666464484
transform 1 0 12880 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1666464484
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_145
timestamp 1666464484
transform 1 0 14444 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_155
timestamp 1666464484
transform 1 0 15364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1666464484
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_182
timestamp 1666464484
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_202
timestamp 1666464484
transform 1 0 19688 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1666464484
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_243
timestamp 1666464484
transform 1 0 23460 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_263
timestamp 1666464484
transform 1 0 25300 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1666464484
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_290
timestamp 1666464484
transform 1 0 27784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1666464484
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_73
timestamp 1666464484
transform 1 0 7820 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_76
timestamp 1666464484
transform 1 0 8096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1666464484
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_91
timestamp 1666464484
transform 1 0 9476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_103
timestamp 1666464484
transform 1 0 10580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_115
timestamp 1666464484
transform 1 0 11684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_129
timestamp 1666464484
transform 1 0 12972 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1666464484
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_154
timestamp 1666464484
transform 1 0 15272 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1666464484
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1666464484
transform 1 0 19596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1666464484
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1666464484
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1666464484
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_291
timestamp 1666464484
transform 1 0 27876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1666464484
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1666464484
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1666464484
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1666464484
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1666464484
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_65
timestamp 1666464484
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_68
timestamp 1666464484
transform 1 0 7360 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_74
timestamp 1666464484
transform 1 0 7912 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_80
timestamp 1666464484
transform 1 0 8464 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_86
timestamp 1666464484
transform 1 0 9016 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1666464484
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_98
timestamp 1666464484
transform 1 0 10120 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_104
timestamp 1666464484
transform 1 0 10672 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1666464484
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_119
timestamp 1666464484
transform 1 0 12052 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_135
timestamp 1666464484
transform 1 0 13524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_146
timestamp 1666464484
transform 1 0 14536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1666464484
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_173
timestamp 1666464484
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_182
timestamp 1666464484
transform 1 0 17848 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_202
timestamp 1666464484
transform 1 0 19688 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1666464484
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1666464484
transform 1 0 23460 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_263
timestamp 1666464484
transform 1 0 25300 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1666464484
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_290
timestamp 1666464484
transform 1 0 27784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_297
timestamp 1666464484
transform 1 0 28428 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_8
timestamp 1666464484
transform 1 0 1840 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1666464484
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_58
timestamp 1666464484
transform 1 0 6440 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_64
timestamp 1666464484
transform 1 0 6992 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_70
timestamp 1666464484
transform 1 0 7544 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_76
timestamp 1666464484
transform 1 0 8096 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1666464484
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_91
timestamp 1666464484
transform 1 0 9476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_94
timestamp 1666464484
transform 1 0 9752 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_100
timestamp 1666464484
transform 1 0 10304 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_108
timestamp 1666464484
transform 1 0 11040 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_117
timestamp 1666464484
transform 1 0 11868 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_127
timestamp 1666464484
transform 1 0 12788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1666464484
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_154
timestamp 1666464484
transform 1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_174
timestamp 1666464484
transform 1 0 17112 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_212
timestamp 1666464484
transform 1 0 20608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1666464484
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1666464484
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1666464484
transform 1 0 26036 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_291
timestamp 1666464484
transform 1 0 27876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_297
timestamp 1666464484
transform 1 0 28428 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1666464484
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_63
timestamp 1666464484
transform 1 0 6900 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_75
timestamp 1666464484
transform 1 0 8004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_87
timestamp 1666464484
transform 1 0 9108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_101
timestamp 1666464484
transform 1 0 10396 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1666464484
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_126
timestamp 1666464484
transform 1 0 12696 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1666464484
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1666464484
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_173
timestamp 1666464484
transform 1 0 17020 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_182
timestamp 1666464484
transform 1 0 17848 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1666464484
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1666464484
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_243
timestamp 1666464484
transform 1 0 23460 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_263
timestamp 1666464484
transform 1 0 25300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp 1666464484
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_291
timestamp 1666464484
transform 1 0 27876 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_297
timestamp 1666464484
transform 1 0 28428 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_8
timestamp 1666464484
transform 1 0 1840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1666464484
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_37
timestamp 1666464484
transform 1 0 4508 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_40
timestamp 1666464484
transform 1 0 4784 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_46
timestamp 1666464484
transform 1 0 5336 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_52
timestamp 1666464484
transform 1 0 5888 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_58
timestamp 1666464484
transform 1 0 6440 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_64
timestamp 1666464484
transform 1 0 6992 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_70
timestamp 1666464484
transform 1 0 7544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_76
timestamp 1666464484
transform 1 0 8096 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1666464484
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 1666464484
transform 1 0 9476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_107
timestamp 1666464484
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_118
timestamp 1666464484
transform 1 0 11960 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1666464484
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_154
timestamp 1666464484
transform 1 0 15272 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_174
timestamp 1666464484
transform 1 0 17112 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1666464484
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_201
timestamp 1666464484
transform 1 0 19596 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_212
timestamp 1666464484
transform 1 0 20608 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_232
timestamp 1666464484
transform 1 0 22448 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1666464484
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_271
timestamp 1666464484
transform 1 0 26036 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_291
timestamp 1666464484
transform 1 0 27876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1666464484
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_33
timestamp 1666464484
transform 1 0 4140 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_36
timestamp 1666464484
transform 1 0 4416 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_42
timestamp 1666464484
transform 1 0 4968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_48
timestamp 1666464484
transform 1 0 5520 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1666464484
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_61
timestamp 1666464484
transform 1 0 6716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_67
timestamp 1666464484
transform 1 0 7268 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_73
timestamp 1666464484
transform 1 0 7820 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_79
timestamp 1666464484
transform 1 0 8372 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_86
timestamp 1666464484
transform 1 0 9016 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_101
timestamp 1666464484
transform 1 0 10396 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1666464484
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_126
timestamp 1666464484
transform 1 0 12696 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_146
timestamp 1666464484
transform 1 0 14536 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1666464484
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1666464484
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_182
timestamp 1666464484
transform 1 0 17848 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_202
timestamp 1666464484
transform 1 0 19688 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1666464484
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_243
timestamp 1666464484
transform 1 0 23460 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_263
timestamp 1666464484
transform 1 0 25300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1666464484
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_291
timestamp 1666464484
transform 1 0 27876 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1666464484
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1666464484
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_20
timestamp 1666464484
transform 1 0 2944 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1666464484
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_33
timestamp 1666464484
transform 1 0 4140 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_39
timestamp 1666464484
transform 1 0 4692 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_45
timestamp 1666464484
transform 1 0 5244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_51
timestamp 1666464484
transform 1 0 5796 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_57
timestamp 1666464484
transform 1 0 6348 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_63
timestamp 1666464484
transform 1 0 6900 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_69
timestamp 1666464484
transform 1 0 7452 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_75
timestamp 1666464484
transform 1 0 8004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1666464484
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_92
timestamp 1666464484
transform 1 0 9568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_100
timestamp 1666464484
transform 1 0 10304 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_108
timestamp 1666464484
transform 1 0 11040 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_117
timestamp 1666464484
transform 1 0 11868 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_127
timestamp 1666464484
transform 1 0 12788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1666464484
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_154
timestamp 1666464484
transform 1 0 15272 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_174
timestamp 1666464484
transform 1 0 17112 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_201
timestamp 1666464484
transform 1 0 19596 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_213
timestamp 1666464484
transform 1 0 20700 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_233
timestamp 1666464484
transform 1 0 22540 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1666464484
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_271
timestamp 1666464484
transform 1 0 26036 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1666464484
transform 1 0 27876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_297
timestamp 1666464484
transform 1 0 28428 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_11
timestamp 1666464484
transform 1 0 2116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_18
timestamp 1666464484
transform 1 0 2760 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_26
timestamp 1666464484
transform 1 0 3496 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_29
timestamp 1666464484
transform 1 0 3772 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_34
timestamp 1666464484
transform 1 0 4232 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_42
timestamp 1666464484
transform 1 0 4968 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_47
timestamp 1666464484
transform 1 0 5428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1666464484
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_61
timestamp 1666464484
transform 1 0 6716 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_68
timestamp 1666464484
transform 1 0 7360 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_75
timestamp 1666464484
transform 1 0 8004 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_82
timestamp 1666464484
transform 1 0 8648 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_85
timestamp 1666464484
transform 1 0 8924 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_91
timestamp 1666464484
transform 1 0 9476 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_97
timestamp 1666464484
transform 1 0 10028 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_102
timestamp 1666464484
transform 1 0 10488 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1666464484
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_119
timestamp 1666464484
transform 1 0 12052 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_128
timestamp 1666464484
transform 1 0 12880 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_138
timestamp 1666464484
transform 1 0 13800 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_141
timestamp 1666464484
transform 1 0 14076 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_146
timestamp 1666464484
transform 1 0 14536 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1666464484
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_174
timestamp 1666464484
transform 1 0 17112 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_194
timestamp 1666464484
transform 1 0 18952 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_197
timestamp 1666464484
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_202
timestamp 1666464484
transform 1 0 19688 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1666464484
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_243
timestamp 1666464484
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_250
timestamp 1666464484
transform 1 0 24104 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_253
timestamp 1666464484
transform 1 0 24380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_271
timestamp 1666464484
transform 1 0 26036 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1666464484
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_290
timestamp 1666464484
transform 1 0 27784 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1666464484
transform 1 0 28428 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 28888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 28888 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 28888 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 28888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 28888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 28888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 3680 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 8832 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 13984 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 19136 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 24288 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _094_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27968 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _095_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1666464484
transform -1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _097_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19780 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _098_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18768 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _099_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26128 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _101_
timestamp 1666464484
transform 1 0 28152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1666464484
transform -1 0 10396 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _103_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26496 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23000 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1666464484
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26588 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 1666464484
transform -1 0 23828 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _108_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27600 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19044 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1666464484
transform 1 0 10028 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27416 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1666464484
transform 1 0 10672 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 1666464484
transform 1 0 22908 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1666464484
transform 1 0 22816 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _115_
timestamp 1666464484
transform 1 0 9568 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _116_
timestamp 1666464484
transform -1 0 27048 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1666464484
transform -1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1666464484
transform -1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _119_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12788 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _120_
timestamp 1666464484
transform 1 0 25668 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _121_
timestamp 1666464484
transform -1 0 20608 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _122_
timestamp 1666464484
transform -1 0 19596 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1666464484
transform 1 0 23736 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _124_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26496 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _125_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _126_
timestamp 1666464484
transform -1 0 22540 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _127_
timestamp 1666464484
transform 1 0 20884 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _128_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _129_
timestamp 1666464484
transform 1 0 11408 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _130_
timestamp 1666464484
transform -1 0 13800 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _131_
timestamp 1666464484
transform -1 0 20700 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _132_
timestamp 1666464484
transform -1 0 16100 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _133_
timestamp 1666464484
transform -1 0 19964 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _134_
timestamp 1666464484
transform 1 0 11316 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _135_
timestamp 1666464484
transform -1 0 10948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _136_
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _137_
timestamp 1666464484
transform 1 0 25668 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _138_
timestamp 1666464484
transform 1 0 23184 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _139_
timestamp 1666464484
transform -1 0 14444 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _140_
timestamp 1666464484
transform 1 0 12052 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _141_
timestamp 1666464484
transform -1 0 23920 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _142_
timestamp 1666464484
transform 1 0 17296 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _143_
timestamp 1666464484
transform 1 0 24564 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _144_
timestamp 1666464484
transform -1 0 27784 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _145_
timestamp 1666464484
transform -1 0 20516 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _146_
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _147_
timestamp 1666464484
transform -1 0 15272 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _148_
timestamp 1666464484
transform 1 0 17112 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _149_
timestamp 1666464484
transform -1 0 25300 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _150_
timestamp 1666464484
transform 1 0 17204 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _151_
timestamp 1666464484
transform 1 0 26404 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _152_
timestamp 1666464484
transform 1 0 27140 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _153_
timestamp 1666464484
transform -1 0 16376 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _154_
timestamp 1666464484
transform 1 0 14628 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _155_
timestamp 1666464484
transform -1 0 13524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _156_
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _157_
timestamp 1666464484
transform 1 0 25668 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _158_
timestamp 1666464484
transform 1 0 17112 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _159_
timestamp 1666464484
transform -1 0 23368 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _160_
timestamp 1666464484
transform 1 0 18308 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _161_
timestamp 1666464484
transform 1 0 12420 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _162_
timestamp 1666464484
transform -1 0 14536 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _163_
timestamp 1666464484
transform -1 0 17756 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _164_
timestamp 1666464484
transform 1 0 14628 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _165_
timestamp 1666464484
transform -1 0 18676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _166_
timestamp 1666464484
transform 1 0 22632 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _167_
timestamp 1666464484
transform 1 0 27140 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _168_
timestamp 1666464484
transform -1 0 20700 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _169_
timestamp 1666464484
transform 1 0 14628 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _170_
timestamp 1666464484
transform -1 0 17112 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1666464484
transform -1 0 18124 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _172_
timestamp 1666464484
transform 1 0 12052 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _173_
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _174_
timestamp 1666464484
transform -1 0 23736 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _175_
timestamp 1666464484
transform -1 0 13800 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _176_
timestamp 1666464484
transform 1 0 19412 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _177_
timestamp 1666464484
transform 1 0 23092 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _178_
timestamp 1666464484
transform 1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _179_
timestamp 1666464484
transform 1 0 11408 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _180_
timestamp 1666464484
transform -1 0 22632 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 1666464484
transform 1 0 25392 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _182_
timestamp 1666464484
transform -1 0 26312 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _183_
timestamp 1666464484
transform -1 0 16928 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _184_
timestamp 1666464484
transform 1 0 13156 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _185_
timestamp 1666464484
transform -1 0 15364 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _186_
timestamp 1666464484
transform -1 0 22264 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _187_
timestamp 1666464484
transform -1 0 17848 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _188_
timestamp 1666464484
transform 1 0 27140 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _189_
timestamp 1666464484
transform 1 0 12144 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _190_
timestamp 1666464484
transform 1 0 20240 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _191_
timestamp 1666464484
transform -1 0 24472 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _192_
timestamp 1666464484
transform 1 0 21160 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _193_
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _194_
timestamp 1666464484
transform -1 0 15272 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _195_
timestamp 1666464484
transform -1 0 12788 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _196_
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _197_
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _198_
timestamp 1666464484
transform -1 0 17848 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _199_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26404 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _200_
timestamp 1666464484
transform -1 0 23460 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _201_
timestamp 1666464484
transform 1 0 24564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _202_
timestamp 1666464484
transform 1 0 18216 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _203_
timestamp 1666464484
transform 1 0 20056 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _204_
timestamp 1666464484
transform 1 0 17480 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _205_
timestamp 1666464484
transform 1 0 14904 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _206_
timestamp 1666464484
transform -1 0 16376 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _207_
timestamp 1666464484
transform 1 0 17480 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _208_
timestamp 1666464484
transform 1 0 21988 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _209_
timestamp 1666464484
transform 1 0 24564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _210_
timestamp 1666464484
transform -1 0 26036 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _211_
timestamp 1666464484
transform -1 0 17112 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _212_
timestamp 1666464484
transform -1 0 18952 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _213_
timestamp 1666464484
transform 1 0 23828 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1666464484
transform 1 0 18216 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1666464484
transform 1 0 21988 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1666464484
transform -1 0 21528 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1666464484
transform 1 0 21988 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1666464484
transform -1 0 25300 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1666464484
transform -1 0 17112 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1666464484
transform -1 0 18952 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1666464484
transform -1 0 26036 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp 1666464484
transform -1 0 26036 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _223_
timestamp 1666464484
transform -1 0 23644 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1666464484
transform -1 0 26036 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _225_
timestamp 1666464484
transform -1 0 23460 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _226_
timestamp 1666464484
transform 1 0 14904 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _227_
timestamp 1666464484
transform 1 0 15640 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _228_
timestamp 1666464484
transform -1 0 21528 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _229_
timestamp 1666464484
transform 1 0 24564 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _230_
timestamp 1666464484
transform -1 0 25300 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _231_
timestamp 1666464484
transform -1 0 19688 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1666464484
transform 1 0 20056 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1666464484
transform 1 0 21988 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1666464484
transform 1 0 24564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1666464484
transform 1 0 23828 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _236_
timestamp 1666464484
transform -1 0 21528 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _237_
timestamp 1666464484
transform -1 0 22540 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1666464484
transform -1 0 18952 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1666464484
transform 1 0 18216 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1666464484
transform -1 0 22448 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _241_
timestamp 1666464484
transform 1 0 21068 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp 1666464484
transform -1 0 22724 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _243_
timestamp 1666464484
transform -1 0 27876 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _244_
timestamp 1666464484
transform -1 0 22448 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _245_
timestamp 1666464484
transform -1 0 23460 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _246_
timestamp 1666464484
transform -1 0 25300 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _247_
timestamp 1666464484
transform 1 0 20056 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _248_
timestamp 1666464484
transform -1 0 23460 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _249_
timestamp 1666464484
transform 1 0 23828 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _250_
timestamp 1666464484
transform -1 0 16376 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _251_
timestamp 1666464484
transform -1 0 27876 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _252_
timestamp 1666464484
transform -1 0 22816 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _253_
timestamp 1666464484
transform 1 0 17480 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _254_
timestamp 1666464484
transform -1 0 21528 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _255_
timestamp 1666464484
transform 1 0 21252 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _256_
timestamp 1666464484
transform -1 0 25300 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _257_
timestamp 1666464484
transform 1 0 26404 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _258_
timestamp 1666464484
transform 1 0 13064 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _259_
timestamp 1666464484
transform -1 0 19688 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _260_
timestamp 1666464484
transform -1 0 20884 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _261_
timestamp 1666464484
transform 1 0 15640 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _262_
timestamp 1666464484
transform 1 0 13064 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _263_
timestamp 1666464484
transform 1 0 26404 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _264_
timestamp 1666464484
transform 1 0 12328 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _265_
timestamp 1666464484
transform 1 0 19504 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _334_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1666464484
transform -1 0 8648 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1666464484
transform 1 0 28152 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp 1666464484
transform 1 0 26404 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1666464484
transform 1 0 16836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1666464484
transform 1 0 14260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp 1666464484
transform 1 0 19412 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1666464484
transform 1 0 9292 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1666464484
transform -1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout17
timestamp 1666464484
transform -1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1666464484
transform 1 0 15180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout19
timestamp 1666464484
transform 1 0 22816 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1666464484
transform 1 0 12604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1666464484
transform 1 0 10672 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout22
timestamp 1666464484
transform 1 0 28152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout23
timestamp 1666464484
transform -1 0 9660 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1666464484
transform 1 0 28152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform 1 0 27508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform 1 0 27508 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform -1 0 28428 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1666464484
transform -1 0 28428 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform 1 0 28152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform 1 0 9936 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform -1 0 11224 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform -1 0 12052 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform -1 0 10488 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform -1 0 9476 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1666464484
transform -1 0 5428 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1666464484
transform -1 0 2116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_24 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_25
timestamp 1666464484
transform 1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_26
timestamp 1666464484
transform 1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_27
timestamp 1666464484
transform 1 0 28152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_28
timestamp 1666464484
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_29
timestamp 1666464484
transform 1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_30
timestamp 1666464484
transform 1 0 28152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_31
timestamp 1666464484
transform 1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_32
timestamp 1666464484
transform 1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_33
timestamp 1666464484
transform 1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_34
timestamp 1666464484
transform 1 0 28152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_35
timestamp 1666464484
transform 1 0 27508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_36
timestamp 1666464484
transform 1 0 26404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_37
timestamp 1666464484
transform 1 0 28152 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_38
timestamp 1666464484
transform 1 0 26864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_39
timestamp 1666464484
transform 1 0 27508 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_40
timestamp 1666464484
transform -1 0 1840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_41
timestamp 1666464484
transform -1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_42
timestamp 1666464484
transform -1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_43
timestamp 1666464484
transform -1 0 1840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_44
timestamp 1666464484
transform -1 0 1840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_45
timestamp 1666464484
transform -1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_46
timestamp 1666464484
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_47
timestamp 1666464484
transform -1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_48
timestamp 1666464484
transform -1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_49
timestamp 1666464484
transform -1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_50
timestamp 1666464484
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_51
timestamp 1666464484
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_52
timestamp 1666464484
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_53
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_54
timestamp 1666464484
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_55
timestamp 1666464484
transform 1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_56
timestamp 1666464484
transform 1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_57
timestamp 1666464484
transform 1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_58
timestamp 1666464484
transform 1 0 28152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_59
timestamp 1666464484
transform 1 0 28152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_60
timestamp 1666464484
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_61
timestamp 1666464484
transform 1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_62
timestamp 1666464484
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_63
timestamp 1666464484
transform 1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_64
timestamp 1666464484
transform 1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_65
timestamp 1666464484
transform 1 0 27508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_66
timestamp 1666464484
transform 1 0 26864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_67
timestamp 1666464484
transform 1 0 26220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_68
timestamp 1666464484
transform 1 0 25576 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_69
timestamp 1666464484
transform -1 0 27416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_70
timestamp 1666464484
transform -1 0 24656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_71
timestamp 1666464484
transform 1 0 7728 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_72
timestamp 1666464484
transform -1 0 24104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_73
timestamp 1666464484
transform 1 0 8372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_74
timestamp 1666464484
transform 1 0 8740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_75
timestamp 1666464484
transform -1 0 7360 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_76
timestamp 1666464484
transform -1 0 4232 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_77
timestamp 1666464484
transform -1 0 2760 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_78
timestamp 1666464484
transform -1 0 1840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_79
timestamp 1666464484
transform -1 0 1840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_80
timestamp 1666464484
transform -1 0 1840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_81
timestamp 1666464484
transform -1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_82
timestamp 1666464484
transform -1 0 1840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_83
timestamp 1666464484
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_84
timestamp 1666464484
transform -1 0 1840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_85
timestamp 1666464484
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_86
timestamp 1666464484
transform -1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_87
timestamp 1666464484
transform -1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_88
timestamp 1666464484
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_89
timestamp 1666464484
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_90
timestamp 1666464484
transform -1 0 1840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tiny_user_project_91
timestamp 1666464484
transform -1 0 1840 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal3 s 29200 1912 30000 2032 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 29200 22312 30000 22432 0 FreeSans 480 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 29200 24352 30000 24472 0 FreeSans 480 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 29200 26392 30000 26512 0 FreeSans 480 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 29200 28432 30000 28552 0 FreeSans 480 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 29200 30472 30000 30592 0 FreeSans 480 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 29274 33200 29330 34000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 25962 33200 26018 34000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 22650 33200 22706 34000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 19338 33200 19394 34000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 16026 33200 16082 34000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 29200 3952 30000 4072 0 FreeSans 480 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 12714 33200 12770 34000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 9402 33200 9458 34000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 6090 33200 6146 34000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 2778 33200 2834 34000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 29200 5992 30000 6112 0 FreeSans 480 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 29200 8032 30000 8152 0 FreeSans 480 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 29200 10072 30000 10192 0 FreeSans 480 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 29200 12112 30000 12232 0 FreeSans 480 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 29200 14152 30000 14272 0 FreeSans 480 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 29200 16192 30000 16312 0 FreeSans 480 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 29200 18232 30000 18352 0 FreeSans 480 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 29200 20272 30000 20392 0 FreeSans 480 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 29200 3272 30000 3392 0 FreeSans 480 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 29200 23672 30000 23792 0 FreeSans 480 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 29200 25712 30000 25832 0 FreeSans 480 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 29200 27752 30000 27872 0 FreeSans 480 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 29200 29792 30000 29912 0 FreeSans 480 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 29200 31832 30000 31952 0 FreeSans 480 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 27066 33200 27122 34000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 23754 33200 23810 34000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 20442 33200 20498 34000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 17130 33200 17186 34000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 13818 33200 13874 34000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 29200 5312 30000 5432 0 FreeSans 480 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 10506 33200 10562 34000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 7194 33200 7250 34000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 3882 33200 3938 34000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 570 33200 626 34000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 29200 7352 30000 7472 0 FreeSans 480 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 29200 9392 30000 9512 0 FreeSans 480 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 29200 11432 30000 11552 0 FreeSans 480 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 29200 13472 30000 13592 0 FreeSans 480 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 29200 15512 30000 15632 0 FreeSans 480 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 29200 17552 30000 17672 0 FreeSans 480 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 29200 19592 30000 19712 0 FreeSans 480 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 29200 21632 30000 21752 0 FreeSans 480 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 29200 2592 30000 2712 0 FreeSans 480 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 29200 22992 30000 23112 0 FreeSans 480 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 29200 25032 30000 25152 0 FreeSans 480 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 29200 27072 30000 27192 0 FreeSans 480 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 29200 29112 30000 29232 0 FreeSans 480 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 29200 31152 30000 31272 0 FreeSans 480 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 28170 33200 28226 34000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 24858 33200 24914 34000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 21546 33200 21602 34000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 18234 33200 18290 34000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 14922 33200 14978 34000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 29200 4632 30000 4752 0 FreeSans 480 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 11610 33200 11666 34000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 8298 33200 8354 34000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 4986 33200 5042 34000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 1674 33200 1730 34000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 0 28160 800 28280 0 FreeSans 480 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s 0 24080 800 24200 0 FreeSans 480 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 29200 6672 30000 6792 0 FreeSans 480 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 29200 8712 30000 8832 0 FreeSans 480 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 29200 10752 30000 10872 0 FreeSans 480 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 29200 12792 30000 12912 0 FreeSans 480 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 29200 14832 30000 14952 0 FreeSans 480 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 29200 16872 30000 16992 0 FreeSans 480 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 29200 18912 30000 19032 0 FreeSans 480 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 29200 20952 30000 21072 0 FreeSans 480 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4417 2128 4737 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 11363 2128 11683 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 18309 2128 18629 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 25255 2128 25575 31600 0 FreeSans 1920 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 7890 2128 8210 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 31600 0 FreeSans 1920 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 14996 31008 14996 31008 0 vccd1
rlabel via1 15076 31552 15076 31552 0 vssd1
rlabel metal1 5014 30362 5014 30362 0 _000_
rlabel metal2 14214 24684 14214 24684 0 _001_
rlabel metal1 15318 23766 15318 23766 0 _002_
rlabel metal2 16790 23800 16790 23800 0 _003_
rlabel via2 17250 25245 17250 25245 0 _004_
rlabel metal1 27186 30226 27186 30226 0 _005_
rlabel metal1 14950 26928 14950 26928 0 _006_
rlabel metal1 16284 23290 16284 23290 0 _007_
rlabel metal2 13662 28764 13662 28764 0 _008_
rlabel metal1 10810 30022 10810 30022 0 _009_
rlabel metal2 19872 29036 19872 29036 0 _010_
rlabel metal1 18357 23562 18357 23562 0 _011_
rlabel metal1 23644 25262 23644 25262 0 _012_
rlabel metal1 16422 27098 16422 27098 0 _013_
rlabel metal1 21804 21658 21804 21658 0 _014_
rlabel metal1 21298 23562 21298 23562 0 _015_
rlabel metal2 13202 29716 13202 29716 0 _016_
rlabel metal4 23460 29240 23460 29240 0 _017_
rlabel metal1 17894 22474 17894 22474 0 _018_
rlabel metal2 23414 26452 23414 26452 0 _019_
rlabel metal2 19550 23001 19550 23001 0 _020_
rlabel via2 11362 29699 11362 29699 0 _021_
rlabel metal3 18860 25704 18860 25704 0 _022_
rlabel metal1 21804 22746 21804 22746 0 _023_
rlabel metal2 23874 26180 23874 26180 0 _024_
rlabel metal1 13340 27098 13340 27098 0 _025_
rlabel metal1 15456 28934 15456 28934 0 _026_
rlabel metal1 23460 22134 23460 22134 0 _027_
rlabel metal1 17296 25398 17296 25398 0 _028_
rlabel metal2 26634 30362 26634 30362 0 _029_
rlabel metal1 23782 31144 23782 31144 0 _030_
rlabel metal2 20286 23919 20286 23919 0 _031_
rlabel metal1 12098 29002 12098 29002 0 _032_
rlabel metal1 17388 29070 17388 29070 0 _033_
rlabel metal1 20369 22508 20369 22508 0 _034_
rlabel metal1 17020 25942 17020 25942 0 _035_
rlabel metal1 27278 25806 27278 25806 0 _036_
rlabel metal3 19780 25840 19780 25840 0 _037_
rlabel metal1 15594 26010 15594 26010 0 _038_
rlabel metal1 16159 30294 16159 30294 0 _039_
rlabel via2 13294 27965 13294 27965 0 _040_
rlabel metal3 18860 30056 18860 30056 0 _041_
rlabel metal2 19458 29903 19458 29903 0 _042_
rlabel metal2 18722 21835 18722 21835 0 _043_
rlabel metal2 20378 30804 20378 30804 0 _044_
rlabel metal1 13846 28050 13846 28050 0 _045_
rlabel metal1 16100 28186 16100 28186 0 _046_
rlabel metal1 16376 24650 16376 24650 0 _047_
rlabel metal1 17388 28730 17388 28730 0 _048_
rlabel via2 18538 24701 18538 24701 0 _049_
rlabel metal2 23046 22151 23046 22151 0 _050_
rlabel metal1 23046 28084 23046 28084 0 _051_
rlabel metal1 16514 26384 16514 26384 0 _052_
rlabel metal1 17112 26486 17112 26486 0 _053_
rlabel metal2 14306 26962 14306 26962 0 _054_
rlabel metal2 20194 27489 20194 27489 0 _055_
rlabel metal1 21390 24208 21390 24208 0 _056_
rlabel metal1 23644 24378 23644 24378 0 _057_
rlabel metal3 18423 31756 18423 31756 0 _058_
rlabel metal1 21482 24378 21482 24378 0 _059_
rlabel via1 20746 25211 20746 25211 0 _060_
rlabel metal4 12052 26520 12052 26520 0 _061_
rlabel metal1 22448 22406 22448 22406 0 _062_
rlabel metal1 25760 23222 25760 23222 0 _063_
rlabel metal1 27278 29138 27278 29138 0 _064_
rlabel metal1 15134 25466 15134 25466 0 _065_
rlabel metal2 13294 28509 13294 28509 0 _066_
rlabel metal1 17526 26792 17526 26792 0 _067_
rlabel metal1 20792 21862 20792 21862 0 _068_
rlabel metal1 17848 27098 17848 27098 0 _069_
rlabel metal2 13110 26061 13110 26061 0 _070_
rlabel metal2 20286 26180 20286 26180 0 _071_
rlabel metal1 23276 22746 23276 22746 0 _072_
rlabel metal1 19412 23154 19412 23154 0 _073_
rlabel metal1 14214 27438 14214 27438 0 _074_
rlabel metal1 15640 27574 15640 27574 0 _075_
rlabel via2 12558 28509 12558 28509 0 _076_
rlabel metal1 21298 23290 21298 23290 0 _077_
rlabel metal1 22146 26996 22146 26996 0 _078_
rlabel metal3 20447 21556 20447 21556 0 _079_
rlabel metal1 19320 28390 19320 28390 0 _080_
rlabel metal4 23828 27404 23828 27404 0 _081_
rlabel metal1 22954 27506 22954 27506 0 _082_
rlabel metal1 22908 28526 22908 28526 0 _083_
rlabel metal1 9384 26758 9384 26758 0 _084_
rlabel metal2 12006 25534 12006 25534 0 _085_
rlabel metal1 26634 23222 26634 23222 0 _086_
rlabel metal1 23322 22678 23322 22678 0 _087_
rlabel metal1 22770 18598 22770 18598 0 _088_
rlabel metal1 11776 25738 11776 25738 0 _089_
rlabel metal2 6854 29002 6854 29002 0 _090_
rlabel metal2 23230 24361 23230 24361 0 _091_
rlabel via2 19090 24803 19090 24803 0 _092_
rlabel metal1 23552 24174 23552 24174 0 _093_
rlabel metal1 28336 22610 28336 22610 0 io_in[10]
rlabel metal1 27692 18394 27692 18394 0 io_in[11]
rlabel metal1 27370 20026 27370 20026 0 io_in[12]
rlabel metal1 27784 17850 27784 17850 0 io_in[13]
rlabel metal2 29348 31756 29348 31756 0 io_in[15]
rlabel via2 28382 18309 28382 18309 0 io_in[8]
rlabel metal2 28382 20383 28382 20383 0 io_in[9]
rlabel metal2 25392 33252 25392 33252 0 io_out[16]
rlabel metal1 16146 30872 16146 30872 0 io_out[17]
rlabel metal2 18262 32489 18262 32489 0 io_out[18]
rlabel metal2 11822 31824 11822 31824 0 io_out[19]
rlabel metal1 10948 31450 10948 31450 0 io_out[20]
rlabel metal1 8786 31450 8786 31450 0 io_out[21]
rlabel metal1 5106 31450 5106 31450 0 io_out[22]
rlabel metal1 1794 31450 1794 31450 0 io_out[23]
rlabel metal2 24886 21267 24886 21267 0 mod.flipflop1.d
rlabel metal1 23920 20910 23920 20910 0 mod.flipflop1.q
rlabel metal2 24610 30464 24610 30464 0 mod.flipflop10.d
rlabel metal1 19228 23086 19228 23086 0 mod.flipflop10.q
rlabel metal1 21804 27846 21804 27846 0 mod.flipflop11.d
rlabel metal1 16524 30226 16524 30226 0 mod.flipflop11.q
rlabel metal1 16698 27846 16698 27846 0 mod.flipflop12.d
rlabel metal2 13386 27319 13386 27319 0 mod.flipflop12.q
rlabel metal2 19182 24888 19182 24888 0 mod.flipflop13.d
rlabel metal3 22724 24344 22724 24344 0 mod.flipflop13.q
rlabel metal1 20792 26214 20792 26214 0 mod.flipflop14.d
rlabel metal1 18814 27472 18814 27472 0 mod.flipflop14.q
rlabel via1 23142 29138 23142 29138 0 mod.flipflop15.q
rlabel metal1 13478 28492 13478 28492 0 mod.flipflop16.q
rlabel via1 20373 26962 20373 26962 0 mod.flipflop17.q
rlabel metal1 22862 26758 22862 26758 0 mod.flipflop18.d
rlabel metal2 21114 27370 21114 27370 0 mod.flipflop18.q
rlabel metal1 11454 30600 11454 30600 0 mod.flipflop19.d
rlabel via2 14674 26299 14674 26299 0 mod.flipflop19.q
rlabel via1 22305 26962 22305 26962 0 mod.flipflop2.q
rlabel metal1 16897 27370 16897 27370 0 mod.flipflop20.d
rlabel metal1 13018 30226 13018 30226 0 mod.flipflop20.q
rlabel metal3 17273 29308 17273 29308 0 mod.flipflop21.q
rlabel metal1 20930 28662 20930 28662 0 mod.flipflop22.q
rlabel metal1 21850 29002 21850 29002 0 mod.flipflop23.q
rlabel metal1 22739 25194 22739 25194 0 mod.flipflop24.q
rlabel metal1 21390 26758 21390 26758 0 mod.flipflop25.q
rlabel metal2 21758 30991 21758 30991 0 mod.flipflop26.q
rlabel metal2 23414 25857 23414 25857 0 mod.flipflop27.q
rlabel metal1 18814 26486 18814 26486 0 mod.flipflop28.q
rlabel metal1 12466 31416 12466 31416 0 mod.flipflop29.q
rlabel metal1 20060 29138 20060 29138 0 mod.flipflop30.q
rlabel metal1 22586 30566 22586 30566 0 mod.flipflop31.q
rlabel metal1 18732 28526 18732 28526 0 mod.flipflop32.q
rlabel metal1 18671 29138 18671 29138 0 mod.flipflop33.q
rlabel metal2 23414 27115 23414 27115 0 mod.flipflop34.q
rlabel via1 22034 28475 22034 28475 0 mod.flipflop35.q
rlabel metal1 26434 26282 26434 26282 0 mod.flipflop36.q
rlabel via1 19821 26350 19821 26350 0 mod.flipflop37.q
rlabel metal1 18722 28934 18722 28934 0 mod.flipflop38.q
rlabel metal2 22310 29631 22310 29631 0 mod.flipflop39.q
rlabel metal1 12190 28084 12190 28084 0 mod.flipflop4.d
rlabel metal1 18088 28390 18088 28390 0 mod.flipflop40.q
rlabel metal1 19550 28934 19550 28934 0 mod.flipflop41.q
rlabel via1 12456 29138 12456 29138 0 mod.flipflop42.q
rlabel metal1 21758 24582 21758 24582 0 mod.flipflop43.q
rlabel via2 8510 29291 8510 29291 0 mod.flipflop44.q
rlabel metal3 22034 21964 22034 21964 0 mod.flipflop45.q
rlabel metal1 21344 30022 21344 30022 0 mod.flipflop46.q
rlabel metal2 23414 29886 23414 29886 0 mod.flipflop47.q
rlabel metal1 26818 31246 26818 31246 0 mod.flipflop48.q
rlabel metal2 24656 28356 24656 28356 0 mod.flipflop49.q
rlabel metal3 18469 31484 18469 31484 0 mod.flipflop5.d
rlabel metal2 13754 29665 13754 29665 0 mod.flipflop50.q
rlabel metal1 19324 28118 19324 28118 0 mod.flipflop51.q
rlabel metal1 14766 30090 14766 30090 0 mod.flipflop52.q
rlabel metal2 16790 27897 16790 27897 0 mod.flipflop53.q
rlabel metal2 20102 28101 20102 28101 0 mod.flipflop54.q
rlabel metal1 23240 28050 23240 28050 0 mod.flipflop55.q
rlabel metal2 23874 27370 23874 27370 0 mod.flipflop56.q
rlabel metal1 19044 23018 19044 23018 0 mod.flipflop57.q
rlabel metal1 19366 25466 19366 25466 0 mod.flipflop58.q
rlabel metal1 18676 28186 18676 28186 0 mod.flipflop59.q
rlabel metal4 14628 27200 14628 27200 0 mod.flipflop60.q
rlabel metal2 20746 26367 20746 26367 0 mod.flipflop61.q
rlabel metal3 18952 21692 18952 21692 0 mod.flipflop65.q
rlabel metal1 26235 23766 26235 23766 0 mod.flipflop66.d
rlabel metal1 23736 23086 23736 23086 0 mod.flipflop66.q
rlabel metal1 24150 21658 24150 21658 0 mod.flipflop68.d
rlabel metal1 20378 28390 20378 28390 0 mod.flipflop68.q
rlabel metal1 7406 28730 7406 28730 0 mod.mux15.out
rlabel metal1 20884 27302 20884 27302 0 mod.mux22.out
rlabel metal2 20654 31144 20654 31144 0 mod.mux29.out
rlabel metal1 17112 30362 17112 30362 0 mod.mux36.out
rlabel metal1 16606 29138 16606 29138 0 mod.mux43.out
rlabel metal1 19642 31382 19642 31382 0 mod.mux50.out
rlabel metal1 9430 30702 9430 30702 0 mod.mux57.out
rlabel metal3 17871 27676 17871 27676 0 mod.mux8.out
rlabel metal1 27048 23630 27048 23630 0 net1
rlabel via2 11178 31331 11178 31331 0 net10
rlabel metal2 12006 31263 12006 31263 0 net11
rlabel metal1 10442 31280 10442 31280 0 net12
rlabel metal1 9430 31246 9430 31246 0 net13
rlabel metal3 15916 30600 15916 30600 0 net14
rlabel metal1 2070 31348 2070 31348 0 net15
rlabel metal2 13386 25772 13386 25772 0 net16
rlabel metal1 13478 26894 13478 26894 0 net17
rlabel metal1 24564 31246 24564 31246 0 net18
rlabel metal1 18308 25874 18308 25874 0 net19
rlabel metal1 26542 23086 26542 23086 0 net2
rlabel metal2 24610 25313 24610 25313 0 net20
rlabel metal1 23322 19210 23322 19210 0 net21
rlabel metal2 18814 21182 18814 21182 0 net22
rlabel metal2 22402 17408 22402 17408 0 net23
rlabel metal3 28850 2652 28850 2652 0 net24
rlabel metal2 28382 4845 28382 4845 0 net25
rlabel via2 28382 6749 28382 6749 0 net26
rlabel via2 28382 9061 28382 9061 0 net27
rlabel via2 28382 11101 28382 11101 0 net28
rlabel metal2 28382 13073 28382 13073 0 net29
rlabel metal1 26220 28118 26220 28118 0 net3
rlabel via2 28382 14875 28382 14875 0 net30
rlabel via2 28382 16949 28382 16949 0 net31
rlabel metal2 28382 19057 28382 19057 0 net32
rlabel metal2 28382 21165 28382 21165 0 net33
rlabel via2 28382 23069 28382 23069 0 net34
rlabel metal3 28451 24820 28451 24820 0 net35
rlabel metal3 28911 26996 28911 26996 0 net36
rlabel metal2 29118 29172 29118 29172 0 net37
rlabel metal2 29164 31212 29164 31212 0 net38
rlabel metal2 28382 33252 28382 33252 0 net39
rlabel metal2 23874 28832 23874 28832 0 net4
rlabel metal3 1142 30260 1142 30260 0 net40
rlabel metal3 1142 28220 1142 28220 0 net41
rlabel metal3 1142 26180 1142 26180 0 net42
rlabel metal3 1142 24140 1142 24140 0 net43
rlabel metal3 1142 22100 1142 22100 0 net44
rlabel metal3 1142 20060 1142 20060 0 net45
rlabel metal3 1142 18020 1142 18020 0 net46
rlabel metal3 1142 15980 1142 15980 0 net47
rlabel metal3 1142 13940 1142 13940 0 net48
rlabel metal3 1142 11900 1142 11900 0 net49
rlabel metal1 26220 21658 26220 21658 0 net5
rlabel metal3 1142 9860 1142 9860 0 net50
rlabel metal3 1142 7820 1142 7820 0 net51
rlabel metal3 1142 5780 1142 5780 0 net52
rlabel metal3 1142 3740 1142 3740 0 net53
rlabel via2 28382 3621 28382 3621 0 net54
rlabel via2 28382 5661 28382 5661 0 net55
rlabel metal2 28382 7633 28382 7633 0 net56
rlabel via2 28382 9435 28382 9435 0 net57
rlabel via2 28382 11509 28382 11509 0 net58
rlabel metal2 28382 13617 28382 13617 0 net59
rlabel metal2 23598 18088 23598 18088 0 net6
rlabel metal2 28382 15725 28382 15725 0 net60
rlabel via2 28382 17629 28382 17629 0 net61
rlabel via2 28382 19805 28382 19805 0 net62
rlabel metal2 28382 21777 28382 21777 0 net63
rlabel via2 28382 23715 28382 23715 0 net64
rlabel metal3 28620 25772 28620 25772 0 net65
rlabel metal1 26358 24854 26358 24854 0 net66
rlabel metal3 28942 29852 28942 29852 0 net67
rlabel metal3 27677 31892 27677 31892 0 net68
rlabel metal1 27508 27370 27508 27370 0 net69
rlabel metal1 28704 25942 28704 25942 0 net7
rlabel metal2 23966 33252 23966 33252 0 net70
rlabel metal2 16422 30090 16422 30090 0 net71
rlabel metal1 21114 30124 21114 30124 0 net72
rlabel metal2 13846 32480 13846 32480 0 net73
rlabel metal1 9752 30158 9752 30158 0 net74
rlabel metal1 7176 31314 7176 31314 0 net75
rlabel metal1 3956 31314 3956 31314 0 net76
rlabel metal1 1564 31246 1564 31246 0 net77
rlabel metal3 1142 29580 1142 29580 0 net78
rlabel metal3 1142 27540 1142 27540 0 net79
rlabel metal1 26450 22610 26450 22610 0 net8
rlabel metal3 1142 25500 1142 25500 0 net80
rlabel metal3 1142 23460 1142 23460 0 net81
rlabel metal3 1142 21420 1142 21420 0 net82
rlabel metal3 1142 19380 1142 19380 0 net83
rlabel metal3 1142 17340 1142 17340 0 net84
rlabel metal3 1142 15300 1142 15300 0 net85
rlabel metal3 1142 13260 1142 13260 0 net86
rlabel metal3 1142 11220 1142 11220 0 net87
rlabel metal3 1142 9180 1142 9180 0 net88
rlabel metal3 1142 7140 1142 7140 0 net89
rlabel metal1 9982 30668 9982 30668 0 net9
rlabel metal3 1142 5100 1142 5100 0 net90
rlabel metal3 1142 3060 1142 3060 0 net91
<< properties >>
string FIXED_BBOX 0 0 30000 34000
<< end >>
