magic
tech sky130A
magscale 1 2
timestamp 1672533679
<< obsli1 >>
rect 1104 2159 31832 32657
<< obsm1 >>
rect 934 2128 32996 33516
<< metal2 >>
rect 938 34350 994 35150
rect 2134 34350 2190 35150
rect 3330 34350 3386 35150
rect 4526 34350 4582 35150
rect 5722 34350 5778 35150
rect 6918 34350 6974 35150
rect 8114 34350 8170 35150
rect 9310 34350 9366 35150
rect 10506 34350 10562 35150
rect 11702 34350 11758 35150
rect 12898 34350 12954 35150
rect 14094 34350 14150 35150
rect 15290 34350 15346 35150
rect 16486 34350 16542 35150
rect 17682 34350 17738 35150
rect 18878 34350 18934 35150
rect 20074 34350 20130 35150
rect 21270 34350 21326 35150
rect 22466 34350 22522 35150
rect 23662 34350 23718 35150
rect 24858 34350 24914 35150
rect 26054 34350 26110 35150
rect 27250 34350 27306 35150
rect 28446 34350 28502 35150
rect 29642 34350 29698 35150
rect 30838 34350 30894 35150
rect 32034 34350 32090 35150
<< obsm2 >>
rect 1050 34294 2078 34921
rect 2246 34294 3274 34921
rect 3442 34294 4470 34921
rect 4638 34294 5666 34921
rect 5834 34294 6862 34921
rect 7030 34294 8058 34921
rect 8226 34294 9254 34921
rect 9422 34294 10450 34921
rect 10618 34294 11646 34921
rect 11814 34294 12842 34921
rect 13010 34294 14038 34921
rect 14206 34294 15234 34921
rect 15402 34294 16430 34921
rect 16598 34294 17626 34921
rect 17794 34294 18822 34921
rect 18990 34294 20018 34921
rect 20186 34294 21214 34921
rect 21382 34294 22410 34921
rect 22578 34294 23606 34921
rect 23774 34294 24802 34921
rect 24970 34294 25998 34921
rect 26166 34294 27194 34921
rect 27362 34294 28390 34921
rect 28558 34294 29586 34921
rect 29754 34294 30782 34921
rect 30950 34294 31978 34921
rect 32146 34294 32996 34921
rect 940 711 32996 34294
<< metal3 >>
rect 0 34144 800 34264
rect 0 33328 800 33448
rect 0 32512 800 32632
rect 32206 32376 33006 32496
rect 0 31696 800 31816
rect 32206 31696 33006 31816
rect 0 30880 800 31000
rect 32206 31016 33006 31136
rect 32206 30336 33006 30456
rect 0 30064 800 30184
rect 32206 29656 33006 29776
rect 0 29248 800 29368
rect 32206 28976 33006 29096
rect 0 28432 800 28552
rect 32206 28296 33006 28416
rect 0 27616 800 27736
rect 32206 27616 33006 27736
rect 0 26800 800 26920
rect 32206 26936 33006 27056
rect 32206 26256 33006 26376
rect 0 25984 800 26104
rect 32206 25576 33006 25696
rect 0 25168 800 25288
rect 32206 24896 33006 25016
rect 0 24352 800 24472
rect 32206 24216 33006 24336
rect 0 23536 800 23656
rect 32206 23536 33006 23656
rect 0 22720 800 22840
rect 32206 22856 33006 22976
rect 32206 22176 33006 22296
rect 0 21904 800 22024
rect 32206 21496 33006 21616
rect 0 21088 800 21208
rect 32206 20816 33006 20936
rect 0 20272 800 20392
rect 32206 20136 33006 20256
rect 0 19456 800 19576
rect 32206 19456 33006 19576
rect 0 18640 800 18760
rect 32206 18776 33006 18896
rect 32206 18096 33006 18216
rect 0 17824 800 17944
rect 32206 17416 33006 17536
rect 0 17008 800 17128
rect 32206 16736 33006 16856
rect 0 16192 800 16312
rect 32206 16056 33006 16176
rect 0 15376 800 15496
rect 32206 15376 33006 15496
rect 0 14560 800 14680
rect 32206 14696 33006 14816
rect 32206 14016 33006 14136
rect 0 13744 800 13864
rect 32206 13336 33006 13456
rect 0 12928 800 13048
rect 32206 12656 33006 12776
rect 0 12112 800 12232
rect 32206 11976 33006 12096
rect 0 11296 800 11416
rect 32206 11296 33006 11416
rect 0 10480 800 10600
rect 32206 10616 33006 10736
rect 32206 9936 33006 10056
rect 0 9664 800 9784
rect 32206 9256 33006 9376
rect 0 8848 800 8968
rect 32206 8576 33006 8696
rect 0 8032 800 8152
rect 32206 7896 33006 8016
rect 0 7216 800 7336
rect 32206 7216 33006 7336
rect 0 6400 800 6520
rect 32206 6536 33006 6656
rect 32206 5856 33006 5976
rect 0 5584 800 5704
rect 32206 5176 33006 5296
rect 0 4768 800 4888
rect 32206 4496 33006 4616
rect 0 3952 800 4072
rect 32206 3816 33006 3936
rect 0 3136 800 3256
rect 32206 3136 33006 3256
rect 0 2320 800 2440
rect 32206 2456 33006 2576
rect 0 1504 800 1624
rect 0 688 800 808
<< obsm3 >>
rect 800 34344 32831 34917
rect 880 34064 32831 34344
rect 800 33528 32831 34064
rect 880 33248 32831 33528
rect 800 32712 32831 33248
rect 880 32576 32831 32712
rect 880 32432 32126 32576
rect 800 32296 32126 32432
rect 800 31896 32831 32296
rect 880 31616 32126 31896
rect 800 31216 32831 31616
rect 800 31080 32126 31216
rect 880 30936 32126 31080
rect 880 30800 32831 30936
rect 800 30536 32831 30800
rect 800 30264 32126 30536
rect 880 30256 32126 30264
rect 880 29984 32831 30256
rect 800 29856 32831 29984
rect 800 29576 32126 29856
rect 800 29448 32831 29576
rect 880 29176 32831 29448
rect 880 29168 32126 29176
rect 800 28896 32126 29168
rect 800 28632 32831 28896
rect 880 28496 32831 28632
rect 880 28352 32126 28496
rect 800 28216 32126 28352
rect 800 27816 32831 28216
rect 880 27536 32126 27816
rect 800 27136 32831 27536
rect 800 27000 32126 27136
rect 880 26856 32126 27000
rect 880 26720 32831 26856
rect 800 26456 32831 26720
rect 800 26184 32126 26456
rect 880 26176 32126 26184
rect 880 25904 32831 26176
rect 800 25776 32831 25904
rect 800 25496 32126 25776
rect 800 25368 32831 25496
rect 880 25096 32831 25368
rect 880 25088 32126 25096
rect 800 24816 32126 25088
rect 800 24552 32831 24816
rect 880 24416 32831 24552
rect 880 24272 32126 24416
rect 800 24136 32126 24272
rect 800 23736 32831 24136
rect 880 23456 32126 23736
rect 800 23056 32831 23456
rect 800 22920 32126 23056
rect 880 22776 32126 22920
rect 880 22640 32831 22776
rect 800 22376 32831 22640
rect 800 22104 32126 22376
rect 880 22096 32126 22104
rect 880 21824 32831 22096
rect 800 21696 32831 21824
rect 800 21416 32126 21696
rect 800 21288 32831 21416
rect 880 21016 32831 21288
rect 880 21008 32126 21016
rect 800 20736 32126 21008
rect 800 20472 32831 20736
rect 880 20336 32831 20472
rect 880 20192 32126 20336
rect 800 20056 32126 20192
rect 800 19656 32831 20056
rect 880 19376 32126 19656
rect 800 18976 32831 19376
rect 800 18840 32126 18976
rect 880 18696 32126 18840
rect 880 18560 32831 18696
rect 800 18296 32831 18560
rect 800 18024 32126 18296
rect 880 18016 32126 18024
rect 880 17744 32831 18016
rect 800 17616 32831 17744
rect 800 17336 32126 17616
rect 800 17208 32831 17336
rect 880 16936 32831 17208
rect 880 16928 32126 16936
rect 800 16656 32126 16928
rect 800 16392 32831 16656
rect 880 16256 32831 16392
rect 880 16112 32126 16256
rect 800 15976 32126 16112
rect 800 15576 32831 15976
rect 880 15296 32126 15576
rect 800 14896 32831 15296
rect 800 14760 32126 14896
rect 880 14616 32126 14760
rect 880 14480 32831 14616
rect 800 14216 32831 14480
rect 800 13944 32126 14216
rect 880 13936 32126 13944
rect 880 13664 32831 13936
rect 800 13536 32831 13664
rect 800 13256 32126 13536
rect 800 13128 32831 13256
rect 880 12856 32831 13128
rect 880 12848 32126 12856
rect 800 12576 32126 12848
rect 800 12312 32831 12576
rect 880 12176 32831 12312
rect 880 12032 32126 12176
rect 800 11896 32126 12032
rect 800 11496 32831 11896
rect 880 11216 32126 11496
rect 800 10816 32831 11216
rect 800 10680 32126 10816
rect 880 10536 32126 10680
rect 880 10400 32831 10536
rect 800 10136 32831 10400
rect 800 9864 32126 10136
rect 880 9856 32126 9864
rect 880 9584 32831 9856
rect 800 9456 32831 9584
rect 800 9176 32126 9456
rect 800 9048 32831 9176
rect 880 8776 32831 9048
rect 880 8768 32126 8776
rect 800 8496 32126 8768
rect 800 8232 32831 8496
rect 880 8096 32831 8232
rect 880 7952 32126 8096
rect 800 7816 32126 7952
rect 800 7416 32831 7816
rect 880 7136 32126 7416
rect 800 6736 32831 7136
rect 800 6600 32126 6736
rect 880 6456 32126 6600
rect 880 6320 32831 6456
rect 800 6056 32831 6320
rect 800 5784 32126 6056
rect 880 5776 32126 5784
rect 880 5504 32831 5776
rect 800 5376 32831 5504
rect 800 5096 32126 5376
rect 800 4968 32831 5096
rect 880 4696 32831 4968
rect 880 4688 32126 4696
rect 800 4416 32126 4688
rect 800 4152 32831 4416
rect 880 4016 32831 4152
rect 880 3872 32126 4016
rect 800 3736 32126 3872
rect 800 3336 32831 3736
rect 880 3056 32126 3336
rect 800 2656 32831 3056
rect 800 2520 32126 2656
rect 880 2376 32126 2520
rect 880 2240 32831 2376
rect 800 1704 32831 2240
rect 880 1424 32831 1704
rect 800 888 32831 1424
rect 880 715 32831 888
<< metal4 >>
rect 4785 2128 5105 32688
rect 8626 2128 8946 32688
rect 12467 2128 12787 32688
rect 16308 2128 16628 32688
rect 20149 2128 20469 32688
rect 23990 2128 24310 32688
rect 27831 2128 28151 32688
rect 31672 2128 31992 32688
<< obsm4 >>
rect 5395 32768 32693 34917
rect 5395 4659 8546 32768
rect 9026 4659 12387 32768
rect 12867 4659 16228 32768
rect 16708 4659 20069 32768
rect 20549 4659 23910 32768
rect 24390 4659 27751 32768
rect 28231 4659 31592 32768
rect 32072 4659 32693 32768
<< labels >>
rlabel metal3 s 32206 2456 33006 2576 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 32206 22856 33006 22976 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 32206 24896 33006 25016 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 32206 26936 33006 27056 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 32206 28976 33006 29096 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 32206 31016 33006 31136 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 32034 34350 32090 35150 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 28446 34350 28502 35150 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 24858 34350 24914 35150 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 21270 34350 21326 35150 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 17682 34350 17738 35150 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 32206 4496 33006 4616 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 14094 34350 14150 35150 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 10506 34350 10562 35150 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 6918 34350 6974 35150 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 3330 34350 3386 35150 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 32206 6536 33006 6656 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 32206 8576 33006 8696 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 32206 10616 33006 10736 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 32206 12656 33006 12776 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 32206 14696 33006 14816 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 32206 16736 33006 16856 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 32206 18776 33006 18896 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 32206 20816 33006 20936 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 32206 3816 33006 3936 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 32206 24216 33006 24336 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 32206 26256 33006 26376 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 32206 28296 33006 28416 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 32206 30336 33006 30456 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 32206 32376 33006 32496 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 29642 34350 29698 35150 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 26054 34350 26110 35150 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 22466 34350 22522 35150 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 18878 34350 18934 35150 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 15290 34350 15346 35150 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 32206 5856 33006 5976 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 11702 34350 11758 35150 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 8114 34350 8170 35150 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 4526 34350 4582 35150 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 938 34350 994 35150 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 32206 7896 33006 8016 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 688 800 808 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 32206 9936 33006 10056 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 32206 11976 33006 12096 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 32206 14016 33006 14136 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 32206 16056 33006 16176 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 32206 18096 33006 18216 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 32206 20136 33006 20256 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 32206 22176 33006 22296 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 32206 3136 33006 3256 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 32206 23536 33006 23656 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 32206 25576 33006 25696 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 32206 27616 33006 27736 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 32206 29656 33006 29776 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 32206 31696 33006 31816 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 30838 34350 30894 35150 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 27250 34350 27306 35150 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 23662 34350 23718 35150 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 20074 34350 20130 35150 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 16486 34350 16542 35150 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 32206 5176 33006 5296 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 12898 34350 12954 35150 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 9310 34350 9366 35150 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 5722 34350 5778 35150 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 2134 34350 2190 35150 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 32206 7216 33006 7336 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 32206 9256 33006 9376 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 32206 11296 33006 11416 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 32206 13336 33006 13456 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 32206 15376 33006 15496 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 32206 17416 33006 17536 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 32206 19456 33006 19576 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 32206 21496 33006 21616 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 4785 2128 5105 32688 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 12467 2128 12787 32688 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 20149 2128 20469 32688 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 27831 2128 28151 32688 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 8626 2128 8946 32688 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 16308 2128 16628 32688 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 23990 2128 24310 32688 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 31672 2128 31992 32688 6 vssd1
port 116 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 33006 35150
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4024100
string GDS_FILE /home/runner/work/tiny_user_project_vgaclock_mpw8/tiny_user_project_vgaclock_mpw8/openlane/tiny_user_project/runs/22_12_31_22_51/results/signoff/tiny_user_project.magic.gds
string GDS_START 509702
<< end >>

